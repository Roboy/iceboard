// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Jan 31 15:26:06 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, INHC_c, INLB_c, INHB_c, 
        INLA_c, INHA_c;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(125[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(127[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(128[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(129[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(130[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(131[22:24])
    
    wire n37492;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(133[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(134[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(135[22:35])
    
    wire n37491, n37168;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(165[22:33])
    
    wire n516;
    wire [7:0]data;   // verilog/TinyFPGA_B.v(228[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(252[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(260[15:20])
    
    wire n49422;
    wire [22:0]pwm_setpoint_22__N_11;
    
    wire RX_N_10;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(124[11:28])
    
    wire n1152;
    wire [31:0]motor_state_23__N_106;
    wire [32:0]encoder0_position_scaled_23__N_34;
    
    wire encoder1_position_scaled_23__N_231;
    wire [31:0]encoder1_position_scaled_23__N_58;
    wire [23:0]displacement_23__N_82;
    
    wire n659, n660, n661, n662, n663, n664, n665, n666, n667, 
        n668, n669, n670, n671, n672, n673, n674, n675, n676, 
        n677, n678, n679, n680, n681, n682, n683, n684, n685, 
        n686, n687, n688, n689, n690, read_N_321, n777, n37490, 
        n37489, n37488, n1193;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(126[11:28])
    
    wire n37487;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n37486, n28292, n28291, n28290, n28289, n28288, n28287, 
        n28286, n28285, n28284, n28283, n28282, n49129, n37485, 
        n37484, n37483, n37482, n37481, n37480, n4227, n37479, 
        n26652, n37478, n43217, n33700, n48495, n33696, n26487, 
        n2, n15, n34613, n28281, n28280, n28279, n28278;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n15_adj_4947, n37477, n37476, n28277, n28276, n3, n4, 
        n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15_adj_4948, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n37475, n49552, n19247;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire tx_active, n40598, n43254, n37474, n48033, n49181, n49096, 
        n28275, n48424, n37184, n37473, n37472, n37471, n37183, 
        n14_adj_4949, n10_adj_4950, n37470, n25_adj_4951, n17_adj_4952, 
        n44198, n5_adj_4953, n6_adj_4954, n7_adj_4955, n8_adj_4956, 
        n9_adj_4957, n10_adj_4958, n11_adj_4959, n12_adj_4960, n13_adj_4961, 
        n14_adj_4962, n15_adj_4963, n16_adj_4964, n17_adj_4965, n18_adj_4966, 
        n19_adj_4967, n20_adj_4968, n21_adj_4969, n22_adj_4970, n23_adj_4971, 
        n24_adj_4972, n25_adj_4973, n37469, n37167, n37468, n37467, 
        n37466, n37465, n37464, n37463, n37462, n37182, n47990, 
        n43213, n37461, n37460, n38496, n38495, n38494, n38493, 
        n38492, n38491, n38490, n34679, n38489, n38488, n38487, 
        n38486, n38485, n38484, n38483, n38482, n43603, n38481, 
        n38480, n38479, n37459, n38478, n38477, n38476, n38475, 
        n38474, n38473, n37458, n37457, n38472, n38471, n38470, 
        n38469, n38468, n38467, n38466, n38465, n38464, n38463, 
        n38462, n38461, n38460, n38459, n38458, n38457, n38456, 
        n38455, n38454, n38453, n38452, n38451, n38450, n38449, 
        n38448, n38447, n38446, n38445, n38444, n37166, n38443, 
        n38442, n37456, n38441, n38440, n38439, n38438, n43181, 
        n38437, n38436, n38435, n37455, n38434, n38433, n38432, 
        n38431, n38430, n38429, n43134, n38428, n49248, n41391, 
        n38427, n38426, n12_adj_4974, n38425, n38424, n38423, n38422, 
        n37454, n37453, n15_adj_4975, n14_adj_4976, n37214, n37452, 
        n38421, n37451, n37450, n38420, n38419, n38418, n38417, 
        n34637, n38416, n38415, n38414, n38413, n38412, n38411, 
        n38410, n38409, n38408, n10_adj_4977, n28274, n4_adj_4978, 
        n38407, n38406, n38405, n38404, n38403, n38402, n30301, 
        n38401, n38400, n38399, n38398, n37213, n38397, n38396, 
        n38668, n38395, n38394, n38393, n38392, n34533, n38391, 
        n38673, n38677, n38390, n38389, n34627, n38388, n38387, 
        n38386, n37181, n38385, n38384, n38383, n48286, n49036, 
        n38382, n38381, n38380, n38379, n38378, n38377, n38376, 
        n38375, n38374, n38373, n38372, n38371, n38370, n38369, 
        n38368, n38367, n38366, n38365, n38364, n38363, n38362, 
        n43242, n12_adj_4979, n38361, n4_adj_4980, n4_adj_4981, n43610, 
        n38360, n38359, n34379, n34377, n34373, n34365, n34363, 
        n34313, n34481, n38358, n34306, n38357, n38356, n38355, 
        n38354, n38353, n38352, n38351, n38350, n38349, n38348, 
        n38347, n38346, n38345, n38344, n38343, n38342, n38341, 
        n38340, n38339, n38338, n38337, n38336, n38335, n38334, 
        n38333, n38332, n38331, n38330, n38329, n38328, n38327, 
        n38326, n38325, n42790, n38324, n38323, n38322, n28747, 
        n28746, n28745, n28744, n28743, n28742, n28741, n28738, 
        n28737, n48769, n8_adj_4982, n28736, n7_adj_4983, n28735, 
        n28734, n28733, n28732, n28731, n28730, n28729, n28728, 
        n28727, n28726, n28725, n28724, n28723, n28722, n28721, 
        n28720, n28719, n28718, n28717, n28716, n28715, n28714, 
        n28713, n28712, n28711, n28710, n28709, n28708, n28707, 
        n28706, n28705, n28704, n4_adj_4984, n28703, n38321, n38320, 
        n38319, n38318, n38317, n38316, n28702, n33, n32, n31, 
        n30, n29, n28, n27, n26, n25_adj_4985, n24_adj_4986, n23_adj_4987, 
        n22_adj_4988, n21_adj_4989, n20_adj_4990, n19_adj_4991, n18_adj_4992, 
        n17_adj_4993, n16_adj_4994, n15_adj_4995, n14_adj_4996, n13_adj_4997, 
        n12_adj_4998, n11_adj_4999, n10_adj_5000, n9_adj_5001, n8_adj_5002, 
        n7_adj_5003, n28701, n28700, n38315, n28698, n28697, n28696, 
        n28695, n28694, n28693, n28692, n3_adj_5004, n4_adj_5005, 
        n28691, n28690, n28689, n28688, n28687, n28686, n28685, 
        n5722, n28684, n28273, n28272, n28271, n28270, n28269, 
        n28268, n28267, n28266, n28265, n28264, n28263, n28262, 
        n28261, n28260, n28259, n28258, n28257, n28256, n28255, 
        n28254, n28253, n28252, n28251, n28250, n28249, n28248, 
        n28247, n28246, n28245, n28244, n28243, n28242, n28241, 
        n28683, n38314, n28682, n28681, n28680, n28679, n28678, 
        n28677, n28676, n28675, n28674, n28673, n28672, n38313, 
        n38312, n28671, n28670, n28669, n28668, n28667, n28666, 
        n28665, n28664, n28663, n28662, n38311, n28661, n28660, 
        n28659, n38310, n28658, n28657, n28656, n28655, n7_adj_5006, 
        n28654, n28653, n28652, n28651, n28650, n28649, n28648, 
        n28647, n28646, n28645, n28644, n28643, n26489, n28642, 
        n28641, n28640, n28639, n28638, n28637, n28636, n28635, 
        n28634, n28633, n28632, n28631, n28630, n28629, n28628, 
        n28627, n28626, n28625, n38309, n4_adj_5007, n5_adj_5008, 
        n38308, n28624, n28623, n28622, n28621, n28620, n28619, 
        n28618, n28617, n28616, n28615, n28614, n28613, n28612, 
        n28611, n28610, n28609, n28608, n28607, n4_adj_5009, n28606, 
        n28605, n28604, n28603, n28602, n28601, n28600;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n28599, n28598, n28597, n28596, n28595, n28594, 
        n28593, n28592, n28591, n28590, n28589, n28588, n28587, 
        n28586, n28585, n28584, n28583, n28582, n28581, n28580, 
        n28579, n28578, direction_N_3807, n28577, n28576, n28575, 
        n28574, n28573, n28572, n28571, n28570, n28569, n28568, 
        n28567, n28566, n28565, n28564, n28563, n28562, n28561, 
        n28560, n28559, n28558, n28557, n28556, n38298, n28555, 
        n28240, n28239, n28554, n28238, n28237, n28236, n28235, 
        n28234, n28233, n28232, n28553, n28552;
    wire [1:0]a_new_adj_5130;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_5011, n28551, n28550, n28549, n28548, n28547, 
        n28546, n28545, n28544, n1419, n2380, n38297, n28543, 
        n28542, n28541, n48206, direction_N_3807_adj_5012, n28539, 
        n38296, n38295, n28538, n4_adj_5013, n28537, n28536, n28535, 
        n28534, n28533, n28532, n28531, n28530, n28529, n28528, 
        n38294, n5855, n38293, n28527, n28526, n6014, n38292, 
        n28525, n28524, n43196, n38291, n28523, n38290, n28522, 
        n28521, n38289, n28224, n28221, n28216, n28215, n28212, 
        n41841, n28520, rw;
    wire [7:0]state_adj_5154;   // verilog/eeprom.v(23[11:16])
    
    wire n28519, n28518, n5_adj_5016, n28517, n28516, n28515, n28514, 
        n5_adj_5017, n38288, n28513, n28512, n28511, n28510, n28509, 
        n28508, n28507, n28506, n38287, n38286, n28505, n28504, 
        n6_adj_5018, n5_adj_5019, n4_adj_5020, n3_adj_5021, n2_adj_5022, 
        r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n38285, n28503, n38284, n38283, n38282, n38281, n42126, 
        n38280, n38279, n28502, n28501;
    wire [2:0]r_SM_Main_2__N_3442;
    
    wire n28500, n28499, n28498, n38278, n38277, n28497, n28496, 
        n28495, n28494, n28493, n28492, n28491, n28490, n28489, 
        n28488, n28487, n28486, n34597;
    wire [2:0]r_SM_Main_adj_5161;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5163;   // verilog/uart_tx.v(33[16:27])
    
    wire n38276, n38275;
    wire [2:0]r_SM_Main_2__N_3513;
    
    wire n38274, n28485, n28484, n38273, n28104, n28483, n28482, 
        n38272, n38271, n38270, n28481, n28480, n28479, n28478, 
        n28477, n28476, n28475, n34595, n38269, n38268, n38267, 
        n28474, n28473, n28472, n28471, n28470, n28469, n28468, 
        n28467, n28466, n28465, n28464, n38266;
    wire [7:0]state_adj_5170;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n38265, n38264, n4_adj_5028, enable_slow_N_4090, n38263, 
        n38262, n34593, n38261, n38260, n38259;
    wire [7:0]state_7__N_3987;
    
    wire n38258, n5538, n38257, n38256, n38255, n38659, n38254;
    wire [7:0]state_7__N_4003;
    
    wire n38661, n38253, n38252, n38251, n38250, n38249, n38248, 
        n38247, n38246, n38245, n38244, n38243, n38242, n28202, 
        n38241, n38663, n621, n622, n623, n625, n626, n627, 
        n628, n629, n630, n631, n632, n633, n634, n635, n636, 
        n637, n638, n639, n640, n641, n642, n643, n644, n645, 
        n646, n647, n648, n649, n650, n651, n652, n38240, n38239, 
        n38238, n38237, n38236, n38235, n38234, n38233, n6542, 
        n6541, n6540, n6539, n6538, n6537, n38232, n828, n829, 
        n830, n831, n832, n833, n38231, n861, n896, n897, n898, 
        n899, n900, n901, n927, n928, n929, n930, n931, n932, 
        n933, n38230, n960, n48208, n995, n996, n997, n998, 
        n999, n1000, n1001, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n38229, n1059, n38665, n1093, n1094, 
        n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1125, 
        n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
        n1158, n1193_adj_5029, n1194, n1195, n1196, n1197, n1198, 
        n1199, n1200, n1201, n1224, n1225, n1226, n1227, n1228, 
        n1229, n1230, n1231, n1232, n1233, n1257, n1292, n1293, 
        n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
        n38228, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
        n1330, n1331, n1332, n1333, n1356, n1391, n1392, n1393, 
        n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
        n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
        n1430, n1431, n1432, n1433, n38227, n1455, n1490, n1491, 
        n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
        n1500, n1501, n1521, n1522, n1523, n1524, n1525, n1526, 
        n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1554, 
        n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
        n1597, n1598, n1599, n1600, n1601, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n1653, n41955, n1688, n1689, n1690, 
        n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
        n1699, n1700, n1701, n38226, n38225, n38666, n1719, n1720, 
        n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
        n1729, n1730, n1731, n1732, n1733, n1752, n38670, n38224, 
        n34587, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
        n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
        n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
        n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
        n38223, n1851, n38222, n1886, n1887, n1888, n1889, n1890, 
        n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
        n1899, n1900, n1901, n1917, n1918, n1919, n1920, n1921, 
        n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
        n1930, n1931, n1932, n1933, n38221, n27824, n1950, n27820, 
        n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
        n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
        n2001, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
        n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
        n2031, n2032, n2033, n2049, n38220, n2084, n2085, n2086, 
        n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
        n2095, n2096, n2097, n2098, n2099, n2100, n2101, n38219, 
        n38218, n2115, n2116, n2117, n2118, n2119, n2120, n2121, 
        n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
        n2130, n2131, n2132, n2133, n2148, n34583, n38217, n43150, 
        n38216, n6_adj_5030, n2183, n2184, n2185, n2186, n2187, 
        n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, 
        n2196, n2197, n2198, n2199, n2200, n2201, n2214, n2215, 
        n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, 
        n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, 
        n2232, n2233, n2247, n38675, n2282, n2283, n2284, n2285, 
        n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
        n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
        n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
        n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
        n2329, n2330, n2331, n2332, n2333, n2346, n38215, n46578, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n2445, n2480, n2481, n2482, n2483, 
        n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, 
        n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
        n2500, n2501, n2511, n2512, n2513, n2514, n2515, n2516, 
        n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
        n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
        n2533, n2544, n2579, n2580, n2581, n2582, n2583, n2584, 
        n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
        n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
        n2601, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
        n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
        n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
        n2633, n48618, n2643, n27784, n2678, n2679, n2680, n2681, 
        n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
        n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
        n2698, n2699, n2700, n2701, n2709, n2710, n2711, n2712, 
        n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
        n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
        n2729, n2730, n2731, n2732, n2733, n2742, n2777, n2778, 
        n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
        n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, 
        n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2808, 
        n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
        n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, 
        n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
        n2833, n2841, n43139, n2876, n2877, n2878, n2879, n2880, 
        n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
        n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
        n2897, n2898, n2899, n2900, n2901, n2907, n2908, n2909, 
        n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, 
        n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
        n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
        n2940, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
        n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
        n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
        n2998, n2999, n3000, n3001, n3006, n3007, n3008, n3009, 
        n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
        n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
        n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
        n3039, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
        n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
        n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, 
        n3096, n3097, n3098, n3099, n3100, n3101, n3105, n3106, 
        n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, 
        n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
        n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, 
        n3131, n3132, n3133, n49040, n3138, n3173, n3174, n3175, 
        n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
        n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
        n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
        n3200, n3201, n3204, n3205, n3206, n3207, n3208, n3209, 
        n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, 
        n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, 
        n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
        n49074, n3237, n3272, n3273, n3274, n3275, n3276, n3277, 
        n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, 
        n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
        n3294, n3295, n3296, n3298, n3299, n3300, n3301, n38214, 
        n38213, n38212, n49368, n49365, n24_adj_5031, n27753, n27752, 
        n62, n26514, n26517, n38211, n26499, n48037, n48229, n38210, 
        n38209, n6_adj_5032, n49002, n48039, n48228, n28195, n28194, 
        n4_adj_5033, n6_adj_5034, n7_adj_5035, n8_adj_5036, n9_adj_5037, 
        n10_adj_5038, n11_adj_5039, n12_adj_5040, n13_adj_5041, n15_adj_5042, 
        n17_adj_5043, n19_adj_5044, n21_adj_5045, n23_adj_5046, n48425, 
        n25_adj_5047, n27_adj_5048, n48370, n29_adj_5049, n30_adj_5050, 
        n31_adj_5051, n33_adj_5052, n48750, n35, n26497, n38649, 
        n45658, n28192, n28191, n26511, n28189, n28188, n45650, 
        n45644, n48366, n48731, n48023, n45638, n45632, n45630, 
        n42123, n42230, n45624, n45620, n45618, n38656, n45604, 
        n12_adj_5053, n45598, n44442, n43224, n45590, n45584, n14_adj_5054, 
        n10_adj_5055, n45578, n45574, n45572, n28187, n28405, n28403, 
        n28402, n28401, n28400, n28399, n28398, n28397, n43159, 
        n49231, n38679, n28186, n28185, n28184, n28183, n28182, 
        n28181, n28180, n28179, n28178, n28177, n28176, n28174, 
        n28170, n28169, n34577, n49207, n45554, n45548, n48717, 
        n12_adj_5056, n34575, n2_adj_5057, n3_adj_5058, n4_adj_5059, 
        n5_adj_5060, n6_adj_5061, n7_adj_5062, n8_adj_5063, n9_adj_5064, 
        n10_adj_5065, n11_adj_5066, n12_adj_5067, n13_adj_5068, n14_adj_5069, 
        n15_adj_5070, n16_adj_5071, n17_adj_5072, n18_adj_5073, n19_adj_5074, 
        n20_adj_5075, n21_adj_5076, n22_adj_5077, n23_adj_5078, n24_adj_5079, 
        n25_adj_5080, n26_adj_5081, n27_adj_5082, n28_adj_5083, n29_adj_5084, 
        n30_adj_5085, n31_adj_5086, n32_adj_5087, n33_adj_5088, n48371, 
        n45542, n41845, n43073, n37180, n38091, n38090, n34557, 
        n38089, n38088, n38087, n43002, n38086, n38085, n38084, 
        n38083, n38082, n38081, n8_adj_5089, n38080, n38079, n38078, 
        n38077, n38076, n38075, n45536, n42897, n38074, n38073, 
        n38072, n45534, n46660, n45526, n48696, n37212, n34525, 
        n48968, n45518, n45512, n37211, n37179, n45506, n45504, 
        n47614, n45498, n42957, n42955, n42953, n42951, n42948, 
        n45496, n34515, n45494, n28168, n37990, n37989, n37988, 
        n37987, n38667, n37986, n37985, n38671, n37210, n37984, 
        n37983, n37982, n37981, n37980, n37979, n37978, n38672, 
        n37977, n37209, n37976, n38676, n37975, n37974, n37973, 
        n37972, n37971, n37970, n37178, n37969, n37968, n45474, 
        n37165, n37967, n37966, n37965, n37964, n37963, n37962, 
        n37961, n37960, n37959, n37958, n37957, n37956, n45468, 
        n37955, n37954, n37953, n37952, n37951, n37950, n45464, 
        n37949, n37948, n37947, n37551, n37946, n37208, n37945, 
        n37550, n37944, n37207, n37943, n37942, n37941, n37940, 
        n37939, n37549, n37938, n37937, n45458, n37936, n47726, 
        n37935, n37548, n45456, n37934, n37177, n37176, n37933, 
        n38650, n37547, n37932, n37931, n37930, n37929, n37928, 
        n37927, n37926, n37925, n37924, n37206, n38651, n37205, 
        n46605, n38652, n38653, n37204, n34501, n38657, n49153, 
        n37923, n37922, n37921, n46598, n37920, n38658, n37919, 
        n48297, n37918, n38660, n34551, n47597, n38662, n37917, 
        n37916, n37915, n37914, n37913, n13_adj_5090, n15_adj_5091, 
        n17_adj_5092, n38664, n19_adj_5093, n21_adj_5094, n34491, 
        n23_adj_5095, n27_adj_5096, n37175, n38669, n43, n37912, 
        n38674, n37203, n59, n48936, n61, n37202, n37911, n46594, 
        n45440, n41813, n45434, n45428, n45424, n37201, n45416, 
        n46588, n45408, n45402, n44044, n46544, n37910, n37909, 
        n44222, n45396, n42541, n45392, n45386, n37908, n37907, 
        n37906, n38678, n37905, n37200, n45376, n34487, n37904, 
        n37903, n37902, n37901, n45370, n45366, n37900, n37899, 
        n48497, n37898, n37897, n37896, n37895, n37894, n37893, 
        n45356, n37174, n45350, n45344, n10_adj_5097, n37892, n48904, 
        n33499, n45332, n26628, n45326, n45318, n45316, n45310, 
        n45308, n47573, n45300, n45290, n26607, n45286, n43755, 
        n47693, n45274, n45270, n37164, n37199, n42229, n45264, 
        n45256, n45250, n45248, n42185, n48859, n37881, n37173, 
        n45242, n45240, n45230, n45224, n42949, n37172, n37880, 
        n37879, n37878, n37877, n37876, n37875, n37874, n37873, 
        n37872, n37871, n47691, n37870, n37869, n47683, n37868, 
        n37867, n37866, n37865, n37864, n37863, n37862, n37861, 
        n37860, n47676, n37859, n37858, n37857, n37856, n37855, 
        n37854, n37853, n37852, n37851, n37850, n37849, n37848, 
        n37847, n37846, n37845, n37844, n37843, n37842, n37841, 
        n37840, n37839, n37838, n37837, n37836, n45218, n37825, 
        n37824, n37823, n37822, n37821, n37820, n37819, n37818, 
        n37817, n37816, n37815, n37814, n37813, n37812, n37811, 
        n37810, n37809, n37808, n37807, n37806, n37805, n37804, 
        n37803, n37802, n45212, n45210, n42551, n45196, n45194, 
        n45188, n48562, n45184, n48496, n37198, n28167, n28166, 
        n28165, n28164, n45174, n45168, n37197, n37196, n45164, 
        n48831, n37163, n45158, n45156, n34571, n45144, n45142, 
        n7_adj_5098, n45140, n45138, n45136, n45134, n45132, n37171, 
        n45130, n45126, n45124, n37195, n45122, n37194, n37193, 
        n37192, n45118, n34447, n45112, n45110, n37191, n47538, 
        n37190, n48439, n37189, n45106, n45104, n45102, n37162, 
        n34439, n45100, n46486, n45094, n45088, n28163, n48478, 
        n45082, n26633, n45072, n37170, n45066, n38654, n37161, 
        n37710, n38655, n37709, n37708, n37707, n45060, n26657, 
        n37706, n37705, n45054, n37188, n23943, n37187, n45048, 
        n45046, n48808, n34507, n45044, n37169, n48288, n45026, 
        n37186, n44886, n45020, n45014, n45012, n47524, n45006, 
        n47523, n45002, n45000, n48291, n44870, n44988, n43282, 
        n37185, n44978, n27554, n44972, n48787, n47518, n43131, 
        n37494, n26488, n44966, n37493;
    
    VCC i2 (.Y(VCC_net));
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_58 (.Q(INLB_c), .C(CLK_c), .D(hall3));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n38079), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[0]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4003[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_82[0]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n38079), .I0(n2226), 
            .I1(VCC_net), .CO(n38080));
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n38222), .I0(n2320), 
            .I1(VCC_net), .CO(n38223));
    SB_LUT4 add_29_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n37163), .O(n687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF h2_57 (.Q(INHB_c), .C(CLK_c), .D(hall2));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n38078), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .CLK_c(CLK_c), .n34515(n34515), .\state[1] (state[1]), .\state[0] (state[0]), 
            .GND_net(GND_net), .n2380(n2380), .n30301(n30301), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n28262(n28262), .neopxl_color({neopxl_color}), .n28261(n28261), 
            .n28260(n28260), .n28259(n28259), .n28258(n28258), .n28257(n28257), 
            .n28256(n28256), .n28255(n28255), .n28254(n28254), .n47523(n47523), 
            .n28253(n28253), .n28252(n28252), .n28251(n28251), .n28250(n28250), 
            .n28249(n28249), .n28248(n28248), .timer({timer}), .VCC_net(VCC_net), 
            .n28247(n28247), .n28246(n28246), .n28245(n28245), .n28244(n28244), 
            .n28243(n28243), .n28242(n28242), .n28241(n28241), .n28240(n28240), 
            .n28239(n28239), .n28238(n28238), .n28237(n28237), .n28236(n28236), 
            .n28235(n28235), .n28234(n28234), .n28233(n28233), .n28232(n28232), 
            .n12(n12_adj_5053), .NEOPXL_c(NEOPXL_c), .n28163(n28163), 
            .LED_c(LED_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n37972), .I0(n2133), 
            .I1(VCC_net), .CO(n37973));
    SB_LUT4 i15120_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_5013), 
            .I3(n26633), .O(n28179));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15120_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33778_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48731));
    defparam i33778_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n640), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_78_8 (.CI(n37197), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n37198));
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n640), 
            .I1(GND_net), .CO(n37972));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n38470), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n37171), .O(n679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n37196), .O(encoder1_position_scaled_23__N_58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n38221), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n38221), .I0(n2321), 
            .I1(VCC_net), .CO(n38222));
    SB_DFF dir_62 (.Q(INHC_c), .C(CLK_c), .D(duty[23]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n38470), .I0(n3207), 
            .I1(VCC_net), .CO(n38471));
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n49129), .I1(n2016), 
            .I2(VCC_net), .I3(n37971), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_84_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[0]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15121_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_5013), 
            .I3(n26628), .O(n28180));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15121_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15523_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n23943), .I3(GND_net), .O(n28582));   // verilog/coms.v(127[12] 300[6])
    defparam i15523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15524_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n23943), .I3(GND_net), .O(n28583));   // verilog/coms.v(127[12] 300[6])
    defparam i15524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15525_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n23943), .I3(GND_net), .O(n28584));   // verilog/coms.v(127[12] 300[6])
    defparam i15525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15526_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n23943), .I3(GND_net), .O(n28585));   // verilog/coms.v(127[12] 300[6])
    defparam i15526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15527_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n23943), .I3(GND_net), .O(n28586));   // verilog/coms.v(127[12] 300[6])
    defparam i15527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33797_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48750));
    defparam i33797_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15528_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n23943), .I3(GND_net), .O(n28587));   // verilog/coms.v(127[12] 300[6])
    defparam i15528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15529_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n23943), .I3(GND_net), .O(n28588));   // verilog/coms.v(127[12] 300[6])
    defparam i15529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15530_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n23943), .I3(GND_net), .O(n28589));   // verilog/coms.v(127[12] 300[6])
    defparam i15530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15531_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n23943), .I3(GND_net), .O(n28590));   // verilog/coms.v(127[12] 300[6])
    defparam i15531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[1]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15532_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n23943), .I3(GND_net), .O(n28591));   // verilog/coms.v(127[12] 300[6])
    defparam i15532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15533_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n23943), .I3(GND_net), .O(n28592));   // verilog/coms.v(127[12] 300[6])
    defparam i15533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15534_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n23943), .I3(GND_net), .O(n28593));   // verilog/coms.v(127[12] 300[6])
    defparam i15534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15535_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n23943), .I3(GND_net), .O(n28594));   // verilog/coms.v(127[12] 300[6])
    defparam i15535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15536_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n23943), .I3(GND_net), .O(n28595));   // verilog/coms.v(127[12] 300[6])
    defparam i15536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_scaled_23__I_2_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_231));   // verilog/TinyFPGA_B.v(223[33:52])
    defparam encoder1_position_scaled_23__I_2_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i33816_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48769));
    defparam i33816_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15189_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n2380), .I3(GND_net), .O(n28248));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15537_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n23943), .I3(GND_net), .O(n28596));   // verilog/coms.v(127[12] 300[6])
    defparam i15537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15538_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n23943), .I3(GND_net), .O(n28597));   // verilog/coms.v(127[12] 300[6])
    defparam i15538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15539_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n23943), .I3(GND_net), .O(n28598));   // verilog/coms.v(127[12] 300[6])
    defparam i15539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15540_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n23943), .I3(GND_net), .O(n28599));   // verilog/coms.v(127[12] 300[6])
    defparam i15540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15541_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n23943), .I3(GND_net), .O(n28600));   // verilog/coms.v(127[12] 300[6])
    defparam i15541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15190_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n2380), .I3(GND_net), .O(n28249));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15191_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n2380), .I3(GND_net), .O(n28250));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15542_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n23943), .I3(GND_net), .O(n28601));   // verilog/coms.v(127[12] 300[6])
    defparam i15542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15543_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n23943), .I3(GND_net), .O(n28602));   // verilog/coms.v(127[12] 300[6])
    defparam i15543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15544_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n23943), .I3(GND_net), .O(n28603));   // verilog/coms.v(127[12] 300[6])
    defparam i15544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15545_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n23943), .I3(GND_net), .O(n28604));   // verilog/coms.v(127[12] 300[6])
    defparam i15545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15546_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n23943), .I3(GND_net), .O(n28605));   // verilog/coms.v(127[12] 300[6])
    defparam i15546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15192_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n2380), .I3(GND_net), .O(n28251));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15547_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n23943), .I3(GND_net), .O(n28606));   // verilog/coms.v(127[12] 300[6])
    defparam i15547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15548_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n23943), .I3(GND_net), .O(n28607));   // verilog/coms.v(127[12] 300[6])
    defparam i15548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15549_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n23943), .I3(GND_net), .O(n28608));   // verilog/coms.v(127[12] 300[6])
    defparam i15549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15550_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n23943), .I3(GND_net), .O(n28609));   // verilog/coms.v(127[12] 300[6])
    defparam i15550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15193_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n2380), .I3(GND_net), .O(n28252));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15194_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n2380), .I3(GND_net), .O(n28253));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15551_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n23943), .I3(GND_net), .O(n28610));   // verilog/coms.v(127[12] 300[6])
    defparam i15551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15552_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n23943), .I3(GND_net), .O(n28611));   // verilog/coms.v(127[12] 300[6])
    defparam i15552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15553_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n23943), .I3(GND_net), .O(n28612));   // verilog/coms.v(127[12] 300[6])
    defparam i15553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15554_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n23943), .I3(GND_net), .O(n28613));   // verilog/coms.v(127[12] 300[6])
    defparam i15554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15555_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n23943), .I3(GND_net), .O(n28614));   // verilog/coms.v(127[12] 300[6])
    defparam i15555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[2]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15556_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n23943), .I3(GND_net), .O(n28615));   // verilog/coms.v(127[12] 300[6])
    defparam i15556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15557_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n23943), .I3(GND_net), .O(n28616));   // verilog/coms.v(127[12] 300[6])
    defparam i15557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15558_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n23943), .I3(GND_net), .O(n28617));   // verilog/coms.v(127[12] 300[6])
    defparam i15558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15559_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n23943), .I3(GND_net), .O(n28618));   // verilog/coms.v(127[12] 300[6])
    defparam i15559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15560_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n23943), .I3(GND_net), .O(n28619));   // verilog/coms.v(127[12] 300[6])
    defparam i15560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15561_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n23943), .I3(GND_net), .O(n28620));   // verilog/coms.v(127[12] 300[6])
    defparam i15561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15562_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n23943), .I3(GND_net), .O(n28621));   // verilog/coms.v(127[12] 300[6])
    defparam i15562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15563_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n23943), .I3(GND_net), .O(n28622));   // verilog/coms.v(127[12] 300[6])
    defparam i15563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15564_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n23943), .I3(GND_net), .O(n28623));   // verilog/coms.v(127[12] 300[6])
    defparam i15564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15565_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n23943), .I3(GND_net), .O(n28624));   // verilog/coms.v(127[12] 300[6])
    defparam i15565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33834_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48787));
    defparam i33834_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15195_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n2380), .I3(GND_net), .O(n28254));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15566_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n23943), .I3(GND_net), .O(n28625));   // verilog/coms.v(127[12] 300[6])
    defparam i15566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15567_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n23943), .I3(GND_net), .O(n28626));   // verilog/coms.v(127[12] 300[6])
    defparam i15567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15568_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n23943), .I3(GND_net), .O(n28627));   // verilog/coms.v(127[12] 300[6])
    defparam i15568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15569_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n23943), .I3(GND_net), .O(n28628));   // verilog/coms.v(127[12] 300[6])
    defparam i15569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15570_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n23943), .I3(GND_net), .O(n28629));   // verilog/coms.v(127[12] 300[6])
    defparam i15570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15196_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n2380), .I3(GND_net), .O(n28255));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15197_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n2380), .I3(GND_net), .O(n28256));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n37970), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15571_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n23943), .I3(GND_net), .O(n28630));   // verilog/coms.v(127[12] 300[6])
    defparam i15571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15572_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n23943), .I3(GND_net), .O(n28631));   // verilog/coms.v(127[12] 300[6])
    defparam i15572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15573_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n23943), .I3(GND_net), .O(n28632));   // verilog/coms.v(127[12] 300[6])
    defparam i15573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15574_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n23943), .I3(GND_net), .O(n28633));   // verilog/coms.v(127[12] 300[6])
    defparam i15574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15575_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n23943), .I3(GND_net), .O(n28634));   // verilog/coms.v(127[12] 300[6])
    defparam i15575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15576_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n23943), .I3(GND_net), .O(n28635));   // verilog/coms.v(127[12] 300[6])
    defparam i15576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15577_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n23943), .I3(GND_net), .O(n28636));   // verilog/coms.v(127[12] 300[6])
    defparam i15577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15578_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n23943), .I3(GND_net), .O(n28637));   // verilog/coms.v(127[12] 300[6])
    defparam i15578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15579_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n23943), .I3(GND_net), .O(n28638));   // verilog/coms.v(127[12] 300[6])
    defparam i15579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15580_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n23943), .I3(GND_net), .O(n28639));   // verilog/coms.v(127[12] 300[6])
    defparam i15580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15581_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n23943), .I3(GND_net), .O(n28640));   // verilog/coms.v(127[12] 300[6])
    defparam i15581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15582_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n23943), .I3(GND_net), .O(n28641));   // verilog/coms.v(127[12] 300[6])
    defparam i15582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15583_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n23943), .I3(GND_net), .O(n28642));   // verilog/coms.v(127[12] 300[6])
    defparam i15583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15584_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n23943), .I3(GND_net), .O(n28643));   // verilog/coms.v(127[12] 300[6])
    defparam i15584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15585_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n23943), .I3(GND_net), .O(n28644));   // verilog/coms.v(127[12] 300[6])
    defparam i15585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15586_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n23943), .I3(GND_net), .O(n28645));   // verilog/coms.v(127[12] 300[6])
    defparam i15586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15587_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n23943), 
            .I3(GND_net), .O(n28646));   // verilog/coms.v(127[12] 300[6])
    defparam i15587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15588_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n23943), 
            .I3(GND_net), .O(n28647));   // verilog/coms.v(127[12] 300[6])
    defparam i15588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15198_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n2380), .I3(GND_net), .O(n28257));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15589_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n23943), 
            .I3(GND_net), .O(n28648));   // verilog/coms.v(127[12] 300[6])
    defparam i15589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15199_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n2380), .I3(GND_net), .O(n28258));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15200_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n2380), .I3(GND_net), .O(n28259));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15201_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n2380), .I3(GND_net), .O(n28260));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15590_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n23943), 
            .I3(GND_net), .O(n28649));   // verilog/coms.v(127[12] 300[6])
    defparam i15590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15591_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n23943), 
            .I3(GND_net), .O(n28650));   // verilog/coms.v(127[12] 300[6])
    defparam i15591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15592_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n23943), 
            .I3(GND_net), .O(n28651));   // verilog/coms.v(127[12] 300[6])
    defparam i15592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15593_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n23943), 
            .I3(GND_net), .O(n28652));   // verilog/coms.v(127[12] 300[6])
    defparam i15593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15202_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n2380), .I3(GND_net), .O(n28261));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34083_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49036));
    defparam i34083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15594_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n23943), 
            .I3(GND_net), .O(n28653));   // verilog/coms.v(127[12] 300[6])
    defparam i15594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15595_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n27752), 
            .I3(GND_net), .O(n28654));   // verilog/coms.v(127[12] 300[6])
    defparam i15595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15596_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n27752), 
            .I3(GND_net), .O(n28655));   // verilog/coms.v(127[12] 300[6])
    defparam i15596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15597_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n27752), 
            .I3(GND_net), .O(n28656));   // verilog/coms.v(127[12] 300[6])
    defparam i15597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15598_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n27752), 
            .I3(GND_net), .O(n28657));   // verilog/coms.v(127[12] 300[6])
    defparam i15598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15599_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n27752), 
            .I3(GND_net), .O(n28658));   // verilog/coms.v(127[12] 300[6])
    defparam i15599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15600_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n27752), 
            .I3(GND_net), .O(n28659));   // verilog/coms.v(127[12] 300[6])
    defparam i15600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15601_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n27752), 
            .I3(GND_net), .O(n28660));   // verilog/coms.v(127[12] 300[6])
    defparam i15601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15602_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n27752), 
            .I3(GND_net), .O(n28661));   // verilog/coms.v(127[12] 300[6])
    defparam i15602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15603_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n27752), 
            .I3(GND_net), .O(n28662));   // verilog/coms.v(127[12] 300[6])
    defparam i15603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15604_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n27752), 
            .I3(GND_net), .O(n28663));   // verilog/coms.v(127[12] 300[6])
    defparam i15604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15605_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n27752), 
            .I3(GND_net), .O(n28664));   // verilog/coms.v(127[12] 300[6])
    defparam i15605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15606_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n27752), 
            .I3(GND_net), .O(n28665));   // verilog/coms.v(127[12] 300[6])
    defparam i15606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15607_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n27752), 
            .I3(GND_net), .O(n28666));   // verilog/coms.v(127[12] 300[6])
    defparam i15607_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n37970), .I0(n2017), 
            .I1(VCC_net), .CO(n37971));
    SB_LUT4 i15608_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n27752), 
            .I3(GND_net), .O(n28667));   // verilog/coms.v(127[12] 300[6])
    defparam i15608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15609_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n27752), 
            .I3(GND_net), .O(n28668));   // verilog/coms.v(127[12] 300[6])
    defparam i15609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[3]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15610_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n27752), 
            .I3(GND_net), .O(n28669));   // verilog/coms.v(127[12] 300[6])
    defparam i15610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n651));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15611_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n27752), 
            .I3(GND_net), .O(n28670));   // verilog/coms.v(127[12] 300[6])
    defparam i15611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15203_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n2380), .I3(GND_net), .O(n28262));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15612_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n27752), 
            .I3(GND_net), .O(n28671));   // verilog/coms.v(127[12] 300[6])
    defparam i15612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n37969), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15613_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n27752), 
            .I3(GND_net), .O(n28672));   // verilog/coms.v(127[12] 300[6])
    defparam i15613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n650), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15614_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n27752), 
            .I3(GND_net), .O(n28673));   // verilog/coms.v(127[12] 300[6])
    defparam i15614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15615_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n27752), 
            .I3(GND_net), .O(n28674));   // verilog/coms.v(127[12] 300[6])
    defparam i15615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15616_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n27752), 
            .I3(GND_net), .O(n28675));   // verilog/coms.v(127[12] 300[6])
    defparam i15616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15617_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n27752), 
            .I3(GND_net), .O(n28676));   // verilog/coms.v(127[12] 300[6])
    defparam i15617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15618_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n27752), 
            .I3(GND_net), .O(n28677));   // verilog/coms.v(127[12] 300[6])
    defparam i15618_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n5722), 
            .D(n659), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15619_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n27752), 
            .I3(GND_net), .O(n28678));   // verilog/coms.v(127[12] 300[6])
    defparam i15619_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n5722), 
            .D(n660), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n5722), 
            .D(n661), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n5722), 
            .D(n662), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i33951_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48904));
    defparam i33951_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15620_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n27752), 
            .I3(GND_net), .O(n28679));   // verilog/coms.v(127[12] 300[6])
    defparam i15620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15621_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n27752), 
            .I3(GND_net), .O(n28680));   // verilog/coms.v(127[12] 300[6])
    defparam i15621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15622_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n27752), 
            .I3(GND_net), .O(n28681));   // verilog/coms.v(127[12] 300[6])
    defparam i15622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15623_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n27752), 
            .I3(GND_net), .O(n28682));   // verilog/coms.v(127[12] 300[6])
    defparam i15623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15204_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n27752), .I3(GND_net), .O(n28263));   // verilog/coms.v(127[12] 300[6])
    defparam i15204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15624_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n27752), 
            .I3(GND_net), .O(n28683));   // verilog/coms.v(127[12] 300[6])
    defparam i15624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15625_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28684));   // verilog/coms.v(127[12] 300[6])
    defparam i15625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15626_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28685));   // verilog/coms.v(127[12] 300[6])
    defparam i15626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15627_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28686));   // verilog/coms.v(127[12] 300[6])
    defparam i15627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15628_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28687));   // verilog/coms.v(127[12] 300[6])
    defparam i15628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15629_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28688));   // verilog/coms.v(127[12] 300[6])
    defparam i15629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15630_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28689));   // verilog/coms.v(127[12] 300[6])
    defparam i15630_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n5722), 
            .D(n663), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n5722), 
            .D(n664), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n5722), 
            .D(n665), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n37969), .I0(n2018), 
            .I1(VCC_net), .CO(n37970));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n37968), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n37968), .I0(n2019), 
            .I1(VCC_net), .CO(n37969));
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n37967), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n37967), .I0(n2020), 
            .I1(VCC_net), .CO(n37968));
    SB_LUT4 i15631_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28690));   // verilog/coms.v(127[12] 300[6])
    defparam i15631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15632_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28691));   // verilog/coms.v(127[12] 300[6])
    defparam i15632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15633_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28692));   // verilog/coms.v(127[12] 300[6])
    defparam i15633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15634_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28693));   // verilog/coms.v(127[12] 300[6])
    defparam i15634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15205_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n27752), .I3(GND_net), .O(n28264));   // verilog/coms.v(127[12] 300[6])
    defparam i15205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15635_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28694));   // verilog/coms.v(127[12] 300[6])
    defparam i15635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15636_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28695));   // verilog/coms.v(127[12] 300[6])
    defparam i15636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15206_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n27752), .I3(GND_net), .O(n28265));   // verilog/coms.v(127[12] 300[6])
    defparam i15206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15637_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28696));   // verilog/coms.v(127[12] 300[6])
    defparam i15637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15638_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28697));   // verilog/coms.v(127[12] 300[6])
    defparam i15638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15639_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28698));   // verilog/coms.v(127[12] 300[6])
    defparam i15639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15207_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n27752), .I3(GND_net), .O(n28266));   // verilog/coms.v(127[12] 300[6])
    defparam i15207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28130_4_lut (.I0(n7_adj_5098), .I1(state_adj_5154[0]), .I2(n6_adj_5032), 
            .I3(state_adj_5170[0]), .O(n43002));
    defparam i28130_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i15208_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n27752), .I3(GND_net), .O(n28267));   // verilog/coms.v(127[12] 300[6])
    defparam i15208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15209_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n27752), .I3(GND_net), .O(n28268));   // verilog/coms.v(127[12] 300[6])
    defparam i15209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33855_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48808));
    defparam i33855_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15210_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n27752), .I3(GND_net), .O(n28269));   // verilog/coms.v(127[12] 300[6])
    defparam i15210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15211_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n27752), .I3(GND_net), .O(n28270));   // verilog/coms.v(127[12] 300[6])
    defparam i15211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15212_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n27752), .I3(GND_net), .O(n28271));   // verilog/coms.v(127[12] 300[6])
    defparam i15212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33878_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48831));
    defparam i33878_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut (.I0(state_adj_5154[1]), .I1(read), .I2(n43073), 
            .I3(GND_net), .O(n12_adj_5056));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n34306), .I1(n12_adj_5056), .I2(state_adj_5154[0]), 
            .I3(n43073), .O(n41845));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut.LUT_INIT = 16'h88a8;
    SB_LUT4 i15641_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28700));   // verilog/coms.v(127[12] 300[6])
    defparam i15641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15642_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28701));   // verilog/coms.v(127[12] 300[6])
    defparam i15642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15643_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28702));   // verilog/coms.v(127[12] 300[6])
    defparam i15643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15644_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28703));   // verilog/coms.v(127[12] 300[6])
    defparam i15644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15645_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28704));   // verilog/coms.v(127[12] 300[6])
    defparam i15645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15646_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28705));   // verilog/coms.v(127[12] 300[6])
    defparam i15646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15647_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28706));   // verilog/coms.v(127[12] 300[6])
    defparam i15647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15648_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28707));   // verilog/coms.v(127[12] 300[6])
    defparam i15648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15649_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28708));   // verilog/coms.v(127[12] 300[6])
    defparam i15649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15650_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28709));   // verilog/coms.v(127[12] 300[6])
    defparam i15650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15651_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28710));   // verilog/coms.v(127[12] 300[6])
    defparam i15651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15652_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28711));   // verilog/coms.v(127[12] 300[6])
    defparam i15652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15653_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28712));   // verilog/coms.v(127[12] 300[6])
    defparam i15653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15654_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28713));   // verilog/coms.v(127[12] 300[6])
    defparam i15654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n37966), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n37966), .I0(n2021), 
            .I1(VCC_net), .CO(n37967));
    SB_LUT4 i15655_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28714));   // verilog/coms.v(127[12] 300[6])
    defparam i15655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n37965), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n37965), .I0(n2022), 
            .I1(VCC_net), .CO(n37966));
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n37964), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n38469), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n38355), .I0(n2811), 
            .I1(VCC_net), .CO(n38356));
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n37964), .I0(n2023), 
            .I1(VCC_net), .CO(n37965));
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n37963), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33324_3_lut (.I0(n1727), .I1(n1794), .I2(n1752), .I3(GND_net), 
            .O(n1826));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15656_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28715));   // verilog/coms.v(127[12] 300[6])
    defparam i15656_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n38469), .I0(n3208), 
            .I1(VCC_net), .CO(n38470));
    SB_LUT4 i15657_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n27752), .I3(GND_net), .O(n28716));   // verilog/coms.v(127[12] 300[6])
    defparam i15657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15658_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n27752), .I3(GND_net), .O(n28717));   // verilog/coms.v(127[12] 300[6])
    defparam i15658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15659_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n27752), .I3(GND_net), .O(n28718));   // verilog/coms.v(127[12] 300[6])
    defparam i15659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15660_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n27752), .I3(GND_net), .O(n28719));   // verilog/coms.v(127[12] 300[6])
    defparam i15660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15661_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n27752), .I3(GND_net), .O(n28720));   // verilog/coms.v(127[12] 300[6])
    defparam i15661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15662_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n27752), .I3(GND_net), .O(n28721));   // verilog/coms.v(127[12] 300[6])
    defparam i15662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15663_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n27752), .I3(GND_net), .O(n28722));   // verilog/coms.v(127[12] 300[6])
    defparam i15663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15664_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n27752), .I3(GND_net), .O(n28723));   // verilog/coms.v(127[12] 300[6])
    defparam i15664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15665_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n27752), .I3(GND_net), .O(n28724));   // verilog/coms.v(127[12] 300[6])
    defparam i15665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15666_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n27752), .I3(GND_net), .O(n28725));   // verilog/coms.v(127[12] 300[6])
    defparam i15666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15667_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n27752), .I3(GND_net), .O(n28726));   // verilog/coms.v(127[12] 300[6])
    defparam i15667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15668_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n27752), .I3(GND_net), .O(n28727));   // verilog/coms.v(127[12] 300[6])
    defparam i15668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15669_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n27752), .I3(GND_net), .O(n28728));   // verilog/coms.v(127[12] 300[6])
    defparam i15669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15670_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n27752), .I3(GND_net), .O(n28729));   // verilog/coms.v(127[12] 300[6])
    defparam i15670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15671_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n27752), .I3(GND_net), .O(n28730));   // verilog/coms.v(127[12] 300[6])
    defparam i15671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[4]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15672_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n27752), .I3(GND_net), .O(n28731));   // verilog/coms.v(127[12] 300[6])
    defparam i15672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28083_3_lut (.I0(n6_adj_5018), .I1(n6541), .I2(n42948), .I3(GND_net), 
            .O(n42955));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28084_3_lut (.I0(encoder0_position[27]), .I1(n42955), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15673_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n27752), .I3(GND_net), .O(n28732));   // verilog/coms.v(127[12] 300[6])
    defparam i15673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15674_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n27752), .I3(GND_net), .O(n28733));   // verilog/coms.v(127[12] 300[6])
    defparam i15674_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n37963), .I0(n2024), 
            .I1(VCC_net), .CO(n37964));
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15675_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n27752), .I3(GND_net), .O(n28734));   // verilog/coms.v(127[12] 300[6])
    defparam i15675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15676_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n27752), .I3(GND_net), .O(n28735));   // verilog/coms.v(127[12] 300[6])
    defparam i15676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[5]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15677_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n27752), .I3(GND_net), .O(n28736));   // verilog/coms.v(127[12] 300[6])
    defparam i15677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15678_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n27752), .I3(GND_net), .O(n28737));   // verilog/coms.v(127[12] 300[6])
    defparam i15678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15679_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n27752), .I3(GND_net), .O(n28738));   // verilog/coms.v(127[12] 300[6])
    defparam i15679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[6]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28079_3_lut (.I0(n4_adj_5020), .I1(n6539), .I2(n42948), .I3(GND_net), 
            .O(n42951));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15682_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n44870), .I3(GND_net), 
            .O(n28741));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15682_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15683_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n44870), .I3(GND_net), 
            .O(n28742));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28080_3_lut (.I0(encoder0_position[29]), .I1(n42951), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15684_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n44870), .I3(GND_net), 
            .O(n28743));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15684_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15685_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n44870), .I3(GND_net), 
            .O(n28744));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15685_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15686_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n44870), .I3(GND_net), 
            .O(n28745));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15686_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15687_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n44870), .I3(GND_net), 
            .O(n28746));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15687_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15688_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n44870), .I3(GND_net), 
            .O(n28747));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15688_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1669 (.I0(n5_adj_5017), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n1419), .I3(read_N_321), .O(n25_adj_4951));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i1_4_lut_adj_1669.LUT_INIT = 16'h7350;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31665_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46544));
    defparam i31665_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33918_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n5855), .I2(n46544), 
            .I3(n25_adj_4951), .O(n17_adj_4952));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i33918_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15213_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n27752), .I3(GND_net), .O(n28272));   // verilog/coms.v(127[12] 300[6])
    defparam i15213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33906_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48859));
    defparam i33906_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15214_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n27752), .I3(GND_net), .O(n28273));   // verilog/coms.v(127[12] 300[6])
    defparam i15214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[7]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15122_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n33696), 
            .I3(n26633), .O(n28181));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15122_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15123_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n33696), 
            .I3(n26628), .O(n28182));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15123_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15215_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n27752), .I3(GND_net), .O(n28274));   // verilog/coms.v(127[12] 300[6])
    defparam i15215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15216_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n27752), .I3(GND_net), .O(n28275));   // verilog/coms.v(127[12] 300[6])
    defparam i15216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_84_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[8]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_5018), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n625));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5_adj_5019), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n516));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_5020), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3_adj_5021), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n622));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4093_2_lut (.I0(n2_adj_5022), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4093_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5088));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5087));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5086));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5085));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n37962), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n38220), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n38354), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n38220), .I0(n2322), 
            .I1(VCC_net), .CO(n38221));
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n37962), .I0(n2025), 
            .I1(VCC_net), .CO(n37963));
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n37961), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n37961), .I0(n2026), 
            .I1(VCC_net), .CO(n37962));
    SB_LUT4 mux_84_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[9]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n38219), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n38219), .I0(n2323), 
            .I1(VCC_net), .CO(n38220));
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n38078), .I0(n2227), 
            .I1(VCC_net), .CO(n38079));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5084));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5083));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5082));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5081));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5080));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5079));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5078));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n37960), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n37960), .I0(n2027), 
            .I1(VCC_net), .CO(n37961));
    SB_CARRY add_78_7 (.CI(n37196), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n37197));
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n38468), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5077));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n37959), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n38468), .I0(n3209), 
            .I1(VCC_net), .CO(n38469));
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n38467), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5076));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5075));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5074));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5073));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(146[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5072));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5071));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5070));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n37959), .I0(n2028), 
            .I1(VCC_net), .CO(n37960));
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n37958), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5069));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5068));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5067));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5066));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5065));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5064));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n38218), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5063));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5062));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5061));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5060));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5059));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5058));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5057));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_84_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[10]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_84_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[11]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n38218), .I0(n2324), 
            .I1(VCC_net), .CO(n38219));
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n38077), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15124_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28183));   // verilog/coms.v(127[12] 300[6])
    defparam i15124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15125_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n27752), 
            .I3(GND_net), .O(n28184));   // verilog/coms.v(127[12] 300[6])
    defparam i15125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15126_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n27752), 
            .I3(GND_net), .O(n28185));   // verilog/coms.v(127[12] 300[6])
    defparam i15126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15127_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n27753), .I3(GND_net), .O(n28186));   // verilog/coms.v(127[12] 300[6])
    defparam i15127_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n38354), .I0(n2812), 
            .I1(VCC_net), .CO(n38355));
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n38353), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n38467), .I0(n3210), 
            .I1(VCC_net), .CO(n38468));
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n38077), .I0(n2228), 
            .I1(VCC_net), .CO(n38078));
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n37958), .I0(n2029), 
            .I1(GND_net), .CO(n37959));
    SB_LUT4 i15128_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n42229), 
            .I3(GND_net), .O(n28187));   // verilog/coms.v(127[12] 300[6])
    defparam i15128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34278_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49231));
    defparam i34278_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33326_3_lut (.I0(n1827), .I1(n1894), .I2(n1851), .I3(GND_net), 
            .O(n1926));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15129_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n27752), .I3(GND_net), .O(n28188));   // verilog/coms.v(127[12] 300[6])
    defparam i15129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n37957), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n37957), .I0(n2030), 
            .I1(GND_net), .CO(n37958));
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n5722), 
            .D(n666), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n38076), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n38466), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n38353), .I0(n2813), 
            .I1(VCC_net), .CO(n38354));
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n38217), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n38217), .I0(n2325), 
            .I1(VCC_net), .CO(n38218));
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n38076), .I0(n2229), 
            .I1(GND_net), .CO(n38077));
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n38075), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n38075), .I0(n2230), 
            .I1(GND_net), .CO(n38076));
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n38074), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n38074), .I0(n2231), 
            .I1(VCC_net), .CO(n38075));
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n37956), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n37956), .I0(n2031), 
            .I1(VCC_net), .CO(n37957));
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n38466), .I0(n3211), 
            .I1(VCC_net), .CO(n38467));
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n38465), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n38352), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n38465), .I0(n3212), 
            .I1(VCC_net), .CO(n38466));
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n38464), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n38352), .I0(n2814), 
            .I1(VCC_net), .CO(n38353));
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n38351), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n38351), .I0(n2815), 
            .I1(VCC_net), .CO(n38352));
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n38350), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n38216), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n38216), .I0(n2326), 
            .I1(VCC_net), .CO(n38217));
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n38215), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n38215), .I0(n2327), 
            .I1(VCC_net), .CO(n38216));
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n38214), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n37955), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n37955), .I0(n2032), 
            .I1(GND_net), .CO(n37956));
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n37954), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n37954), .I0(n2033), 
            .I1(VCC_net), .CO(n37955));
    SB_LUT4 encoder0_position_31__I_0_i1245_3_lut (.I0(n46594), .I1(n1628), 
            .I2(n48039), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34206_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n45256), 
            .O(n2148));
    defparam i34206_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n639), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n5722), 
            .D(n667), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n639), 
            .I1(GND_net), .CO(n37954));
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n49096), .I1(n1917), 
            .I2(VCC_net), .I3(n37953), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n38350), .I0(n2816), 
            .I1(VCC_net), .CO(n38351));
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n38073), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n38349), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n38464), .I0(n3213), 
            .I1(VCC_net), .CO(n38465));
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n38463), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n37952), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n38463), .I0(n3214), 
            .I1(VCC_net), .CO(n38464));
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n37952), .I0(n1918), 
            .I1(VCC_net), .CO(n37953));
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n38462), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n38214), .I0(n2328), 
            .I1(VCC_net), .CO(n38215));
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n38462), .I0(n3215), 
            .I1(VCC_net), .CO(n38463));
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n38349), .I0(n2817), 
            .I1(VCC_net), .CO(n38350));
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n37951), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n37951), .I0(n1919), 
            .I1(VCC_net), .CO(n37952));
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n37950), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n37950), .I0(n1920), 
            .I1(VCC_net), .CO(n37951));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n37949), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n38461), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n38461), .I0(n3216), 
            .I1(VCC_net), .CO(n38462));
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n38460), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n38348), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n38460), .I0(n3217), 
            .I1(VCC_net), .CO(n38461));
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n38213), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n38213), .I0(n2329), 
            .I1(GND_net), .CO(n38214));
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n38459), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n38459), .I0(n3218), 
            .I1(VCC_net), .CO(n38460));
    SB_LUT4 add_78_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n37195), .O(encoder1_position_scaled_23__N_58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n38073), .I0(n2232), 
            .I1(GND_net), .CO(n38074));
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n38458), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n38072), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n38072), .I0(n2233), 
            .I1(VCC_net), .CO(n38073));
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n641), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n38212), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n37949), .I0(n1921), 
            .I1(VCC_net), .CO(n37950));
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n641), 
            .I1(GND_net), .CO(n38072));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n37948), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n37948), .I0(n1922), 
            .I1(VCC_net), .CO(n37949));
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n38348), .I0(n2818), 
            .I1(VCC_net), .CO(n38349));
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n38347), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n37947), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n37947), .I0(n1923), 
            .I1(VCC_net), .CO(n37948));
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n37946), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n37946), .I0(n1924), 
            .I1(VCC_net), .CO(n37947));
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n37945), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15130_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n27752), .I3(GND_net), .O(n28189));   // verilog/coms.v(127[12] 300[6])
    defparam i15130_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n38458), .I0(n3219), 
            .I1(VCC_net), .CO(n38459));
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n38347), .I0(n2819), 
            .I1(VCC_net), .CO(n38348));
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n38457), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n38457), .I0(n3220), 
            .I1(VCC_net), .CO(n38458));
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n38212), .I0(n2330), 
            .I1(GND_net), .CO(n38213));
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n38346), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n38456), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n37945), .I0(n1925), 
            .I1(VCC_net), .CO(n37946));
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n37944), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_78_6 (.CI(n37195), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n37196));
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n37944), .I0(n1926), 
            .I1(VCC_net), .CO(n37945));
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n37943), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n38211), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n37943), .I0(n1927), 
            .I1(VCC_net), .CO(n37944));
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n38456), .I0(n3221), 
            .I1(VCC_net), .CO(n38457));
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n38211), .I0(n2331), 
            .I1(VCC_net), .CO(n38212));
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n38455), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n38210), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n37194), .O(encoder1_position_scaled_23__N_58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n38346), .I0(n2820), 
            .I1(VCC_net), .CO(n38347));
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n5722), 
            .D(n685), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n37942), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n5722), 
            .D(n668), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n37942), .I0(n1928), 
            .I1(VCC_net), .CO(n37943));
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n37941), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n5722), 
            .D(n686), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n37941), .I0(n1929), 
            .I1(GND_net), .CO(n37942));
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n38345), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_22__N_11[0]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n38210), .I0(n2332), 
            .I1(GND_net), .CO(n38211));
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n38209), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n38345), .I0(n2821), 
            .I1(VCC_net), .CO(n38346));
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n38344), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n38455), .I0(n3222), 
            .I1(VCC_net), .CO(n38456));
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n38344), .I0(n2822), 
            .I1(VCC_net), .CO(n38345));
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n38209), .I0(n2333), 
            .I1(VCC_net), .CO(n38210));
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n642), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n642), 
            .I1(GND_net), .CO(n38209));
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n38454), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n38343), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n38343), .I0(n2823), 
            .I1(VCC_net), .CO(n38344));
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n37940), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n38454), .I0(n3223), 
            .I1(VCC_net), .CO(n38455));
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n38342), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(enable_slow_N_4090), .I1(data_ready), 
            .I2(state_adj_5154[1]), .I3(state_adj_5154[0]), .O(n41955));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'hccd0;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n37940), .I0(n1930), 
            .I1(GND_net), .CO(n37941));
    SB_CARRY add_78_5 (.CI(n37194), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n37195));
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n37939), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n37939), .I0(n1931), 
            .I1(VCC_net), .CO(n37940));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n38453), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n37938), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n37938), .I0(n1932), 
            .I1(GND_net), .CO(n37939));
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n38342), .I0(n2824), 
            .I1(VCC_net), .CO(n38343));
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n38453), .I0(n3224), 
            .I1(VCC_net), .CO(n38454));
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n37937), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n38341), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n38341), .I0(n2825), 
            .I1(VCC_net), .CO(n38342));
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n37937), .I0(n1933), 
            .I1(VCC_net), .CO(n37938));
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n38452), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n638), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n5722), 
            .D(n669), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n638), 
            .I1(GND_net), .CO(n37937));
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n5722), 
            .D(n670), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n38340), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n38452), .I0(n3225), 
            .I1(VCC_net), .CO(n38453));
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n48859), .I1(n1818), 
            .I2(VCC_net), .I3(n37936), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n37935), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n38340), .I0(n2826), 
            .I1(VCC_net), .CO(n38341));
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n38451), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n37935), .I0(n1819), 
            .I1(VCC_net), .CO(n37936));
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n37934), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n37934), .I0(n1820), 
            .I1(VCC_net), .CO(n37935));
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n37933), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n37933), .I0(n1821), 
            .I1(VCC_net), .CO(n37934));
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n38339), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n38339), .I0(n2827), 
            .I1(VCC_net), .CO(n38340));
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n37932), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n37193), .O(encoder1_position_scaled_23__N_58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n37932), .I0(n1822), 
            .I1(VCC_net), .CO(n37933));
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n38451), .I0(n3226), 
            .I1(VCC_net), .CO(n38452));
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n38450), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n37931), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n37931), .I0(n1823), 
            .I1(VCC_net), .CO(n37932));
    SB_CARRY add_78_4 (.CI(n37193), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n37194));
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n37930), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n37930), .I0(n1824), 
            .I1(VCC_net), .CO(n37931));
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n37929), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n37929), .I0(n1825), 
            .I1(VCC_net), .CO(n37930));
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n38338), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n37928), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n37928), .I0(n1826), 
            .I1(VCC_net), .CO(n37929));
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n37927), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n38450), .I0(n3227), 
            .I1(VCC_net), .CO(n38451));
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n37927), .I0(n1827), 
            .I1(VCC_net), .CO(n37928));
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n37926), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n37926), .I0(n1828), 
            .I1(VCC_net), .CO(n37927));
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n38338), .I0(n2828), 
            .I1(VCC_net), .CO(n38339));
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n38449), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n38449), .I0(n3228), 
            .I1(VCC_net), .CO(n38450));
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n38448), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n37925), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n38337), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n37925), .I0(n1829), 
            .I1(GND_net), .CO(n37926));
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n37924), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n37924), .I0(n1830), 
            .I1(GND_net), .CO(n37925));
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n37923), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n38337), .I0(n2829), 
            .I1(GND_net), .CO(n38338));
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n37923), .I0(n1831), 
            .I1(VCC_net), .CO(n37924));
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n38336), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n37922), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n37922), .I0(n1832), 
            .I1(GND_net), .CO(n37923));
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n37921), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n37921), .I0(n1833), 
            .I1(VCC_net), .CO(n37922));
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n637), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n637), 
            .I1(GND_net), .CO(n37921));
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n48831), .I1(n1719), 
            .I2(VCC_net), .I3(n37920), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n37919), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n37919), .I0(n1720), 
            .I1(VCC_net), .CO(n37920));
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n37918), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n37918), .I0(n1721), 
            .I1(VCC_net), .CO(n37919));
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n37917), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n37917), .I0(n1722), 
            .I1(VCC_net), .CO(n37918));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n37916), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n38336), .I0(n2830), 
            .I1(GND_net), .CO(n38337));
    SB_LUT4 mux_84_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[12]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i34015_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48968));
    defparam i34015_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15217_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n27752), .I3(GND_net), .O(n28276));   // verilog/coms.v(127[12] 300[6])
    defparam i15217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n37916), .I0(n1723), 
            .I1(VCC_net), .CO(n37917));
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n37915), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n37915), .I0(n1724), 
            .I1(VCC_net), .CO(n37916));
    SB_LUT4 i15218_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n27752), .I3(GND_net), .O(n28277));   // verilog/coms.v(127[12] 300[6])
    defparam i15218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n5722), 
            .D(n687), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i34143_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49096));
    defparam i34143_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n37914), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n5722), 
            .D(n688), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n37914), .I0(n1725), 
            .I1(VCC_net), .CO(n37915));
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n37913), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n37913), .I0(n1726), 
            .I1(VCC_net), .CO(n37914));
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n37912), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n37912), .I0(n1727), 
            .I1(VCC_net), .CO(n37913));
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n37911), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n37911), .I0(n1728), 
            .I1(VCC_net), .CO(n37912));
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n37910), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n37910), .I0(n1729), 
            .I1(GND_net), .CO(n37911));
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n37909), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n37909), .I0(n1730), 
            .I1(GND_net), .CO(n37910));
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n37908), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n37908), .I0(n1731), 
            .I1(VCC_net), .CO(n37909));
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n37907), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n37907), .I0(n1732), 
            .I1(GND_net), .CO(n37908));
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n37906), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n37906), .I0(n1733), 
            .I1(VCC_net), .CO(n37907));
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n636), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n636), 
            .I1(GND_net), .CO(n37906));
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n48808), .I1(n1620), 
            .I2(VCC_net), .I3(n37905), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n37904), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n37904), .I0(n1621), 
            .I1(VCC_net), .CO(n37905));
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n37903), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n37903), .I0(n1622), 
            .I1(VCC_net), .CO(n37904));
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n37902), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n37902), .I0(n1623), 
            .I1(VCC_net), .CO(n37903));
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n37901), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n37901), .I0(n1624), 
            .I1(VCC_net), .CO(n37902));
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n37900), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17_adj_4993), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n636));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n37900), .I0(n1625), 
            .I1(VCC_net), .CO(n37901));
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n636), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n37899), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n37899), .I0(n1626), 
            .I1(VCC_net), .CO(n37900));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n37898), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n37898), .I0(n1627), 
            .I1(VCC_net), .CO(n37899));
    SB_LUT4 i34200_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49153));
    defparam i34200_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15219_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n27752), .I3(GND_net), .O(n28278));   // verilog/coms.v(127[12] 300[6])
    defparam i15219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15220_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n27752), .I3(GND_net), .O(n28279));   // verilog/coms.v(127[12] 300[6])
    defparam i15220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15221_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n27752), .I3(GND_net), .O(n28280));   // verilog/coms.v(127[12] 300[6])
    defparam i15221_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n38448), .I0(n3229), 
            .I1(GND_net), .CO(n38449));
    SB_LUT4 i15222_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n27752), .I3(GND_net), .O(n28281));   // verilog/coms.v(127[12] 300[6])
    defparam i15222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n38447), .O(n47538)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_84_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[13]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n37897), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n38335), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n38335), .I0(n2831), 
            .I1(VCC_net), .CO(n38336));
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n37897), .I0(n1628), 
            .I1(VCC_net), .CO(n37898));
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n38447), .I0(n3230), 
            .I1(GND_net), .CO(n38448));
    SB_LUT4 encoder0_position_31__I_0_i1313_3_lut (.I0(n46588), .I1(n1728), 
            .I2(n48037), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15223_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n27752), .I3(GND_net), .O(n28282));   // verilog/coms.v(127[12] 300[6])
    defparam i15223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_84_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[14]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n5722), 
            .D(n671), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n37896), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n37896), .I0(n1629), 
            .I1(GND_net), .CO(n37897));
    SB_LUT4 LessThan_700_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5037));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i9_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n5722), 
            .D(n672), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 LessThan_700_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5039));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n37895), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28085_3_lut (.I0(n7_adj_5003), .I1(n6542), .I2(n42948), .I3(GND_net), 
            .O(n42957));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28086_3_lut (.I0(encoder0_position[26]), .I1(n42957), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n38446), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n37895), .I0(n1630), 
            .I1(GND_net), .CO(n37896));
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_700_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5043));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n37894), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n37894), .I0(n1631), 
            .I1(VCC_net), .CO(n37895));
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n38334), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n38446), .I0(n3231), 
            .I1(VCC_net), .CO(n38447));
    SB_LUT4 LessThan_700_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5048));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n37893), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n37893), .I0(n1632), 
            .I1(GND_net), .CO(n37894));
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n5722), 
            .D(n689), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 LessThan_700_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5042));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n37892), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n37892), .I0(n1633), 
            .I1(VCC_net), .CO(n37893));
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n635), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_700_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5041));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_84_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[15]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n38334), .I0(n2832), 
            .I1(GND_net), .CO(n38335));
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n38333), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n38333), .I0(n2833), 
            .I1(VCC_net), .CO(n38334));
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n635), 
            .I1(GND_net), .CO(n37892));
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n38445), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n647), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15224_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n27752), .I3(GND_net), .O(n28283));   // verilog/coms.v(127[12] 300[6])
    defparam i15224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n647), 
            .I1(GND_net), .CO(n38333));
    SB_LUT4 LessThan_700_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5035));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(n48904), .I1(n2709), 
            .I2(VCC_net), .I3(n38332), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n38445), .I0(n3232), 
            .I1(GND_net), .CO(n38446));
    SB_LUT4 LessThan_700_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5045));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_78_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n37192), .O(encoder1_position_scaled_23__N_58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_700_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5046));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n38331), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_700_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5044));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n38331), .I0(n2710), 
            .I1(VCC_net), .CO(n38332));
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n38444), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n38444), .I0(n3233), 
            .I1(VCC_net), .CO(n38445));
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n38330), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n651), 
            .I2(GND_net), .I3(n38443), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_700_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5049));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15132_4_lut (.I0(rw), .I1(state_adj_5154[0]), .I2(state_adj_5154[1]), 
            .I3(n4227), .O(n28191));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15132_4_lut.LUT_INIT = 16'hacaa;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n38443), .I0(n651), 
            .I1(GND_net), .CO(n38444));
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n38330), .I0(n2711), 
            .I1(VCC_net), .CO(n38331));
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n38329), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_700_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5051));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(delay_counter[12]), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4978));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_700_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5052));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_4978), .I2(delay_counter[10]), 
            .I3(n26517), .O(n43755));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1671 (.I0(n43755), .I1(n26511), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n44222));
    defparam i2_4_lut_adj_1671.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_4982));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n38329), .I0(n2712), 
            .I1(VCC_net), .CO(n38330));
    SB_LUT4 i2_4_lut_adj_1672 (.I0(delay_counter[22]), .I1(n44222), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_4983));
    defparam i2_4_lut_adj_1672.LUT_INIT = 16'ha8a0;
    SB_CARRY add_78_3 (.CI(n37192), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n37193));
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n652), 
            .I1(VCC_net), .CO(n38443));
    SB_LUT4 i20766_4_lut (.I0(n7_adj_4983), .I1(delay_counter[31]), .I2(n26514), 
            .I3(n8_adj_4982), .O(n777));   // verilog/TinyFPGA_B.v(280[14:38])
    defparam i20766_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_4974));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n38328), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n49036), .I1(n3105), 
            .I2(VCC_net), .I3(n38442), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n38328), .I0(n2713), 
            .I1(VCC_net), .CO(n38329));
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12_adj_4974), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n26514));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n38441), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n38441), .I0(n3106), 
            .I1(VCC_net), .CO(n38442));
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n38440), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n5722), 
            .D(n690), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n5722), 
            .D(n673), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n37978), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15133_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5161[1]), .I2(n19247), 
            .I3(n4_adj_5007), .O(n28192));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15133_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_4976));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15135_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_3987[0]), 
            .I3(enable_slow_N_4090), .O(n28194));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15135_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i6_4_lut_adj_1673 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_4975));
    defparam i6_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n37978), .I0(n2127), 
            .I1(VCC_net), .CO(n37979));
    SB_LUT4 i2_3_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n44870));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 mux_84_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[17]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15136_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n44870), .I3(GND_net), 
            .O(n28195));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n37977), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4975), .I1(delay_counter[2]), .I2(n14_adj_4976), 
            .I3(delay_counter[6]), .O(n26517));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1674 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n26511));
    defparam i2_3_lut_adj_1674.LUT_INIT = 16'hfefe;
    SB_LUT4 i3764_4_lut (.I0(n26517), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5031));
    defparam i3764_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1675 (.I0(n24_adj_5031), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n44044));
    defparam i2_4_lut_adj_1675.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1676 (.I0(n44044), .I1(delay_counter[18]), .I2(n26511), 
            .I3(GND_net), .O(n44198));
    defparam i2_3_lut_adj_1676.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1677 (.I0(n5_adj_5008), .I1(n3_adj_5021), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n45386));
    defparam i1_3_lut_adj_1677.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1678 (.I0(delay_counter[23]), .I1(n44198), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5006));
    defparam i2_4_lut_adj_1678.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut (.I0(n7_adj_5006), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n26514), .O(n62));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20763_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_321));   // verilog/TinyFPGA_B.v(265[12:35])
    defparam i20763_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4950));   // verilog/TinyFPGA_B.v(278[12:17])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1679 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_4949));   // verilog/TinyFPGA_B.v(278[12:17])
    defparam i6_4_lut_adj_1679.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(ID[3]), .I1(n14_adj_4949), .I2(n10_adj_4950), 
            .I3(ID[6]), .O(n26487));   // verilog/TinyFPGA_B.v(278[12:17])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 \ID_READOUT_FSM.state_2__I_0_i5_2_lut  (.I0(\ID_READOUT_FSM.state [0]), 
            .I1(\ID_READOUT_FSM.state [1]), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_5017));   // verilog/TinyFPGA_B.v(277[7:11])
    defparam \ID_READOUT_FSM.state_2__I_0_i5_2_lut .LUT_INIT = 16'hbbbb;
    SB_LUT4 i15074_4_lut (.I0(n5722), .I1(n777), .I2(n47518), .I3(n26488), 
            .O(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15074_4_lut.LUT_INIT = 16'ha088;
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n37977), .I0(n2128), 
            .I1(VCC_net), .CO(n37978));
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut (.I0(n2_adj_5022), .I1(n6537), 
            .I2(n45386), .I3(encoder0_position[31]), .O(n828));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 i4_4_lut_adj_1680 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4977));   // verilog/TinyFPGA_B.v(169[5:22])
    defparam i4_4_lut_adj_1680.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1681 (.I0(control_mode[6]), .I1(n10_adj_4977), 
            .I2(control_mode[2]), .I3(GND_net), .O(n26607));   // verilog/TinyFPGA_B.v(169[5:22])
    defparam i5_3_lut_adj_1681.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n48787), .I1(n1521), 
            .I2(VCC_net), .I3(n37881), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n38327), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1682 (.I0(n26489), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4947));   // verilog/TinyFPGA_B.v(170[5:22])
    defparam i1_2_lut_adj_1682.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n37880), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n37880), .I0(n1522), 
            .I1(VCC_net), .CO(n37881));
    SB_LUT4 i2_3_lut_adj_1683 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n26607), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(169[5:22])
    defparam i2_3_lut_adj_1683.LUT_INIT = 16'hfdfd;
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n37879), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_84_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[16]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n37879), .I0(n1523), 
            .I1(VCC_net), .CO(n37880));
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n37878), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_84_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[18]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n37976), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n37878), .I0(n1524), 
            .I1(VCC_net), .CO(n37879));
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n37877), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n37877), .I0(n1525), 
            .I1(VCC_net), .CO(n37878));
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n37976), .I0(n2129), 
            .I1(GND_net), .CO(n37977));
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n38440), .I0(n3107), 
            .I1(VCC_net), .CO(n38441));
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n37876), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n37975), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n37975), .I0(n2130), 
            .I1(GND_net), .CO(n37976));
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n37876), .I0(n1526), 
            .I1(VCC_net), .CO(n37877));
    SB_LUT4 mux_84_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[19]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n38439), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n37875), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n38327), .I0(n2714), 
            .I1(VCC_net), .CO(n38328));
    SB_CARRY add_29_13 (.CI(n37171), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n37172));
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n37875), .I0(n1527), 
            .I1(VCC_net), .CO(n37876));
    SB_LUT4 i34087_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49040));
    defparam i34087_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_84_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[20]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n37874), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n38326), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n38439), .I0(n3108), 
            .I1(VCC_net), .CO(n38440));
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n37874), .I0(n1528), 
            .I1(VCC_net), .CO(n37875));
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n37873), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n38326), .I0(n2715), 
            .I1(VCC_net), .CO(n38327));
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n38438), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n37873), .I0(n1529), 
            .I1(GND_net), .CO(n37874));
    SB_LUT4 mux_84_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[21]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n37872), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n37872), .I0(n1530), 
            .I1(GND_net), .CO(n37873));
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n37871), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n37973), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n37871), .I0(n1531), 
            .I1(VCC_net), .CO(n37872));
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n38325), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n37870), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n37870), .I0(n1532), 
            .I1(GND_net), .CO(n37871));
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n37869), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n37869), .I0(n1533), 
            .I1(VCC_net), .CO(n37870));
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n634), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n634), 
            .I1(GND_net), .CO(n37869));
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(n48769), .I1(n1422), 
            .I2(VCC_net), .I3(n37868), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n37867), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n37867), .I0(n1423), 
            .I1(VCC_net), .CO(n37868));
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n37866), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n37866), .I0(n1424), 
            .I1(VCC_net), .CO(n37867));
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n37865), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n37865), .I0(n1425), 
            .I1(VCC_net), .CO(n37866));
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n37864), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n37864), .I0(n1426), 
            .I1(VCC_net), .CO(n37865));
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n37863), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_231), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n37863), .I0(n1427), 
            .I1(VCC_net), .CO(n37864));
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n37862), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n37862), .I0(n1428), 
            .I1(VCC_net), .CO(n37863));
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n38438), .I0(n3109), 
            .I1(VCC_net), .CO(n38439));
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n38437), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n37861), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n38325), .I0(n2716), 
            .I1(VCC_net), .CO(n38326));
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n38324), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34121_1_lut (.I0(n34679), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49074));
    defparam i34121_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5094));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n37861), .I0(n1429), 
            .I1(GND_net), .CO(n37862));
    SB_LUT4 encoder0_position_31__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5096));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_78_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n37197), .O(encoder1_position_scaled_23__N_58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n37860), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n37860), .I0(n1430), 
            .I1(GND_net), .CO(n37861));
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n37859), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n37859), .I0(n1431), 
            .I1(VCC_net), .CO(n37860));
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n37858), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n37858), .I0(n1432), 
            .I1(GND_net), .CO(n37859));
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n37857), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n37857), .I0(n1433), 
            .I1(VCC_net), .CO(n37858));
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n633), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5092));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n633), 
            .I1(GND_net), .CO(n37857));
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n48750), .I1(n1323), 
            .I2(VCC_net), .I3(n37856), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n37855), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n37855), .I0(n1324), 
            .I1(VCC_net), .CO(n37856));
    SB_LUT4 encoder0_position_31__I_0_i2195_3_lut (.I0(n3224), .I1(n3291), 
            .I2(n3237), .I3(GND_net), .O(n23_adj_5095));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n37854), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n37854), .I0(n1325), 
            .I1(VCC_net), .CO(n37855));
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n37853), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n3221), .I1(n23_adj_5095), .I2(n3288), 
            .I3(n3237), .O(n45106));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n37853), .I0(n1326), 
            .I1(VCC_net), .CO(n37854));
    SB_CARRY add_78_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_231), 
            .CO(n37192));
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n38437), .I0(n3110), 
            .I1(VCC_net), .CO(n38438));
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n38324), .I0(n2717), 
            .I1(VCC_net), .CO(n38325));
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n37852), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n37191), .O(n659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n37852), .I0(n1327), 
            .I1(VCC_net), .CO(n37853));
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n37851), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21270_4_lut (.I0(n652), .I1(n651), .I2(n3301), .I3(n3237), 
            .O(n34313));
    defparam i21270_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i21433_4_lut (.I0(n34313), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n34481));
    defparam i21433_4_lut.LUT_INIT = 16'h88a0;
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n37851), .I0(n1328), 
            .I1(VCC_net), .CO(n37852));
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n38436), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n37850), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n37850), .I0(n1329), 
            .I1(GND_net), .CO(n37851));
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n38323), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n37849), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n37190), .O(n660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5091));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n37974), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5093));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n37849), .I0(n1330), 
            .I1(GND_net), .CO(n37850));
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n37848), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n37848), .I0(n1331), 
            .I1(VCC_net), .CO(n37849));
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n3220), .I1(n21_adj_5094), .I2(n3287), 
            .I3(n3237), .O(n45100));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n37847), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n37847), .I0(n1332), 
            .I1(GND_net), .CO(n37848));
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n37846), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n37846), .I0(n1333), 
            .I1(VCC_net), .CO(n37847));
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n632), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n38436), .I0(n3111), 
            .I1(VCC_net), .CO(n38437));
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n38323), .I0(n2718), 
            .I1(VCC_net), .CO(n38324));
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n632), 
            .I1(GND_net), .CO(n37846));
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n38435), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n48731), .I1(n1224), 
            .I2(VCC_net), .I3(n37845), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n3219), .I1(n27_adj_5096), .I2(n3286), 
            .I3(n3237), .O(n45110));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n37844), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n37844), .I0(n1225), 
            .I1(VCC_net), .CO(n37845));
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n37843), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_32 (.CI(n37190), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n37191));
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n37843), .I0(n1226), 
            .I1(VCC_net), .CO(n37844));
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n37842), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n37842), .I0(n1227), 
            .I1(VCC_net), .CO(n37843));
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n37841), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n37841), .I0(n1228), 
            .I1(VCC_net), .CO(n37842));
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n37840), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n38435), .I0(n3112), 
            .I1(VCC_net), .CO(n38436));
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n37840), .I0(n1229), 
            .I1(GND_net), .CO(n37841));
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n37839), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n38322), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n38434), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n38434), .I0(n3113), 
            .I1(VCC_net), .CO(n38435));
    SB_LUT4 encoder0_position_31__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5090));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n37839), .I0(n1230), 
            .I1(GND_net), .CO(n37840));
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n3223), .I1(n17_adj_5092), .I2(n3290), 
            .I3(n3237), .O(n45104));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n37838), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n37838), .I0(n1231), 
            .I1(VCC_net), .CO(n37839));
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n37837), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n5722), 
            .D(n674), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n37837), .I0(n1232), 
            .I1(GND_net), .CO(n37838));
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n37836), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n37836), .I0(n1233), 
            .I1(VCC_net), .CO(n37837));
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n38433), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n631), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n631), 
            .I1(GND_net), .CO(n37836));
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n37974), .I0(n2131), 
            .I1(VCC_net), .CO(n37975));
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n38322), .I0(n2719), 
            .I1(VCC_net), .CO(n38323));
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n38321), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n38321), .I0(n2720), 
            .I1(VCC_net), .CO(n38322));
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n38320), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(n45106), .I1(n3217), .I2(n3284), .I3(n3237), 
            .O(n45112));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'heefa;
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n38320), .I0(n2721), 
            .I1(VCC_net), .CO(n38321));
    SB_LUT4 i1_4_lut_adj_1689 (.I0(n13_adj_5090), .I1(n45110), .I2(n45100), 
            .I3(n19_adj_5093), .O(n45118));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n38319), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n38319), .I0(n2722), 
            .I1(VCC_net), .CO(n38320));
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n38433), .I0(n3114), 
            .I1(VCC_net), .CO(n38434));
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n38318), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n38318), .I0(n2723), 
            .I1(VCC_net), .CO(n38319));
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n38317), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n38317), .I0(n2724), 
            .I1(VCC_net), .CO(n38318));
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n38432), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n38432), .I0(n3115), 
            .I1(VCC_net), .CO(n38433));
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n38431), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n38316), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n3218), .I1(n15_adj_5091), .I2(n3285), 
            .I3(n3237), .O(n45102));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n38431), .I0(n3116), 
            .I1(VCC_net), .CO(n38432));
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n38430), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n38316), .I0(n2725), 
            .I1(VCC_net), .CO(n38317));
    SB_LUT4 add_78_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n37198), .O(encoder1_position_scaled_23__N_58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n38430), .I0(n3117), 
            .I1(VCC_net), .CO(n38431));
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n38429), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n38429), .I0(n3118), 
            .I1(VCC_net), .CO(n38430));
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n38315), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n38428), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n48717), .I1(n1125), 
            .I2(VCC_net), .I3(n37825), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n45102), .I1(n45118), .I2(n45112), 
            .I3(n45104), .O(n45122));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n45122), .I1(n3216), .I2(n3283), .I3(n3237), 
            .O(n45124));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'heefa;
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n38428), .I0(n3119), 
            .I1(VCC_net), .CO(n38429));
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n38427), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n37824), .O(n1193_adj_5029)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n37824), .I0(n1126), 
            .I1(VCC_net), .CO(n37825));
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n37823), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n38315), .I0(n2726), 
            .I1(VCC_net), .CO(n38316));
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n38314), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n38314), .I0(n2727), 
            .I1(VCC_net), .CO(n38315));
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n37823), .I0(n1127), 
            .I1(VCC_net), .CO(n37824));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n38313), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n38427), .I0(n3120), 
            .I1(VCC_net), .CO(n38428));
    SB_LUT4 i33609_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48562));
    defparam i33609_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n37822), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n37822), .I0(n1128), 
            .I1(VCC_net), .CO(n37823));
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n38426), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n37821), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n37821), .I0(n1129), 
            .I1(GND_net), .CO(n37822));
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n37820), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n38313), .I0(n2728), 
            .I1(VCC_net), .CO(n38314));
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n37820), .I0(n1130), 
            .I1(GND_net), .CO(n37821));
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n47538), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5016));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n37819), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(n3215), .I1(n45124), .I2(n3282), .I3(n3237), 
            .O(n45126));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n37819), .I0(n1131), 
            .I1(VCC_net), .CO(n37820));
    SB_LUT4 encoder0_position_31__I_0_i2185_3_lut (.I0(n3214), .I1(n3281), 
            .I2(n3237), .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n37818), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n38312), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21533_4_lut (.I0(n34481), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n34583));
    defparam i21533_4_lut.LUT_INIT = 16'heefa;
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n37818), .I0(n1132), 
            .I1(GND_net), .CO(n37819));
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n34583), .I1(n43), .I2(n45126), .I3(n5_adj_5016), 
            .O(n45130));
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'hfefc;
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n37817), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n3213), .I1(n45130), .I2(n3280), .I3(n3237), 
            .O(n45132));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n37817), .I0(n1133), 
            .I1(VCC_net), .CO(n37818));
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n630), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n38312), .I0(n2729), 
            .I1(GND_net), .CO(n38313));
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n630), 
            .I1(GND_net), .CO(n37817));
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n37816), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n37815), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n37815), .I0(n1027), 
            .I1(VCC_net), .CO(n37816));
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n38426), .I0(n3121), 
            .I1(VCC_net), .CO(n38427));
    SB_LUT4 i1_4_lut_adj_1696 (.I0(n3212), .I1(n45132), .I2(n3279), .I3(n3237), 
            .O(n45134));
    defparam i1_4_lut_adj_1696.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n38425), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n37170), .O(n680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n37814), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(n3211), .I1(n45134), .I2(n3278), .I3(n3237), 
            .O(n45136));
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n37814), .I0(n1028), 
            .I1(VCC_net), .CO(n37815));
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n37813), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n37813), .I0(n1029), 
            .I1(GND_net), .CO(n37814));
    SB_LUT4 add_29_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n37189), .O(n661)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n38425), .I0(n3122), 
            .I1(VCC_net), .CO(n38426));
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n3210), .I1(n45136), .I2(n3277), .I3(n3237), 
            .O(n45138));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n38424), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n3209), .I1(n45138), .I2(n3276), .I3(n3237), 
            .O(n45140));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'heefc;
    SB_CARRY add_29_5 (.CI(n37163), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n37164));
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n37812), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n37812), .I0(n1030), 
            .I1(GND_net), .CO(n37813));
    SB_CARRY add_29_12 (.CI(n37170), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n37171));
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n38311), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n38311), .I0(n2730), 
            .I1(GND_net), .CO(n38312));
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n38310), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n38310), .I0(n2731), 
            .I1(VCC_net), .CO(n38311));
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n37811), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n37811), .I0(n1031), 
            .I1(VCC_net), .CO(n37812));
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n37810), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n37169), .O(n681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n38309), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n3208), .I1(n45140), .I2(n3275), .I3(n3237), 
            .O(n45142));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n38424), .I0(n3123), 
            .I1(VCC_net), .CO(n38425));
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n3207), .I1(n45142), .I2(n3274), .I3(n3237), 
            .O(n45144));
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n38309), .I0(n2732), 
            .I1(GND_net), .CO(n38310));
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n37810), .I0(n1032), 
            .I1(GND_net), .CO(n37811));
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n37809), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n37809), .I0(n1033), 
            .I1(VCC_net), .CO(n37810));
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n629), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n38308), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n38423), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n38423), .I0(n3124), 
            .I1(VCC_net), .CO(n38424));
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n629), 
            .I1(GND_net), .CO(n37809));
    SB_LUT4 i34124_4_lut (.I0(n61), .I1(n46486), .I2(n59), .I3(n45144), 
            .O(n34679));
    defparam i34124_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i33983_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48936));
    defparam i33983_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_84_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[22]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_84_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15), .I3(n15_adj_4947), .O(motor_state_23__N_106[23]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_84_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n37808), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n38422), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n37807), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n38422), .I0(n3125), 
            .I1(VCC_net), .CO(n38423));
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n37807), .I0(n928), 
            .I1(VCC_net), .CO(n37808));
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n38308), .I0(n2733), 
            .I1(VCC_net), .CO(n38309));
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n646), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n37806), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n37806), .I0(n929), 
            .I1(GND_net), .CO(n37807));
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n3222), .I1(n3225), .I2(n3220), .I3(n3227), 
            .O(n45620));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n37805), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n3224), .I1(n3226), .I2(n3228), .I3(n3221), 
            .O(n45618));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n45618), .I1(n45620), .I2(n3219), .I3(n3223), 
            .O(n45624));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i21537_4_lut (.I0(n651), .I1(n3231), .I2(n3232), .I3(n3233), 
            .O(n34587));
    defparam i21537_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n37805), .I0(n930), 
            .I1(GND_net), .CO(n37806));
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n3216), .I1(n3217), .I2(n45624), .I3(n3218), 
            .O(n45630));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n45630), .I1(n3229), .I2(n34587), .I3(n3230), 
            .O(n45632));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'heaaa;
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n37804), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(n3213), .I1(n3214), .I2(n3215), .I3(n45632), 
            .O(n45638));
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n45638), 
            .O(n45644));
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n37804), .I0(n931), 
            .I1(VCC_net), .CO(n37805));
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n37803), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n37803), .I0(n932), 
            .I1(GND_net), .CO(n37804));
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n646), 
            .I1(GND_net), .CO(n38308));
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n37802), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n38421), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_78_11 (.CI(n37200), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n37201));
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n45644), 
            .O(n45650));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_CARRY add_29_31 (.CI(n37189), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n37190));
    SB_LUT4 i34120_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n45650), 
            .O(n3237));
    defparam i34120_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i34049_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49002));
    defparam i34049_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n37802), .I0(n933), 
            .I1(VCC_net), .CO(n37803));
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n628), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n38421), .I0(n3126), 
            .I1(VCC_net), .CO(n38422));
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n628), 
            .I1(GND_net), .CO(n37802));
    SB_LUT4 i33665_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48618));
    defparam i33665_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34254_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49207));
    defparam i34254_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34228_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49181));
    defparam i34228_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n38420), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n38420), .I0(n3127), 
            .I1(VCC_net), .CO(n38421));
    SB_LUT4 i34176_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49129));
    defparam i34176_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n38419), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33764_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48717));
    defparam i33764_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33743_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48696));
    defparam i33743_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n38419), .I0(n3128), 
            .I1(VCC_net), .CO(n38420));
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n38418), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n38418), .I0(n3129), 
            .I1(GND_net), .CO(n38419));
    SB_LUT4 i32822_2_lut (.I0(n49422), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47614));
    defparam i32822_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31707_4_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n46660));
    defparam i31707_4_lut.LUT_INIT = 16'hc00a;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n41391));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i15225_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n27752), .I3(GND_net), .O(n28284));   // verilog/coms.v(127[12] 300[6])
    defparam i15225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15226_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n27752), .I3(GND_net), .O(n28285));   // verilog/coms.v(127[12] 300[6])
    defparam i15226_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 mux_82_i18_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[17]), 
            .I3(encoder0_position_scaled[17]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_82_i19_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[18]), 
            .I3(encoder0_position_scaled[18]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15227_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n27752), .I3(GND_net), .O(n28286));   // verilog/coms.v(127[12] 300[6])
    defparam i15227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_29_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n37188), .O(n662)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n38417), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15228_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n27752), .I3(GND_net), .O(n28287));   // verilog/coms.v(127[12] 300[6])
    defparam i15228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2041_3_lut (.I0(n3006), .I1(n3073), 
            .I2(n3039), .I3(GND_net), .O(n3105));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n38417), .I0(n3130), 
            .I1(GND_net), .CO(n38418));
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n38416), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n38416), .I0(n3131), 
            .I1(VCC_net), .CO(n38417));
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n38415), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n38415), .I0(n3132), 
            .I1(GND_net), .CO(n38416));
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n38414), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_11 (.CI(n37169), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n37170));
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n38414), .I0(n3133), 
            .I1(VCC_net), .CO(n38415));
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n650), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n650), 
            .I1(GND_net), .CO(n38414));
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(GND_net), .I1(n3006), 
            .I2(VCC_net), .I3(n38413), .O(n3073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n38412), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(n48618), .I1(n2610), 
            .I2(VCC_net), .I3(n38298), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n38297), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n38297), .I0(n2611), 
            .I1(VCC_net), .CO(n38298));
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n38412), .I0(n3007), 
            .I1(VCC_net), .CO(n38413));
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n38296), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n38411), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n38411), .I0(n3008), 
            .I1(VCC_net), .CO(n38412));
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n38410), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n38296), .I0(n2612), 
            .I1(VCC_net), .CO(n38297));
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n38295), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n38295), .I0(n2613), 
            .I1(VCC_net), .CO(n38296));
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n38410), .I0(n3009), 
            .I1(VCC_net), .CO(n38411));
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n38409), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n38294), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n649), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n38294), .I0(n2614), 
            .I1(VCC_net), .CO(n38295));
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n38293), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n650));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n38409), .I0(n3010), 
            .I1(VCC_net), .CO(n38410));
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n38293), .I0(n2615), 
            .I1(VCC_net), .CO(n38294));
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n38292), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n38408), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n38292), .I0(n2616), 
            .I1(VCC_net), .CO(n38293));
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n38408), .I0(n3011), 
            .I1(VCC_net), .CO(n38409));
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n38407), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n38407), .I0(n3012), 
            .I1(VCC_net), .CO(n38408));
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n38291), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n38291), .I0(n2617), 
            .I1(VCC_net), .CO(n38292));
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n38290), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n38406), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n38290), .I0(n2618), 
            .I1(VCC_net), .CO(n38291));
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n38406), .I0(n3013), 
            .I1(VCC_net), .CO(n38407));
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n38289), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n38289), .I0(n2619), 
            .I1(VCC_net), .CO(n38290));
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n37162), .O(n688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n38405), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n38405), .I0(n3014), 
            .I1(VCC_net), .CO(n38406));
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n38288), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i20_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[19]), 
            .I3(encoder0_position_scaled[19]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_82_i21_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[20]), 
            .I3(encoder0_position_scaled[20]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n38404), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n38288), .I0(n2620), 
            .I1(VCC_net), .CO(n38289));
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n38287), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_82[23]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 encoder0_position_31__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i22_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[21]), 
            .I3(encoder0_position_scaled[21]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_82[22]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n38287), .I0(n2621), 
            .I1(VCC_net), .CO(n38288));
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n38404), .I0(n3015), 
            .I1(VCC_net), .CO(n38405));
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n38286), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n38403), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n38286), .I0(n2622), 
            .I1(VCC_net), .CO(n38287));
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n38403), .I0(n3016), 
            .I1(VCC_net), .CO(n38404));
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n38285), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_82[21]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_82[20]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_82[19]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_82[18]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_82[17]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_82[16]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_82[15]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_82[14]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_82[13]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_82[12]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_82[11]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_82[10]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_82[9]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_82[8]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_82[7]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_82[6]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_82[5]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_82[4]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_82[3]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_82[2]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_82[1]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[23]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[22]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[21]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[20]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[19]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[18]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[17]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[16]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[15]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[14]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[13]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[12]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[11]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[10]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[9]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[8]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[7]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[6]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[5]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[4]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[3]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[2]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[1]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i23_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[22]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n5722), 
            .D(n675), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n38402), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n38402), .I0(n3017), 
            .I1(VCC_net), .CO(n38403));
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n38285), .I0(n2623), 
            .I1(VCC_net), .CO(n38286));
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n38401), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n38401), .I0(n3018), 
            .I1(VCC_net), .CO(n38402));
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n647), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i24_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[23]), 
            .I3(encoder0_position_scaled[23]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7_adj_5003), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n626));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_adj_1710 (.I0(pwm_counter[27]), .I1(pwm_counter[28]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5055));
    defparam i2_2_lut_adj_1710.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1711 (.I0(pwm_counter[23]), .I1(pwm_counter[29]), 
            .I2(pwm_counter[25]), .I3(pwm_counter[26]), .O(n14_adj_5054));
    defparam i6_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1712 (.I0(pwm_counter[30]), .I1(n14_adj_5054), 
            .I2(n10_adj_5055), .I3(pwm_counter[24]), .O(n26497));
    defparam i7_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n646), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n647));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33239_3_lut (.I0(n2624), .I1(n2691), .I2(n2643), .I3(GND_net), 
            .O(n2723));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33240_3_lut (.I0(n2723), .I1(n2790), .I2(n2742), .I3(GND_net), 
            .O(n2822));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33245_3_lut (.I0(n2628), .I1(n2695), .I2(n2643), .I3(GND_net), 
            .O(n2727));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n4_adj_5020), .I1(n5_adj_5019), .I2(n626), 
            .I3(n6_adj_5018), .O(n5_adj_5008));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'heeea;
    SB_LUT4 i33246_3_lut (.I0(n2727), .I1(n2794), .I2(n2742), .I3(GND_net), 
            .O(n2826));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n645), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_DFF read_66 (.Q(read), .C(CLK_c), .D(n44886));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n646));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n38400), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n38400), .I0(n3019), 
            .I1(VCC_net), .CO(n38401));
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n38399), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n38399), .I0(n3020), 
            .I1(VCC_net), .CO(n38400));
    SB_LUT4 i33235_3_lut (.I0(n2522), .I1(n2589), .I2(n2544), .I3(GND_net), 
            .O(n2621));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33235_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33236_3_lut (.I0(n2621), .I1(n2688), .I2(n2643), .I3(GND_net), 
            .O(n2720));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33236_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i1_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[23]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n38284), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n38284), .I0(n2624), 
            .I1(VCC_net), .CO(n38285));
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n38283), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n38398), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33237_3_lut (.I0(n2523), .I1(n2590), .I2(n2544), .I3(GND_net), 
            .O(n2622));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33238_3_lut (.I0(n2622), .I1(n2689), .I2(n2643), .I3(GND_net), 
            .O(n2721));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_4_lut_adj_1714 (.I0(\data_out_frame[19] [6]), .I1(n42541), 
            .I2(\data_out_frame[24] [1]), .I3(n43610), .O(n12_adj_4979));
    defparam i5_4_lut_adj_1714.LUT_INIT = 16'h9669;
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n38398), .I0(n3021), 
            .I1(VCC_net), .CO(n38399));
    SB_LUT4 mux_82_i2_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i6_4_lut_adj_1715 (.I0(n40598), .I1(n12_adj_4979), .I2(n42790), 
            .I3(\data_out_frame[24] [0]), .O(n43603));
    defparam i6_4_lut_adj_1715.LUT_INIT = 16'h9669;
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[22]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n38397), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[21]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[20]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[19]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_22__N_11[22]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_22__N_11[21]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_22__N_11[20]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_22__N_11[19]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_22__N_11[18]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_22__N_11[17]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_22__N_11[16]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_22__N_11[15]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_22__N_11[14]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_22__N_11[13]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_22__N_11[12]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_22__N_11[11]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_22__N_11[10]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_22__N_11[9]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_22__N_11[8]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_22__N_11[7]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_22__N_11[6]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_22__N_11[5]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_22__N_11[4]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_22__N_11[3]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_22__N_11[2]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_22__N_11[1]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i15233_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n27752), .I3(GND_net), .O(n28292));   // verilog/coms.v(127[12] 300[6])
    defparam i15233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n38283), .I0(n2625), 
            .I1(VCC_net), .CO(n38284));
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n38282), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n38397), .I0(n3022), 
            .I1(VCC_net), .CO(n38398));
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n38396), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n38282), .I0(n2626), 
            .I1(VCC_net), .CO(n38283));
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n38396), .I0(n3023), 
            .I1(VCC_net), .CO(n38397));
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n38395), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n38395), .I0(n3024), 
            .I1(VCC_net), .CO(n38396));
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n38281), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n38281), .I0(n2627), 
            .I1(VCC_net), .CO(n38282));
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n38280), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n38280), .I0(n2628), 
            .I1(VCC_net), .CO(n38281));
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n38279), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n38279), .I0(n2629), 
            .I1(GND_net), .CO(n38280));
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n38394), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n38278), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n38278), .I0(n2630), 
            .I1(GND_net), .CO(n38279));
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n38394), .I0(n3025), 
            .I1(VCC_net), .CO(n38395));
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n38277), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n38277), .I0(n2631), 
            .I1(VCC_net), .CO(n38278));
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n38393), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n38393), .I0(n3026), 
            .I1(VCC_net), .CO(n38394));
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n38392), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n38276), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n38276), .I0(n2632), 
            .I1(GND_net), .CO(n38277));
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n38392), .I0(n3027), 
            .I1(VCC_net), .CO(n38393));
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n38275), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n38275), .I0(n2633), 
            .I1(VCC_net), .CO(n38276));
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n38391), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n645), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n38391), .I0(n3028), 
            .I1(VCC_net), .CO(n38392));
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n38390), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n645), 
            .I1(GND_net), .CO(n38275));
    SB_LUT4 mux_82_i3_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n38390), .I0(n3029), 
            .I1(GND_net), .CO(n38391));
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n48562), .I1(n2511), 
            .I2(VCC_net), .I3(n38274), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n38273), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_30 (.CI(n37188), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n37189));
    SB_LUT4 encoder0_position_31__I_0_i1729_3_lut (.I0(n644), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n38389), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n38273), .I0(n2512), 
            .I1(VCC_net), .CO(n38274));
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n38389), .I0(n3030), 
            .I1(GND_net), .CO(n38390));
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n38272), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n38272), .I0(n2513), 
            .I1(VCC_net), .CO(n38273));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n645));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1723_rep_11_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1723_rep_11_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_4 (.CI(n37162), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n37163));
    SB_LUT4 mux_82_i4_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n38388), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i1661_3_lut (.I0(n643), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25_adj_4985), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n644));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1650_rep_23_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1650_rep_23_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i5_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1651_rep_25_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1651_rep_25_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n38388), .I0(n3031), 
            .I1(VCC_net), .CO(n38389));
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n38387), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n38271), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n38271), .I0(n2514), 
            .I1(VCC_net), .CO(n38272));
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n37710), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n38270), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n37709), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n37709), .I0(n829), 
            .I1(GND_net), .CO(n37710));
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n37708), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n37708), .I0(n830), 
            .I1(GND_net), .CO(n37709));
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n38387), .I0(n3032), 
            .I1(GND_net), .CO(n38388));
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n37707), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n37707), .I0(n831), 
            .I1(VCC_net), .CO(n37708));
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n37706), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n37706), .I0(n832), 
            .I1(GND_net), .CO(n37707));
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n37705), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n37705), .I0(n833), 
            .I1(VCC_net), .CO(n37706));
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n627), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n627), 
            .I1(GND_net), .CO(n37705));
    SB_LUT4 i1_3_lut_adj_1716 (.I0(n3_adj_5021), .I1(n2_adj_5022), .I2(n5_adj_5008), 
            .I3(GND_net), .O(n42948));
    defparam i1_3_lut_adj_1716.LUT_INIT = 16'h8080;
    SB_LUT4 i28081_3_lut (.I0(n5_adj_5019), .I1(n6540), .I2(n42948), .I3(GND_net), 
            .O(n42953));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28082_3_lut (.I0(encoder0_position[28]), .I1(n42953), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n38386), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n28195));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n5722), 
            .D(n676), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n38270), .I0(n2515), 
            .I1(VCC_net), .CO(n38271));
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n38269), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n27554), .I1(n42897), .I2(\data_out_frame[20] [0]), 
            .I3(n4_adj_5028), .O(n42541));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1718 (.I0(\data_out_frame[23] [6]), .I1(n42551), 
            .I2(GND_net), .I3(GND_net), .O(n42790));
    defparam i1_2_lut_adj_1718.LUT_INIT = 16'h9999;
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n38269), .I0(n2516), 
            .I1(VCC_net), .CO(n38270));
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1593_3_lut (.I0(n642), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24_adj_4986), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n643));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n38268), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n38386), .I0(n3033), 
            .I1(VCC_net), .CO(n38387));
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n38268), .I0(n2517), 
            .I1(VCC_net), .CO(n38269));
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33233_3_lut (.I0(n2126), .I1(n2193), .I2(n2148), .I3(GND_net), 
            .O(n2225));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33233_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33234_3_lut (.I0(n2225), .I1(n2292), .I2(n2247), .I3(GND_net), 
            .O(n2324));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33234_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n649), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n38267), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n49153), .I1(n2115), 
            .I2(VCC_net), .I3(n37990), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n37989), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n37168), .O(n682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n38267), .I0(n2518), 
            .I1(VCC_net), .CO(n38268));
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n37989), .I0(n2116), 
            .I1(VCC_net), .CO(n37990));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n37988), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_700_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5047));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_700_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1719 (.I0(n26497), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n26499));
    defparam i1_2_lut_adj_1719.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n37988), .I0(n2117), 
            .I1(VCC_net), .CO(n37989));
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n649), 
            .I1(GND_net), .CO(n38386));
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n38266), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n37987), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n37987), .I0(n2118), 
            .I1(VCC_net), .CO(n37988));
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n37986), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n48968), .I1(n2907), 
            .I2(VCC_net), .I3(n38385), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_82_i6_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n38266), .I0(n2519), 
            .I1(VCC_net), .CO(n38267));
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n37986), .I0(n2119), 
            .I1(VCC_net), .CO(n37987));
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n37985), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n38265), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n37985), .I0(n2120), 
            .I1(VCC_net), .CO(n37986));
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32738_4_lut (.I0(n27_adj_5048), .I1(n15_adj_5042), .I2(n13_adj_5041), 
            .I3(n11_adj_5039), .O(n47691));
    defparam i32738_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34396 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n49365));
    defparam byte_transmit_counter_0__bdd_4_lut_34396.LUT_INIT = 16'he4aa;
    SB_LUT4 n49365_bdd_4_lut (.I0(n49365), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n49368));
    defparam n49365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i33080_4_lut (.I0(n9_adj_5037), .I1(n7_adj_5035), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n48033));
    defparam i33080_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i33255_4_lut (.I0(n15_adj_5042), .I1(n13_adj_5041), .I2(n11_adj_5039), 
            .I3(n48033), .O(n48208));
    defparam i33255_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33253_4_lut (.I0(n21_adj_5045), .I1(n19_adj_5044), .I2(n17_adj_5043), 
            .I3(n48208), .O(n48206));
    defparam i33253_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32740_4_lut (.I0(n27_adj_5048), .I1(n25_adj_5047), .I2(n23_adj_5046), 
            .I3(n48206), .O(n47693));
    defparam i32740_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_700_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_5033));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n37984), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33029_3_lut (.I0(n2226), .I1(n2293), .I2(n2247), .I3(GND_net), 
            .O(n2325));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n38384), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n38265), .I0(n2520), 
            .I1(VCC_net), .CO(n38266));
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n37984), .I0(n2121), 
            .I1(VCC_net), .CO(n37985));
    SB_LUT4 i33231_3_lut (.I0(n2125), .I1(n2192), .I2(n2148), .I3(GND_net), 
            .O(n2224));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33231_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33232_3_lut (.I0(n2224), .I1(n2291), .I2(n2247), .I3(GND_net), 
            .O(n2323));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33232_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1525_3_lut (.I0(n641), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n37983), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n38384), .I0(n2908), 
            .I1(VCC_net), .CO(n38385));
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n38264), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n37187), .O(n663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n37983), .I0(n2122), 
            .I1(VCC_net), .CO(n37984));
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n38264), .I0(n2521), 
            .I1(VCC_net), .CO(n38265));
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n37982), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23_adj_4987), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n642));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n37982), .I0(n2123), 
            .I1(VCC_net), .CO(n37983));
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n2323), .I1(n2327), .I2(n2326), .I3(n2325), 
            .O(n45156));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_CARRY add_29_29 (.CI(n37187), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n37188));
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n37981), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1721 (.I0(n2322), .I1(n2328), .I2(n2324), .I3(GND_net), 
            .O(n45158));
    defparam i1_3_lut_adj_1721.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n38383), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n38263), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21574_4_lut (.I0(n642), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n34627));
    defparam i21574_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 add_29_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n37186), .O(n664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n37981), .I0(n2124), 
            .I1(VCC_net), .CO(n37982));
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n2320), .I1(n2321), .I2(n45158), .I3(n45156), 
            .O(n45164));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n38263), .I0(n2522), 
            .I1(VCC_net), .CO(n38264));
    SB_LUT4 i1_2_lut_adj_1723 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n45416));
    defparam i1_2_lut_adj_1723.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n45416), .I1(n2319), .I2(n45164), .I3(n34627), 
            .O(n45168));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n45168), 
            .O(n45174));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n37980), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n37980), .I0(n2125), 
            .I1(VCC_net), .CO(n37981));
    SB_LUT4 i34257_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n45174), 
            .O(n2346));
    defparam i34257_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n37979), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n37972), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_28 (.CI(n37186), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n37187));
    SB_LUT4 encoder0_position_31__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n2423), .I1(n2427), .I2(n2422), .I3(n2425), 
            .O(n45456));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n38383), .I0(n2909), 
            .I1(VCC_net), .CO(n38384));
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n2426), .I1(n45456), .I2(n2428), .I3(n2424), 
            .O(n45458));
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n38262), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n38382), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n38262), .I0(n2523), 
            .I1(VCC_net), .CO(n38263));
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n38261), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21560_4_lut (.I0(n643), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n34613));
    defparam i21560_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n38382), .I0(n2910), 
            .I1(VCC_net), .CO(n38383));
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n2419), .I1(n2420), .I2(n45458), .I3(n2421), 
            .O(n45464));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1729 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n45658));
    defparam i1_2_lut_adj_1729.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n2418), .I1(n45658), .I2(n45464), .I3(n34613), 
            .O(n45468));
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n45468), 
            .O(n45474));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_LUT4 i34284_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n45474), 
            .O(n2445));
    defparam i34284_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n38261), .I0(n2524), 
            .I1(VCC_net), .CO(n38262));
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n38260), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n38381), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n38260), .I0(n2525), 
            .I1(VCC_net), .CO(n38261));
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n38381), .I0(n2911), 
            .I1(VCC_net), .CO(n38382));
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n38259), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n37185), .O(n665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n38380), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n38259), .I0(n2526), 
            .I1(VCC_net), .CO(n38260));
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n38258), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33417_3_lut (.I0(n4_adj_5033), .I1(pwm_setpoint[13]), .I2(n27_adj_5048), 
            .I3(GND_net), .O(n48370));   // verilog/pwm.v(21[8:24])
    defparam i33417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n2524), .I1(n2525), .I2(n2526), .I3(n2527), 
            .O(n45210));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(n2523), .I1(n2521), .I2(n2528), .I3(n2522), 
            .O(n45212));
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i21459_3_lut (.I0(n644), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n34507));
    defparam i21459_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(n2519), .I1(n2520), .I2(n45212), .I3(n45210), 
            .O(n45218));
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_CARRY add_29_10 (.CI(n37168), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n37169));
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n38380), .I0(n2912), 
            .I1(VCC_net), .CO(n38381));
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n38258), .I0(n2527), 
            .I1(VCC_net), .CO(n38259));
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n38257), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n38379), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n38257), .I0(n2528), 
            .I1(VCC_net), .CO(n38258));
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n38256), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n2529), .I1(n34507), .I2(n2530), .I3(n2531), 
            .O(n43213));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n2517), .I1(n43213), .I2(n2518), .I3(n45218), 
            .O(n45224));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n45224), 
            .O(n45230));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hfffe;
    SB_LUT4 i33616_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n45230), 
            .O(n2544));
    defparam i33616_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY add_29_27 (.CI(n37185), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n37186));
    SB_LUT4 encoder0_position_31__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1720_rep_18_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1720_rep_18_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n37184), .O(n666)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_26 (.CI(n37184), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n37185));
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n38379), .I0(n2913), 
            .I1(VCC_net), .CO(n38380));
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n38378), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1724_rep_14_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1724_rep_14_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n38256), .I0(n2529), 
            .I1(GND_net), .CO(n38257));
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n38255), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1738 (.I0(n2626), .I1(n2628), .I2(GND_net), .I3(GND_net), 
            .O(n45526));
    defparam i1_2_lut_adj_1738.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n2622), .I1(n2621), .I2(n2623), .I3(n2624), 
            .O(n45534));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n2627), .I1(n45534), .I2(n45526), .I3(n2625), 
            .O(n45536));
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'hfffe;
    SB_LUT4 i21453_3_lut (.I0(n645), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n34501));
    defparam i21453_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n2618), .I1(n2619), .I2(n45536), .I3(n2620), 
            .O(n45542));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n38378), .I0(n2914), 
            .I1(VCC_net), .CO(n38379));
    SB_LUT4 i1_4_lut_adj_1742 (.I0(n2629), .I1(n34501), .I2(n2630), .I3(n2631), 
            .O(n43254));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n38255), .I0(n2530), 
            .I1(GND_net), .CO(n38256));
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n2616), .I1(n2617), .I2(n43254), .I3(n45542), 
            .O(n45548));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n45548), 
            .O(n45554));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'hfffe;
    SB_LUT4 i33670_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n45554), 
            .O(n2643));
    defparam i33670_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1722_rep_20_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1722_rep_20_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n38254), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1745 (.I0(n2727), .I1(n2725), .I2(GND_net), .I3(GND_net), 
            .O(n45000));
    defparam i1_2_lut_adj_1745.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1746 (.I0(n2724), .I1(n2721), .I2(n2722), .I3(n2728), 
            .O(n45002));
    defparam i1_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n2723), .I1(n2720), .I2(n45000), .I3(n2726), 
            .O(n45006));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'hfffe;
    SB_LUT4 i21547_4_lut (.I0(n646), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n34597));
    defparam i21547_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n2718), .I1(n2719), .I2(n45006), .I3(n45002), 
            .O(n45012));
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 add_29_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n37161), .O(n689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n38377), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n38254), .I0(n2531), 
            .I1(VCC_net), .CO(n38255));
    SB_LUT4 i1_4_lut_adj_1749 (.I0(n2729), .I1(n45012), .I2(n34597), .I3(n2730), 
            .O(n45014));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n2715), .I1(n2716), .I2(n45014), .I3(n2717), 
            .O(n45020));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_LUT4 add_29_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n37183), .O(n667)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n38377), .I0(n2915), 
            .I1(VCC_net), .CO(n38378));
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n38253), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n38253), .I0(n2532), 
            .I1(GND_net), .CO(n38254));
    SB_LUT4 i1_4_lut_adj_1751 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n45020), 
            .O(n45026));
    defparam i1_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_LUT4 i33956_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n45026), 
            .O(n2742));
    defparam i33956_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i7_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i33244_3_lut (.I0(n2726), .I1(n2793), .I2(n2742), .I3(GND_net), 
            .O(n2825));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n37167), .O(n683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33242_3_lut (.I0(n2725), .I1(n2792), .I2(n2742), .I3(GND_net), 
            .O(n2824));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n2824), .I1(n2825), .I2(n2823), .I3(n2827), 
            .O(n45494));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1753 (.I0(n45494), .I1(n2820), .I2(n2828), .I3(GND_net), 
            .O(n45496));
    defparam i1_3_lut_adj_1753.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n2819), .I1(n2826), .I2(n2822), .I3(n2821), 
            .O(n45498));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 i21545_4_lut (.I0(n647), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n34595));
    defparam i21545_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n2817), .I1(n2818), .I2(n45498), .I3(n45496), 
            .O(n45504));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n2829), .I1(n45504), .I2(n34595), .I3(n2830), 
            .O(n45506));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n45506), 
            .O(n45512));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n45512), 
            .O(n45518));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n38376), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n38252), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33987_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n45518), 
            .O(n2841));
    defparam i33987_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_9 (.CI(n37167), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n37168));
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n5722), 
            .D(n677), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n38376), .I0(n2916), 
            .I1(VCC_net), .CO(n38377));
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1759 (.I0(n2920), .I1(n2927), .I2(GND_net), .I3(GND_net), 
            .O(n45300));
    defparam i1_2_lut_adj_1759.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n2921), .I1(n2928), .I2(n2923), .I3(n2926), 
            .O(n45308));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n2924), .I1(n2919), .I2(n45300), .I3(n2922), 
            .O(n45310));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hfffe;
    SB_CARRY add_29_25 (.CI(n37183), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n37184));
    SB_LUT4 i21543_4_lut (.I0(n648), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n34593));
    defparam i21543_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 add_29_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n37166), .O(n684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n2917), .I1(n2918), .I2(n45310), .I3(n45308), 
            .O(n45316));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n38375), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n38252), .I0(n2533), 
            .I1(VCC_net), .CO(n38253));
    SB_LUT4 add_29_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n37182), .O(n668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n2929), .I1(n45316), .I2(n34593), .I3(n2930), 
            .O(n45318));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_adj_1764 (.I0(n2915), .I1(n2916), .I2(n2925), .I3(GND_net), 
            .O(n44972));
    defparam i1_3_lut_adj_1764.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n2912), .I1(n2910), .I2(n2914), .I3(n45318), 
            .O(n44442));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n2909), .I1(n2911), .I2(n2913), .I3(n44972), 
            .O(n44978));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hfffe;
    SB_LUT4 i34019_4_lut (.I0(n2908), .I1(n2907), .I2(n44978), .I3(n44442), 
            .O(n2940));
    defparam i34019_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n648));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n644), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n38375), .I0(n2917), 
            .I1(VCC_net), .CO(n38376));
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n644), 
            .I1(GND_net), .CO(n38252));
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n38374), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n648), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_24 (.CI(n37182), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n37183));
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n49231), .I1(n2412), 
            .I2(VCC_net), .I3(n38251), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_82_i8_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n649));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_82_i9_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i21443_3_lut (.I0(n649), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n34491));
    defparam i21443_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n3020), .I1(n3023), .I2(n3028), .I3(n3027), 
            .O(n45574));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1768 (.I0(n3021), .I1(n3019), .I2(n3024), .I3(GND_net), 
            .O(n45572));
    defparam i1_3_lut_adj_1768.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_82_i10_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[9]), 
            .I3(encoder0_position_scaled[9]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n38374), .I0(n2918), 
            .I1(VCC_net), .CO(n38375));
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n38250), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n45572), .I1(n45574), .I2(n3025), .I3(n3022), 
            .O(n45578));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n38250), .I0(n2413), 
            .I1(VCC_net), .CO(n38251));
    SB_CARRY add_29_3 (.CI(n37161), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n37162));
    SB_LUT4 i1_4_lut_adj_1770 (.I0(n3029), .I1(n34491), .I2(n3030), .I3(n3031), 
            .O(n43282));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(n3013), .I1(n3015), .I2(n43282), .I3(n45578), 
            .O(n45584));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n3016), .I1(n3017), .I2(n3018), .I3(n3026), 
            .O(n45598));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n3009), .I1(n3011), .I2(n3012), .I3(n45584), 
            .O(n45590));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n3008), .I1(n3010), .I2(n3014), .I3(n45598), 
            .O(n45604));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i34052_4_lut (.I0(n3007), .I1(n45604), .I2(n45590), .I3(n3006), 
            .O(n3039));
    defparam i34052_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n3125), .I1(n3119), .I2(n3118), .I3(n3120), 
            .O(n45044));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n3117), .I1(n3124), .I2(n3121), .I3(n3122), 
            .O(n45048));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n3126), .I1(n3123), .I2(n3127), .I3(n3128), 
            .O(n45046));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_LUT4 i21439_3_lut (.I0(n650), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n34487));
    defparam i21439_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n45046), .I1(n3116), .I2(n45048), .I3(n45044), 
            .O(n45054));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n3129), .I1(n34487), .I2(n3130), .I3(n3131), 
            .O(n43242));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n3114), .I1(n43242), .I2(n3115), .I3(n45054), 
            .O(n45060));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n45060), 
            .O(n45066));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n45066), 
            .O(n45072));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'hfffe;
    SB_LUT4 i34086_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n45072), 
            .O(n3138));
    defparam i34086_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i11_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[10]), 
            .I3(encoder0_position_scaled[10]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_5001), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n628));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_82_i12_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[11]), 
            .I3(encoder0_position_scaled[11]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i641_3_lut (.I0(n628), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n38249), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_8 (.CI(n37166), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n37167));
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n38249), .I0(n2414), 
            .I1(VCC_net), .CO(n38250));
    SB_LUT4 i15338_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n42230), 
            .I3(GND_net), .O(n28397));   // verilog/coms.v(127[12] 300[6])
    defparam i15338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15339_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n42230), 
            .I3(GND_net), .O(n28398));   // verilog/coms.v(127[12] 300[6])
    defparam i15339_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n38373), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n38248), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_700_i30_3_lut (.I0(n12_adj_5040), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30_adj_5050));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n38373), .I0(n2919), 
            .I1(VCC_net), .CO(n38374));
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n38372), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13_adj_4997), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n632));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i913_3_lut (.I0(n632), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_5002), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n627));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i573_3_lut (.I0(n627), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i13_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[12]), 
            .I3(encoder0_position_scaled[12]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33418_3_lut (.I0(n48370), .I1(pwm_setpoint[14]), .I2(n29_adj_5049), 
            .I3(GND_net), .O(n48371));   // verilog/pwm.v(21[8:24])
    defparam i33418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15340_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n42230), 
            .I3(GND_net), .O(n28399));   // verilog/coms.v(127[12] 300[6])
    defparam i15340_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15341_3_lut (.I0(\data_in_frame[8] [4]), .I1(rx_data[4]), .I2(n42230), 
            .I3(GND_net), .O(n28400));   // verilog/coms.v(127[12] 300[6])
    defparam i15341_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32730_4_lut (.I0(n33_adj_5052), .I1(n31_adj_5051), .I2(n29_adj_5049), 
            .I3(n47691), .O(n47683));
    defparam i32730_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i15342_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n42230), 
            .I3(GND_net), .O(n28401));   // verilog/coms.v(127[12] 300[6])
    defparam i15342_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i14_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[13]), 
            .I3(encoder0_position_scaled[13]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i33486_4_lut (.I0(n30_adj_5050), .I1(n10_adj_5038), .I2(n35), 
            .I3(n47676), .O(n48439));   // verilog/pwm.v(21[8:24])
    defparam i33486_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i21527_4_lut (.I0(n627), .I1(n831), .I2(n832), .I3(n833), 
            .O(n34577));
    defparam i21527_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i33338_3_lut (.I0(n48371), .I1(pwm_setpoint[15]), .I2(n31_adj_5051), 
            .I3(GND_net), .O(n48291));   // verilog/pwm.v(21[8:24])
    defparam i33338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21634_4_lut (.I0(n829), .I1(n828), .I2(n34577), .I3(n830), 
            .O(n861));
    defparam i21634_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15343_3_lut (.I0(\data_in_frame[8] [2]), .I1(rx_data[2]), .I2(n42230), 
            .I3(GND_net), .O(n28402));   // verilog/coms.v(127[12] 300[6])
    defparam i15343_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15344_3_lut (.I0(\data_in_frame[8] [1]), .I1(rx_data[1]), .I2(n42230), 
            .I3(GND_net), .O(n28403));   // verilog/coms.v(127[12] 300[6])
    defparam i15344_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19_adj_4991), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n638));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1321_3_lut (.I0(n638), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18_adj_4992), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n637));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1253_3_lut (.I0(n637), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15156_4_lut (.I0(n27824), .I1(r_Bit_Index[0]), .I2(n42126), 
            .I3(r_SM_Main[1]), .O(n28215));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15156_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_82_i15_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[14]), 
            .I3(encoder0_position_scaled[14]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_82_i16_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[15]), 
            .I3(encoder0_position_scaled[15]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_4995), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n634));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n634), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15346_3_lut (.I0(\data_in_frame[8] [0]), .I1(rx_data[0]), .I2(n42230), 
            .I3(GND_net), .O(n28405));   // verilog/coms.v(127[12] 300[6])
    defparam i15346_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_5000), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n629));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28077_3_lut (.I0(n3_adj_5021), .I1(n6538), .I2(n42948), .I3(GND_net), 
            .O(n42949));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i709_3_lut (.I0(n629), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33275_3_lut (.I0(n6_adj_5034), .I1(pwm_setpoint[10]), .I2(n21_adj_5045), 
            .I3(GND_net), .O(n48228));   // verilog/pwm.v(21[8:24])
    defparam i33275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33086_3_lut (.I0(n1851), .I1(n1752), .I2(n1653), .I3(GND_net), 
            .O(n48039));
    defparam i33086_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 encoder0_position_31__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1111_rep_61_3_lut (.I0(n1695), .I1(n1794), 
            .I2(n1752), .I3(GND_net), .O(n46605));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1111_rep_61_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1178_rep_50_3_lut (.I0(n46605), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n46594));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1178_rep_50_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28078_3_lut (.I0(encoder0_position[30]), .I1(n42949), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i28078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33276_3_lut (.I0(n48228), .I1(pwm_setpoint[11]), .I2(n23_adj_5046), 
            .I3(GND_net), .O(n48229));   // verilog/pwm.v(21[8:24])
    defparam i33276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_29_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n37181), .O(n669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n38248), .I0(n2415), 
            .I1(VCC_net), .CO(n38249));
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n38247), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33328_3_lut (.I0(n1925), .I1(n1992), .I2(n1950), .I3(GND_net), 
            .O(n2024));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33328_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n5722), 
            .D(n678), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i21525_4_lut (.I0(n628), .I1(n931), .I2(n932), .I3(n933), 
            .O(n34575));
    defparam i21525_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 mux_82_i17_3_lut_4_lut (.I0(n26489), .I1(control_mode[1]), .I2(motor_state_23__N_106[16]), 
            .I3(encoder0_position_scaled[16]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_82_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15153_4_lut (.I0(n27820), .I1(r_Bit_Index_adj_5163[0]), .I2(n42123), 
            .I3(r_SM_Main_adj_5161[1]), .O(n28212));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15153_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_4999), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n630));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n34306), .I1(n43073), .I2(state_adj_5154[0]), 
            .I3(read), .O(n41841));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'h8280;
    SB_LUT4 encoder0_position_31__I_0_i777_3_lut (.I0(n630), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n38247), .I0(n2416), 
            .I1(VCC_net), .CO(n38248));
    SB_CARRY add_29_23 (.CI(n37181), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n37182));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5057), .I3(n38679), .O(n2_adj_5022)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5058), .I3(n38678), .O(n3_adj_5021)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n38678), 
            .I0(GND_net), .I1(n3_adj_5058), .CO(n38679));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5059), .I3(n38677), .O(n4_adj_5020)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n38677), 
            .I0(GND_net), .I1(n4_adj_5059), .CO(n38678));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5060), .I3(n38676), .O(n5_adj_5019)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n38676), 
            .I0(GND_net), .I1(n5_adj_5060), .CO(n38677));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5061), .I3(n38675), .O(n6_adj_5018)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n38675), 
            .I0(GND_net), .I1(n6_adj_5061), .CO(n38676));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5062), .I3(n38674), .O(n7_adj_5003)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n38372), .I0(n2920), 
            .I1(VCC_net), .CO(n38373));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n38674), 
            .I0(GND_net), .I1(n7_adj_5062), .CO(n38675));
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n38246), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5063), .I3(n38673), .O(n8_adj_5002)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n38673), 
            .I0(GND_net), .I1(n8_adj_5063), .CO(n38674));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5064), .I3(n38672), .O(n9_adj_5001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n38672), 
            .I0(GND_net), .I1(n9_adj_5064), .CO(n38673));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5065), .I3(n38671), .O(n10_adj_5000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n38671), 
            .I0(GND_net), .I1(n10_adj_5065), .CO(n38672));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5066), .I3(n38670), .O(n11_adj_4999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n38670), 
            .I0(GND_net), .I1(n11_adj_5066), .CO(n38671));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5067), .I3(n38669), .O(n12_adj_4998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n38246), .I0(n2417), 
            .I1(VCC_net), .CO(n38247));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n38669), 
            .I0(GND_net), .I1(n12_adj_5067), .CO(n38670));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5068), .I3(n38668), .O(n13_adj_4997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n38668), 
            .I0(GND_net), .I1(n13_adj_5068), .CO(n38669));
    SB_LUT4 add_78_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n37214), .O(encoder1_position_scaled_23__N_58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5069), .I3(n38667), .O(n14_adj_4996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n38667), 
            .I0(GND_net), .I1(n14_adj_5069), .CO(n38668));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5070), .I3(n38666), .O(n15_adj_4995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n37180), .O(n670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n38666), 
            .I0(GND_net), .I1(n15_adj_5070), .CO(n38667));
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n38371), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5071), .I3(n38665), .O(n16_adj_4994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n38245), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n38665), 
            .I0(GND_net), .I1(n16_adj_5071), .CO(n38666));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5072), .I3(n38664), .O(n17_adj_4993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n38664), 
            .I0(GND_net), .I1(n17_adj_5072), .CO(n38665));
    SB_LUT4 add_78_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n37213), .O(encoder1_position_scaled_23__N_58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5073), .I3(n38663), .O(n18_adj_4992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n38663), 
            .I0(GND_net), .I1(n18_adj_5073), .CO(n38664));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5074), .I3(n38662), .O(n19_adj_4991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n38662), 
            .I0(GND_net), .I1(n19_adj_5074), .CO(n38663));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5075), .I3(n38661), .O(n20_adj_4990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n38661), 
            .I0(GND_net), .I1(n20_adj_5075), .CO(n38662));
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n38245), .I0(n2418), 
            .I1(VCC_net), .CO(n38246));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5076), .I3(n38660), .O(n21_adj_4989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n38660), 
            .I0(GND_net), .I1(n21_adj_5076), .CO(n38661));
    SB_CARRY add_78_24 (.CI(n37213), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n37214));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5077), .I3(n38659), .O(n22_adj_4988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n38659), 
            .I0(GND_net), .I1(n22_adj_5077), .CO(n38660));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5078), .I3(n38658), .O(n23_adj_4987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n38658), 
            .I0(GND_net), .I1(n23_adj_5078), .CO(n38659));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5079), .I3(n38657), .O(n24_adj_4986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n38657), 
            .I0(GND_net), .I1(n24_adj_5079), .CO(n38658));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5080), .I3(n38656), .O(n25_adj_4985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n38371), .I0(n2921), 
            .I1(VCC_net), .CO(n38372));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n38656), 
            .I0(GND_net), .I1(n25_adj_5080), .CO(n38657));
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n38244), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5081), .I3(n38655), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n38655), 
            .I0(GND_net), .I1(n26_adj_5081), .CO(n38656));
    SB_CARRY add_29_22 (.CI(n37180), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n37181));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5082), .I3(n38654), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n38654), 
            .I0(GND_net), .I1(n27_adj_5082), .CO(n38655));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5083), .I3(n38653), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n38653), 
            .I0(GND_net), .I1(n28_adj_5083), .CO(n38654));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5084), .I3(n38652), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n38652), 
            .I0(GND_net), .I1(n29_adj_5084), .CO(n38653));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5085), .I3(n38651), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n38370), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n38651), 
            .I0(GND_net), .I1(n30_adj_5085), .CO(n38652));
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n38244), .I0(n2419), 
            .I1(VCC_net), .CO(n38245));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5086), .I3(n38650), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n38650), 
            .I0(GND_net), .I1(n31_adj_5086), .CO(n38651));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5087), .I3(n38649), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n38649), 
            .I0(GND_net), .I1(n32_adj_5087), .CO(n38650));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5088), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5088), .CO(n38649));
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n38243), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n37212), .O(encoder1_position_scaled_23__N_58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33084_3_lut (.I0(n1950), .I1(n1851), .I2(n1752), .I3(GND_net), 
            .O(n48037));
    defparam i33084_3_lut.LUT_INIT = 16'h7f7f;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n38370), .I0(n2922), 
            .I1(VCC_net), .CO(n38371));
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n38243), .I0(n2420), 
            .I1(VCC_net), .CO(n38244));
    SB_LUT4 add_1894_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n37551), 
            .O(n6537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1894_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1894_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n37550), 
            .O(n6538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1894_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1894_6 (.CI(n37550), .I0(n622), .I1(GND_net), .CO(n37551));
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n38242), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n27784), 
            .I3(rx_data_ready), .O(n41813));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_CARRY add_78_23 (.CI(n37212), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n37213));
    SB_LUT4 add_29_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1894_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n37549), 
            .O(n6539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1894_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1894_5 (.CI(n37549), .I0(n623), .I1(VCC_net), .CO(n37550));
    SB_LUT4 i33028_3_lut_4_lut (.I0(n2148), .I1(n2049), .I2(n2028), .I3(n46578), 
            .O(n2226));
    defparam i33028_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 add_1894_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n37548), 
            .O(n6540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1894_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1179_rep_54_3_lut (.I0(n1795), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n46598));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1179_rep_54_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1246_rep_44_3_lut (.I0(n46598), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n46588));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1246_rep_44_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n38369), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1894_4 (.CI(n37548), .I0(n516), .I1(GND_net), .CO(n37549));
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n38242), .I0(n2421), 
            .I1(VCC_net), .CO(n38243));
    SB_LUT4 i33332_3_lut (.I0(n2025), .I1(n2092), .I2(n2049), .I3(GND_net), 
            .O(n2124));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1894_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n37547), 
            .O(n6541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1894_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1894_3 (.CI(n37547), .I0(n625), .I1(VCC_net), .CO(n37548));
    SB_LUT4 add_1894_2_lut (.I0(GND_net), .I1(n626), .I2(GND_net), .I3(VCC_net), 
            .O(n6542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1894_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1894_2 (.CI(VCC_net), .I0(n626), .I1(GND_net), .CO(n37547));
    SB_LUT4 encoder0_position_31__I_0_i1384_rep_32_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1384_rep_32_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20_adj_4990), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n639));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33070_4_lut (.I0(n23_adj_5046), .I1(n21_adj_5045), .I2(n19_adj_5044), 
            .I3(n47726), .O(n48023));
    defparam i33070_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 encoder0_position_31__I_0_i1389_3_lut (.I0(n639), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21_adj_4989), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n640));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n640), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n17_adj_4952));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22_adj_4988), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n641));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n28747));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n28746));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n28745));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n28744));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n28743));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n28742));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n28741));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1784 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n45184));
    defparam i1_2_lut_adj_1784.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_4998), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n631));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i845_3_lut (.I0(n631), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33335_3_lut (.I0(n8_adj_5036), .I1(pwm_setpoint[9]), .I2(n19_adj_5044), 
            .I3(GND_net), .O(n48288));   // verilog/pwm.v(21[8:24])
    defparam i33335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1180_rep_52_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1180_rep_52_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33330_3_lut (.I0(n1927), .I1(n1994), .I2(n1950), .I3(GND_net), 
            .O(n2026));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i33330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1452_rep_30_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1452_rep_30_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n2225), .I1(n2228), .I2(n2226), .I3(n2224), 
            .O(n45424));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n927), .I1(n45184), .I2(n928), .I3(n34575), 
            .O(n960));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hfefa;
    SB_LUT4 i33037_3_lut (.I0(n48229), .I1(pwm_setpoint[12]), .I2(n25_adj_5047), 
            .I3(GND_net), .O(n47990));   // verilog/pwm.v(21[8:24])
    defparam i33037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33333_4_lut (.I0(n33_adj_5052), .I1(n31_adj_5051), .I2(n29_adj_5049), 
            .I3(n47693), .O(n48286));
    defparam i33333_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21400_3_lut (.I0(n629), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n34447));
    defparam i21400_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i21476_3_lut (.I0(n641), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n34525));
    defparam i21476_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n2222), .I1(n45424), .I2(n2223), .I3(n2227), 
            .O(n45428));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'hfffe;
    SB_LUT4 i33525_4_lut (.I0(n48291), .I1(n48439), .I2(n35), .I3(n47683), 
            .O(n48478));   // verilog/pwm.v(21[8:24])
    defparam i33525_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n2229), .I1(n34525), .I2(n2230), .I3(n2231), 
            .O(n43224));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n2220), .I1(n43224), .I2(n2221), .I3(n45428), 
            .O(n45434));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n45434), 
            .O(n45440));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 i34231_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n45440), 
            .O(n2247));
    defparam i34231_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15229_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n27752), .I3(GND_net), .O(n28288));   // verilog/coms.v(127[12] 300[6])
    defparam i15229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15230_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n27752), .I3(GND_net), .O(n28289));   // verilog/coms.v(127[12] 300[6])
    defparam i15230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15231_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n27752), .I3(GND_net), .O(n28290));   // verilog/coms.v(127[12] 300[6])
    defparam i15231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15232_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n27752), .I3(GND_net), .O(n28291));   // verilog/coms.v(127[12] 300[6])
    defparam i15232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n1029), .I1(n34447), .I2(n1030), .I3(n1031), 
            .O(n43139));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'ha080;
    SB_LUT4 i33413_4_lut (.I0(n47990), .I1(n48288), .I2(n25_adj_5047), 
            .I3(n48023), .O(n48366));   // verilog/pwm.v(21[8:24])
    defparam i33413_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33746_4_lut (.I0(n1026), .I1(n43139), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i33746_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33543_4_lut (.I0(n48366), .I1(n48478), .I2(n35), .I3(n48286), 
            .O(n48496));   // verilog/pwm.v(21[8:24])
    defparam i33543_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i21521_4_lut (.I0(n630), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n34571));
    defparam i21521_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i33544_3_lut (.I0(n48496), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n48497));   // verilog/pwm.v(21[8:24])
    defparam i33544_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1792 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n44966));
    defparam i1_3_lut_adj_1792.LUT_INIT = 16'hfefe;
    SB_LUT4 i33542_3_lut (.I0(n48497), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n48495));   // verilog/pwm.v(21[8:24])
    defparam i33542_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n38241), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n38241), .I0(n2422), 
            .I1(VCC_net), .CO(n38242));
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n38240), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n38369), .I0(n2923), 
            .I1(VCC_net), .CO(n38370));
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n38240), .I0(n2423), 
            .I1(VCC_net), .CO(n38241));
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n5722), 
            .D(n679), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 add_29_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n37179), .O(n671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n38368), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n38368), .I0(n2924), 
            .I1(VCC_net), .CO(n38369));
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n38239), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n38239), .I0(n2424), 
            .I1(VCC_net), .CO(n38240));
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5030));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n38367), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1400_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n777), .I3(n26487), .O(n5855));   // verilog/TinyFPGA_B.v(262[5] 286[12])
    defparam i1400_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n38238), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15162_3_lut_4_lut (.I0(n1152), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_3807), .O(n28221));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15162_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i26_4_lut (.I0(n47524), .I1(n47523), .I2(state[1]), .I3(n30301), 
            .O(n12_adj_5053));   // verilog/neopixel.v(35[12] 117[6])
    defparam i26_4_lut.LUT_INIT = 16'h3530;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n38238), .I0(n2425), 
            .I1(VCC_net), .CO(n38239));
    SB_LUT4 i15157_3_lut_4_lut (.I0(n1193), .I1(b_prev_adj_5011), .I2(a_new_adj_5130[1]), 
            .I3(direction_N_3807_adj_5012), .O(n28216));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15157_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n38367), .I0(n2925), 
            .I1(VCC_net), .CO(n38368));
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n38237), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15143_4_lut (.I0(state_7__N_4003[3]), .I1(data[0]), .I2(n10_adj_5097), 
            .I3(n26652), .O(n28202));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15143_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n44886));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n38237), .I0(n2426), 
            .I1(VCC_net), .CO(n38238));
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n38366), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n38366), .I0(n2926), 
            .I1(VCC_net), .CO(n38367));
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n38236), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n37211), .O(encoder1_position_scaled_23__N_58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1793 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n45286));
    defparam i1_2_lut_adj_1793.LUT_INIT = 16'h8888;
    SB_LUT4 i33767_4_lut (.I0(n45286), .I1(n1125), .I2(n44966), .I3(n34571), 
            .O(n1158));
    defparam i33767_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_31__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21393_3_lut (.I0(n631), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n34439));
    defparam i21393_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1794 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n45290));
    defparam i1_3_lut_adj_1794.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n1229), .I1(n34439), .I2(n1230), .I3(n1231), 
            .O(n43134));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'ha080;
    SB_LUT4 i33471_3_lut (.I0(n48495), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n48424));   // verilog/pwm.v(21[8:24])
    defparam i33471_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33782_4_lut (.I0(n1225), .I1(n1224), .I2(n43134), .I3(n45290), 
            .O(n1257));
    defparam i33782_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i769_3_lut (.I0(n1126), .I1(n1193_adj_5029), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21334_3_lut (.I0(n632), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n34379));
    defparam i21334_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n44988));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n1329), .I1(n34379), .I2(n1330), .I3(n1331), 
            .O(n43131));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'ha080;
    SB_LUT4 i33801_4_lut (.I0(n43131), .I1(n1323), .I2(n1324), .I3(n44988), 
            .O(n1356));
    defparam i33801_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21332_3_lut (.I0(n633), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n34377));
    defparam i21332_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i33472_3_lut (.I0(n48424), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n48425));   // verilog/pwm.v(21[8:24])
    defparam i33472_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1798 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n45326));
    defparam i1_2_lut_adj_1798.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n1429), .I1(n34377), .I2(n1430), .I3(n1431), 
            .O(n43150));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n45326), 
            .O(n45332));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'hfffe;
    SB_LUT4 i33820_4_lut (.I0(n1423), .I1(n1422), .I2(n45332), .I3(n43150), 
            .O(n1455));
    defparam i33820_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1801 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n45188));
    defparam i1_2_lut_adj_1801.LUT_INIT = 16'heeee;
    SB_LUT4 i21508_4_lut (.I0(n634), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n34557));
    defparam i21508_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i33344_3_lut (.I0(n48425), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n48297));   // verilog/pwm.v(21[8:24])
    defparam i33344_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1802 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n45188), 
            .O(n45194));
    defparam i1_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n1529), .I1(n45194), .I2(n34557), .I3(n1530), 
            .O(n45196));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'heccc;
    SB_LUT4 i33838_4_lut (.I0(n1522), .I1(n1521), .I2(n45196), .I3(n1523), 
            .O(n1554));
    defparam i33838_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21328_3_lut (.I0(n635), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n34373));
    defparam i21328_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n45344));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n1629), .I1(n34373), .I2(n1630), .I3(n1631), 
            .O(n43159));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_4996), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n633));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n1623), .I1(n43159), .I2(n1624), .I3(n45344), 
            .O(n45350));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 i33860_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n45350), 
            .O(n1653));
    defparam i33860_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n38365), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1807 (.I0(n1728), .I1(n1726), .I2(n1727), .I3(GND_net), 
            .O(n45264));
    defparam i1_3_lut_adj_1807.LUT_INIT = 16'hfefe;
    SB_LUT4 i21502_4_lut (.I0(n636), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n34551));
    defparam i21502_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n1723), .I1(n1724), .I2(n45264), .I3(n1725), 
            .O(n45270));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1809 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n45356));
    defparam i1_2_lut_adj_1809.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i981_3_lut (.I0(n633), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n45356), .I1(n1722), .I2(n45270), .I3(n34551), 
            .O(n45274));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hfefc;
    SB_LUT4 i33886_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n45274), 
            .O(n1752));
    defparam i33886_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n38236), .I0(n2427), 
            .I1(VCC_net), .CO(n38237));
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position_scaled[23]), 
            .I2(n2), .I3(n37494), .O(displacement_23__N_82[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n1825), .I1(n1826), .I2(n1827), .I3(n1828), 
            .O(n45366));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position_scaled[22]), 
            .I2(n3_adj_5004), .I3(n37493), .O(displacement_23__N_82[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_24 (.CI(n37493), .I0(encoder1_position_scaled[22]), 
            .I1(n3_adj_5004), .CO(n37494));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position_scaled[21]), 
            .I2(n4_adj_5005), .I3(n37492), .O(displacement_23__N_82[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_23 (.CI(n37492), .I0(encoder1_position_scaled[21]), 
            .I1(n4_adj_5005), .CO(n37493));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position_scaled[20]), 
            .I2(n5_adj_4953), .I3(n37491), .O(displacement_23__N_82[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_22 (.CI(n37491), .I0(encoder1_position_scaled[20]), 
            .I1(n5_adj_4953), .CO(n37492));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position_scaled[19]), 
            .I2(n6_adj_4954), .I3(n37490), .O(displacement_23__N_82[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_21 (.CI(n37490), .I0(encoder1_position_scaled[19]), 
            .I1(n6_adj_4954), .CO(n37491));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position_scaled[18]), 
            .I2(n7_adj_4955), .I3(n37489), .O(displacement_23__N_82[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_20 (.CI(n37489), .I0(encoder1_position_scaled[18]), 
            .I1(n7_adj_4955), .CO(n37490));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n38235), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n38365), .I0(n2927), 
            .I1(VCC_net), .CO(n38366));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position_scaled[17]), 
            .I2(n8_adj_4956), .I3(n37488), .O(displacement_23__N_82[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_19 (.CI(n37488), .I0(encoder1_position_scaled[17]), 
            .I1(n8_adj_4956), .CO(n37489));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position_scaled[16]), 
            .I2(n9_adj_4957), .I3(n37487), .O(displacement_23__N_82[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_18 (.CI(n37487), .I0(encoder1_position_scaled[16]), 
            .I1(n9_adj_4957), .CO(n37488));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position_scaled[15]), 
            .I2(n10_adj_4958), .I3(n37486), .O(displacement_23__N_82[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF h1_56 (.Q(INLA_c), .C(CLK_c), .D(hall1));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_17 (.CI(n37486), .I0(encoder1_position_scaled[15]), 
            .I1(n10_adj_4958), .CO(n37487));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position_scaled[14]), 
            .I2(n11_adj_4959), .I3(n37485), .O(displacement_23__N_82[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_16 (.CI(n37485), .I0(encoder1_position_scaled[14]), 
            .I1(n11_adj_4959), .CO(n37486));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position_scaled[13]), 
            .I2(n12_adj_4960), .I3(n37484), .O(displacement_23__N_82[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_15 (.CI(n37484), .I0(encoder1_position_scaled[13]), 
            .I1(n12_adj_4960), .CO(n37485));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position_scaled[12]), 
            .I2(n13_adj_4961), .I3(n37483), .O(displacement_23__N_82[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_14 (.CI(n37483), .I0(encoder1_position_scaled[12]), 
            .I1(n13_adj_4961), .CO(n37484));
    SB_LUT4 i21320_3_lut (.I0(n637), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n34365));
    defparam i21320_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position_scaled[11]), 
            .I2(n14_adj_4962), .I3(n37482), .O(displacement_23__N_82[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_13 (.CI(n37482), .I0(encoder1_position_scaled[11]), 
            .I1(n14_adj_4962), .CO(n37483));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position_scaled[10]), 
            .I2(n15_adj_4963), .I3(n37481), .O(displacement_23__N_82[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_12 (.CI(n37481), .I0(encoder1_position_scaled[10]), 
            .I1(n15_adj_4963), .CO(n37482));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position_scaled[9]), 
            .I2(n16_adj_4964), .I3(n37480), .O(displacement_23__N_82[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_11 (.CI(n37480), .I0(encoder1_position_scaled[9]), 
            .I1(n16_adj_4964), .CO(n37481));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position_scaled[8]), 
            .I2(n17_adj_4965), .I3(n37479), .O(displacement_23__N_82[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_10 (.CI(n37479), .I0(encoder1_position_scaled[8]), 
            .I1(n17_adj_4965), .CO(n37480));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position_scaled[7]), 
            .I2(n18_adj_4966), .I3(n37478), .O(displacement_23__N_82[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_9 (.CI(n37478), .I0(encoder1_position_scaled[7]), 
            .I1(n18_adj_4966), .CO(n37479));
    SB_CARRY add_78_22 (.CI(n37211), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n37212));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position_scaled[6]), 
            .I2(n19_adj_4967), .I3(n37477), .O(displacement_23__N_82[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_8 (.CI(n37477), .I0(encoder1_position_scaled[6]), 
            .I1(n19_adj_4967), .CO(n37478));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position_scaled[5]), 
            .I2(n20_adj_4968), .I3(n37476), .O(displacement_23__N_82[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_7 (.CI(n37476), .I0(encoder1_position_scaled[5]), 
            .I1(n20_adj_4968), .CO(n37477));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position_scaled[4]), 
            .I2(n21_adj_4969), .I3(n37475), .O(displacement_23__N_82[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_21 (.CI(n37179), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n37180));
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_6 (.CI(n37475), .I0(encoder1_position_scaled[4]), 
            .I1(n21_adj_4969), .CO(n37476));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position_scaled[3]), 
            .I2(n22_adj_4970), .I3(n37474), .O(displacement_23__N_82[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_5 (.CI(n37474), .I0(encoder1_position_scaled[3]), 
            .I1(n22_adj_4970), .CO(n37475));
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n38235), .I0(n2428), 
            .I1(VCC_net), .CO(n38236));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position_scaled[2]), 
            .I2(n23_adj_4971), .I3(n37473), .O(displacement_23__N_82[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n37210), .O(encoder1_position_scaled_23__N_58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_78_21 (.CI(n37210), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n37211));
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_4 (.CI(n37473), .I0(encoder1_position_scaled[2]), 
            .I1(n23_adj_4971), .CO(n37474));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position_scaled[1]), 
            .I2(n24_adj_4972), .I3(n37472), .O(displacement_23__N_82[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_3 (.CI(n37472), .I0(encoder1_position_scaled[1]), 
            .I1(n24_adj_4972), .CO(n37473));
    SB_LUT4 encoder1_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position_scaled[0]), 
            .I2(n25_adj_4973), .I3(VCC_net), .O(displacement_23__N_82[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position_scaled[0]), 
            .I1(n25_adj_4973), .CO(n37472));
    SB_LUT4 add_674_24_lut (.I0(duty[22]), .I1(n49248), .I2(n3), .I3(n37471), 
            .O(pwm_setpoint_22__N_11[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n38364), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n38234), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n38364), .I0(n2928), 
            .I1(VCC_net), .CO(n38365));
    SB_LUT4 add_674_23_lut (.I0(duty[21]), .I1(n49248), .I2(n4), .I3(n37470), 
            .O(pwm_setpoint_22__N_11[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n38234), .I0(n2429), 
            .I1(GND_net), .CO(n38235));
    SB_CARRY add_674_23 (.CI(n37470), .I0(n49248), .I1(n4), .CO(n37471));
    SB_LUT4 add_674_22_lut (.I0(duty[20]), .I1(n49248), .I2(n5), .I3(n37469), 
            .O(pwm_setpoint_22__N_11[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_22 (.CI(n37469), .I0(n49248), .I1(n5), .CO(n37470));
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n38363), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n38233), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n38363), .I0(n2929), 
            .I1(GND_net), .CO(n38364));
    SB_LUT4 add_674_21_lut (.I0(duty[19]), .I1(n49248), .I2(n6), .I3(n37468), 
            .O(pwm_setpoint_22__N_11[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_21_lut.LUT_INIT = 16'h8BB8;
    GND i1 (.Y(GND_net));
    SB_CARRY add_674_21 (.CI(n37468), .I0(n49248), .I1(n6), .CO(n37469));
    SB_LUT4 add_78_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n37209), .O(encoder1_position_scaled_23__N_58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_674_20_lut (.I0(duty[18]), .I1(n49248), .I2(n7), .I3(n37467), 
            .O(pwm_setpoint_22__N_11[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_20 (.CI(n37467), .I0(n49248), .I1(n7), .CO(n37468));
    SB_LUT4 add_674_19_lut (.I0(duty[17]), .I1(n49248), .I2(n8), .I3(n37466), 
            .O(pwm_setpoint_22__N_11[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_19 (.CI(n37466), .I0(n49248), .I1(n8), .CO(n37467));
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n38233), .I0(n2430), 
            .I1(GND_net), .CO(n38234));
    SB_LUT4 add_29_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n37178), .O(n672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_674_18_lut (.I0(duty[16]), .I1(n49248), .I2(n9), .I3(n37465), 
            .O(pwm_setpoint_22__N_11[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_78_20 (.CI(n37209), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n37210));
    SB_CARRY add_674_18 (.CI(n37465), .I0(n49248), .I1(n9), .CO(n37466));
    SB_LUT4 add_78_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n37208), .O(encoder1_position_scaled_23__N_58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n38362), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n38232), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_674_17_lut (.I0(duty[15]), .I1(n49248), .I2(n10), .I3(n37464), 
            .O(pwm_setpoint_22__N_11[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_17 (.CI(n37464), .I0(n49248), .I1(n10), .CO(n37465));
    SB_LUT4 add_674_16_lut (.I0(duty[14]), .I1(n49248), .I2(n11), .I3(n37463), 
            .O(pwm_setpoint_22__N_11[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_3_lut_adj_1812 (.I0(n1823), .I1(n1824), .I2(n45366), .I3(GND_net), 
            .O(n45370));
    defparam i1_3_lut_adj_1812.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n38362), .I0(n2930), 
            .I1(GND_net), .CO(n38363));
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n38232), .I0(n2431), 
            .I1(VCC_net), .CO(n38233));
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_78_19 (.CI(n37208), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n37209));
    SB_CARRY add_674_16 (.CI(n37463), .I0(n49248), .I1(n11), .CO(n37464));
    SB_LUT4 add_674_15_lut (.I0(duty[13]), .I1(n49248), .I2(n12), .I3(n37462), 
            .O(pwm_setpoint_22__N_11[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n38231), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_674_15 (.CI(n37462), .I0(n49248), .I1(n12), .CO(n37463));
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n5722), 
            .D(n680), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 add_674_14_lut (.I0(duty[12]), .I1(n49248), .I2(n13), .I3(n37461), 
            .O(pwm_setpoint_22__N_11[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_14 (.CI(n37461), .I0(n49248), .I1(n13), .CO(n37462));
    SB_LUT4 add_674_13_lut (.I0(duty[11]), .I1(n49248), .I2(n14), .I3(n37460), 
            .O(pwm_setpoint_22__N_11[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_13 (.CI(n37460), .I0(n49248), .I1(n14), .CO(n37461));
    SB_LUT4 i1_2_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3442[2]), .O(n42185));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(n49181), .I1(n2214), 
            .I2(VCC_net), .I3(n38091), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_29_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n37165), .O(n685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_674_12_lut (.I0(duty[10]), .I1(n49248), .I2(n15_adj_4948), 
            .I3(n37459), .O(pwm_setpoint_22__N_11[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_12_lut.LUT_INIT = 16'h8BB8;
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n5722), 
            .D(n681), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n5722), 
            .D(n682), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY add_674_12 (.CI(n37459), .I0(n49248), .I1(n15_adj_4948), 
            .CO(n37460));
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n38361), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n5722), 
            .D(n683), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 add_674_11_lut (.I0(duty[9]), .I1(n49248), .I2(n16), .I3(n37458), 
            .O(pwm_setpoint_22__N_11[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n38231), .I0(n2432), 
            .I1(GND_net), .CO(n38232));
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n5722), 
            .D(n684), .R(n28104));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n38090), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_20 (.CI(n37178), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n37179));
    SB_LUT4 add_78_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n37207), .O(encoder1_position_scaled_23__N_58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_674_11 (.CI(n37458), .I0(n49248), .I1(n16), .CO(n37459));
    SB_LUT4 i16_4_lut_adj_1813 (.I0(state_adj_5170[0]), .I1(n47597), .I2(n5538), 
            .I3(n33499), .O(n8_adj_5089));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_adj_1813.LUT_INIT = 16'h3afa;
    SB_LUT4 add_674_10_lut (.I0(duty[8]), .I1(n49248), .I2(n17), .I3(n37457), 
            .O(pwm_setpoint_22__N_11[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_29_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n37161));
    SB_LUT4 add_29_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n37177), .O(n673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_674_10 (.CI(n37457), .I0(n49248), .I1(n17), .CO(n37458));
    SB_CARRY add_78_18 (.CI(n37207), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n37208));
    SB_LUT4 add_674_9_lut (.I0(duty[7]), .I1(n49248), .I2(n18), .I3(n37456), 
            .O(pwm_setpoint_22__N_11[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n38361), .I0(n2931), 
            .I1(VCC_net), .CO(n38362));
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n38230), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n38230), .I0(n2433), 
            .I1(VCC_net), .CO(n38231));
    SB_LUT4 add_78_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n37206), .O(encoder1_position_scaled_23__N_58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n38090), .I0(n2215), 
            .I1(VCC_net), .CO(n38091));
    SB_CARRY add_29_7 (.CI(n37165), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n37166));
    SB_CARRY add_29_19 (.CI(n37177), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n37178));
    SB_CARRY add_674_9 (.CI(n37456), .I0(n49248), .I1(n18), .CO(n37457));
    SB_LUT4 add_674_8_lut (.I0(duty[6]), .I1(n49248), .I2(n19), .I3(n37455), 
            .O(pwm_setpoint_22__N_11[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_8 (.CI(n37455), .I0(n49248), .I1(n19), .CO(n37456));
    SB_LUT4 add_29_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n37176), .O(n674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_674_7_lut (.I0(duty[5]), .I1(n49248), .I2(n20), .I3(n37454), 
            .O(pwm_setpoint_22__N_11[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_7 (.CI(n37454), .I0(n49248), .I1(n20), .CO(n37455));
    SB_CARRY add_78_17 (.CI(n37206), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n37207));
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n643), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n37205), .O(encoder1_position_scaled_23__N_58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_674_6_lut (.I0(duty[4]), .I1(n49248), .I2(n21), .I3(n37453), 
            .O(pwm_setpoint_22__N_11[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_78_16 (.CI(n37205), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n37206));
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_674_6 (.CI(n37453), .I0(n49248), .I1(n21), .CO(n37454));
    SB_LUT4 add_674_5_lut (.I0(duty[3]), .I1(n49248), .I2(n22), .I3(n37452), 
            .O(pwm_setpoint_22__N_11[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_29_18 (.CI(n37176), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n37177));
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n38360), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_674_5 (.CI(n37452), .I0(n49248), .I1(n22), .CO(n37453));
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n1829), .I1(n34365), .I2(n1830), .I3(n1831), 
            .O(n43196));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'ha080;
    SB_LUT4 add_674_4_lut (.I0(duty[2]), .I1(n49248), .I2(n23), .I3(n37451), 
            .O(pwm_setpoint_22__N_11[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_674_4 (.CI(n37451), .I0(n49248), .I1(n23), .CO(n37452));
    SB_LUT4 add_674_3_lut (.I0(duty[1]), .I1(n49248), .I2(n24), .I3(n37450), 
            .O(pwm_setpoint_22__N_11[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16_adj_4994), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n635));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_674_3 (.CI(n37450), .I0(n49248), .I1(n24), .CO(n37451));
    SB_LUT4 add_674_2_lut (.I0(duty[0]), .I1(n49248), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_11[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_674_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i32728_3_lut_4_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n34515), .I3(state[1]), .O(n47524));   // verilog/neopixel.v(35[12] 117[6])
    defparam i32728_3_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1815 (.I0(n1821), .I1(n1822), .I2(n43196), .I3(n45370), 
            .O(n45376));
    defparam i1_4_lut_adj_1815.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1117_3_lut (.I0(n635), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33911_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n45376), 
            .O(n1851));
    defparam i33911_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_674_2 (.CI(VCC_net), .I0(n49248), .I1(n25), .CO(n37450));
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n38089), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_78_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n37204), .O(encoder1_position_scaled_23__N_58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_78_15 (.CI(n37204), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n37205));
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n38360), .I0(n2932), 
            .I1(GND_net), .CO(n38361));
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n643), 
            .I1(GND_net), .CO(n38230));
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n38089), .I0(n2216), 
            .I1(VCC_net), .CO(n38090));
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n37973), .I0(n2132), 
            .I1(GND_net), .CO(n37974));
    SB_LUT4 add_78_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n37203), .O(encoder1_position_scaled_23__N_58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n37164), .O(n686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_700_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_5034));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n38088), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n37979), .I0(n2126), 
            .I1(VCC_net), .CO(n37980));
    SB_CARRY add_78_14 (.CI(n37203), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n37204));
    SB_LUT4 add_29_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n37175), .O(n675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_700_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_5038));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_78_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n37202), .O(encoder1_position_scaled_23__N_58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_78_13 (.CI(n37202), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n37203));
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n38359), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n49207), .I1(n2313), 
            .I2(VCC_net), .I3(n38229), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n38088), .I0(n2217), 
            .I1(VCC_net), .CO(n38089));
    SB_LUT4 encoder0_position_31__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15405_3_lut (.I0(\data_in_frame[0] [7]), .I1(rx_data[7]), .I2(n42229), 
            .I3(GND_net), .O(n28464));   // verilog/coms.v(127[12] 300[6])
    defparam i15405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15406_3_lut (.I0(\data_in_frame[0] [6]), .I1(rx_data[6]), .I2(n42229), 
            .I3(GND_net), .O(n28465));   // verilog/coms.v(127[12] 300[6])
    defparam i15406_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n38359), .I0(n2933), 
            .I1(VCC_net), .CO(n38360));
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n38228), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n38087), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n38087), .I0(n2218), 
            .I1(VCC_net), .CO(n38088));
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n38228), .I0(n2314), 
            .I1(VCC_net), .CO(n38229));
    SB_LUT4 add_78_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n37201), .O(encoder1_position_scaled_23__N_58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_78_12 (.CI(n37201), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n37202));
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_78_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n37200), .O(encoder1_position_scaled_23__N_58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15407_3_lut (.I0(\data_in_frame[0] [5]), .I1(rx_data[5]), .I2(n42229), 
            .I3(GND_net), .O(n28466));   // verilog/coms.v(127[12] 300[6])
    defparam i15407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n38086), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n648), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n38227), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n38086), .I0(n2219), 
            .I1(VCC_net), .CO(n38087));
    SB_CARRY add_29_17 (.CI(n37175), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n37176));
    SB_CARRY add_78_9 (.CI(n37198), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n37199));
    SB_LUT4 encoder0_position_31__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15408_3_lut (.I0(\data_in_frame[0] [4]), .I1(rx_data[4]), .I2(n42229), 
            .I3(GND_net), .O(n28467));   // verilog/coms.v(127[12] 300[6])
    defparam i15408_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n38227), .I0(n2315), 
            .I1(VCC_net), .CO(n38228));
    SB_LUT4 i32723_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n47676));
    defparam i32723_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n38085), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1944_25_lut (.I0(n48696), .I1(n2_adj_5057), .I2(n1059), 
            .I3(n38496), .O(encoder0_position_scaled_23__N_34[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1944_24_lut (.I0(n48717), .I1(n2_adj_5057), .I2(n1158), 
            .I3(n38495), .O(encoder0_position_scaled_23__N_34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_24 (.CI(n38495), .I0(n2_adj_5057), .I1(n1158), .CO(n38496));
    SB_LUT4 add_1944_23_lut (.I0(n48731), .I1(n2_adj_5057), .I2(n1257), 
            .I3(n38494), .O(encoder0_position_scaled_23__N_34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_23 (.CI(n38494), .I0(n2_adj_5057), .I1(n1257), .CO(n38495));
    SB_LUT4 add_1944_22_lut (.I0(n48750), .I1(n2_adj_5057), .I2(n1356), 
            .I3(n38493), .O(encoder0_position_scaled_23__N_34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_22 (.CI(n38493), .I0(n2_adj_5057), .I1(n1356), .CO(n38494));
    SB_LUT4 add_1944_21_lut (.I0(n48769), .I1(n2_adj_5057), .I2(n1455), 
            .I3(n38492), .O(encoder0_position_scaled_23__N_34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n38085), .I0(n2220), 
            .I1(VCC_net), .CO(n38086));
    SB_CARRY add_1944_21 (.CI(n38492), .I0(n2_adj_5057), .I1(n1455), .CO(n38493));
    SB_LUT4 add_1944_20_lut (.I0(n48787), .I1(n2_adj_5057), .I2(n1554), 
            .I3(n38491), .O(encoder0_position_scaled_23__N_34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_20 (.CI(n38491), .I0(n2_adj_5057), .I1(n1554), .CO(n38492));
    SB_LUT4 add_78_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n37199), .O(encoder1_position_scaled_23__N_58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_78_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1944_19_lut (.I0(n48808), .I1(n2_adj_5057), .I2(n1653), 
            .I3(n38490), .O(encoder0_position_scaled_23__N_34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_19 (.CI(n38490), .I0(n2_adj_5057), .I1(n1653), .CO(n38491));
    SB_LUT4 add_1944_18_lut (.I0(n48831), .I1(n2_adj_5057), .I2(n1752), 
            .I3(n38489), .O(encoder0_position_scaled_23__N_34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_18 (.CI(n38489), .I0(n2_adj_5057), .I1(n1752), .CO(n38490));
    SB_LUT4 add_1944_17_lut (.I0(n48859), .I1(n2_adj_5057), .I2(n1851), 
            .I3(n38488), .O(encoder0_position_scaled_23__N_34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_17 (.CI(n38488), .I0(n2_adj_5057), .I1(n1851), .CO(n38489));
    SB_LUT4 add_29_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n37174), .O(n676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1944_16_lut (.I0(n49096), .I1(n2_adj_5057), .I2(n1950), 
            .I3(n38487), .O(encoder0_position_scaled_23__N_34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n38226), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1944_16 (.CI(n38487), .I0(n2_adj_5057), .I1(n1950), .CO(n38488));
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n38084), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_700_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_5040));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_1944_15_lut (.I0(n49129), .I1(n2_adj_5057), .I2(n2049), 
            .I3(n38486), .O(encoder0_position_scaled_23__N_34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_15 (.CI(n38486), .I0(n2_adj_5057), .I1(n2049), .CO(n38487));
    SB_LUT4 add_1944_14_lut (.I0(n49153), .I1(n2_adj_5057), .I2(n2148), 
            .I3(n38485), .O(encoder0_position_scaled_23__N_34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_14 (.CI(n38485), .I0(n2_adj_5057), .I1(n2148), .CO(n38486));
    SB_LUT4 add_1944_13_lut (.I0(n49181), .I1(n2_adj_5057), .I2(n2247), 
            .I3(n38484), .O(encoder0_position_scaled_23__N_34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_13 (.CI(n38484), .I0(n2_adj_5057), .I1(n2247), .CO(n38485));
    SB_LUT4 add_1944_12_lut (.I0(n49207), .I1(n2_adj_5057), .I2(n2346), 
            .I3(n38483), .O(encoder0_position_scaled_23__N_34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_12 (.CI(n38483), .I0(n2_adj_5057), .I1(n2346), .CO(n38484));
    SB_LUT4 add_1944_11_lut (.I0(n49231), .I1(n2_adj_5057), .I2(n2445), 
            .I3(n38482), .O(encoder0_position_scaled_23__N_34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_11 (.CI(n38482), .I0(n2_adj_5057), .I1(n2445), .CO(n38483));
    SB_LUT4 add_1944_10_lut (.I0(n48562), .I1(n2_adj_5057), .I2(n2544), 
            .I3(n38481), .O(encoder0_position_scaled_23__N_34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_10 (.CI(n38481), .I0(n2_adj_5057), .I1(n2544), .CO(n38482));
    SB_LUT4 add_1944_9_lut (.I0(n48618), .I1(n2_adj_5057), .I2(n2643), 
            .I3(n38480), .O(encoder0_position_scaled_23__N_34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_9 (.CI(n38480), .I0(n2_adj_5057), .I1(n2643), .CO(n38481));
    SB_CARRY add_29_16 (.CI(n37174), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n37175));
    SB_LUT4 add_1944_8_lut (.I0(n48904), .I1(n2_adj_5057), .I2(n2742), 
            .I3(n38479), .O(encoder0_position_scaled_23__N_34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_8 (.CI(n38479), .I0(n2_adj_5057), .I1(n2742), .CO(n38480));
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n38084), .I0(n2221), 
            .I1(VCC_net), .CO(n38085));
    SB_LUT4 add_1944_7_lut (.I0(n48936), .I1(n2_adj_5057), .I2(n2841), 
            .I3(n38478), .O(encoder0_position_scaled_23__N_34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_29_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n37173), .O(n677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1944_7 (.CI(n38478), .I0(n2_adj_5057), .I1(n2841), .CO(n38479));
    SB_CARRY add_78_10 (.CI(n37199), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n37200));
    SB_LUT4 add_1944_6_lut (.I0(n48968), .I1(n2_adj_5057), .I2(n2940), 
            .I3(n38477), .O(encoder0_position_scaled_23__N_34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_6 (.CI(n38477), .I0(n2_adj_5057), .I1(n2940), .CO(n38478));
    SB_LUT4 add_1944_5_lut (.I0(n49002), .I1(n2_adj_5057), .I2(n3039), 
            .I3(n38476), .O(encoder0_position_scaled_23__N_34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_5 (.CI(n38476), .I0(n2_adj_5057), .I1(n3039), .CO(n38477));
    SB_LUT4 add_1944_4_lut (.I0(n49036), .I1(n2_adj_5057), .I2(n3138), 
            .I3(n38475), .O(encoder0_position_scaled_23__N_34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1944_4 (.CI(n38475), .I0(n2_adj_5057), .I1(n3138), .CO(n38476));
    SB_LUT4 add_1944_3_lut (.I0(n49040), .I1(n2_adj_5057), .I2(n3237), 
            .I3(n38474), .O(encoder0_position_scaled_23__N_34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n38083), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15409_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n42229), 
            .I3(GND_net), .O(n28468));   // verilog/coms.v(127[12] 300[6])
    defparam i15409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15410_3_lut (.I0(\data_in_frame[0] [2]), .I1(rx_data[2]), .I2(n42229), 
            .I3(GND_net), .O(n28469));   // verilog/coms.v(127[12] 300[6])
    defparam i15410_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n38226), .I0(n2316), 
            .I1(VCC_net), .CO(n38227));
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n38083), .I0(n2222), 
            .I1(VCC_net), .CO(n38084));
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n648), 
            .I1(GND_net), .CO(n38359));
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n38225), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_15 (.CI(n37173), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n37174));
    SB_LUT4 add_29_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n37172), .O(n678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1944_3 (.CI(n38474), .I0(n2_adj_5057), .I1(n3237), .CO(n38475));
    SB_LUT4 i15411_3_lut (.I0(\data_in_frame[0] [1]), .I1(rx_data[1]), .I2(n42229), 
            .I3(GND_net), .O(n28470));   // verilog/coms.v(127[12] 300[6])
    defparam i15411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n48936), .I1(n2808), 
            .I2(VCC_net), .I3(n38358), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1944_2_lut (.I0(n49074), .I1(n2_adj_5057), .I2(n34679), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_34[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1944_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n38082), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1944_2 (.CI(VCC_net), .I0(n2_adj_5057), .I1(n34679), 
            .CO(n38474));
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n38225), .I0(n2317), 
            .I1(VCC_net), .CO(n38226));
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n38357), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n38224), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15412_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n27753), .I3(GND_net), .O(n28471));   // verilog/coms.v(127[12] 300[6])
    defparam i15412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n38357), .I0(n2809), 
            .I1(VCC_net), .CO(n38358));
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n38224), .I0(n2318), 
            .I1(VCC_net), .CO(n38225));
    SB_CARRY add_29_6 (.CI(n37164), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n37165));
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n38082), .I0(n2223), 
            .I1(VCC_net), .CO(n38083));
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n38356), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15413_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n27753), .I3(GND_net), .O(n28472));   // verilog/coms.v(127[12] 300[6])
    defparam i15413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(n49040), .I1(n3204), 
            .I2(VCC_net), .I3(n38473), .O(n46486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n38472), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n38356), .I0(n2810), 
            .I1(VCC_net), .CO(n38357));
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n38223), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n38081), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_700_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_5036));   // verilog/pwm.v(21[8:24])
    defparam LessThan_700_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32773_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n47726));
    defparam i32773_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15414_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n27753), .I3(GND_net), .O(n28473));   // verilog/coms.v(127[12] 300[6])
    defparam i15414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15415_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n27753), .I3(GND_net), .O(n28474));   // verilog/coms.v(127[12] 300[6])
    defparam i15415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15416_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n27753), .I3(GND_net), .O(n28475));   // verilog/coms.v(127[12] 300[6])
    defparam i15416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15417_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n27753), .I3(GND_net), .O(n28476));   // verilog/coms.v(127[12] 300[6])
    defparam i15417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15418_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n27753), .I3(GND_net), .O(n28477));   // verilog/coms.v(127[12] 300[6])
    defparam i15418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n38355), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n38223), .I0(n2319), 
            .I1(VCC_net), .CO(n38224));
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n38081), .I0(n2224), 
            .I1(VCC_net), .CO(n38082));
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n38472), .I0(n3205), 
            .I1(VCC_net), .CO(n38473));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n38080), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n38222), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_14 (.CI(n37172), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n37173));
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n38080), .I0(n2225), 
            .I1(VCC_net), .CO(n38081));
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n38471), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15419_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n27753), .I3(GND_net), .O(n28478));   // verilog/coms.v(127[12] 300[6])
    defparam i15419_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n38471), .I0(n3206), 
            .I1(VCC_net), .CO(n38472));
    SB_LUT4 i15420_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n27753), .I3(GND_net), .O(n28479));   // verilog/coms.v(127[12] 300[6])
    defparam i15420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15421_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n27753), .I3(GND_net), .O(n28480));   // verilog/coms.v(127[12] 300[6])
    defparam i15421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15422_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n27753), .I3(GND_net), .O(n28481));   // verilog/coms.v(127[12] 300[6])
    defparam i15422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15423_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n27753), .I3(GND_net), .O(n28482));   // verilog/coms.v(127[12] 300[6])
    defparam i15423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15424_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n27753), .I3(GND_net), .O(n28483));   // verilog/coms.v(127[12] 300[6])
    defparam i15424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15425_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n27753), .I3(GND_net), .O(n28484));   // verilog/coms.v(127[12] 300[6])
    defparam i15425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15426_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n27753), .I3(GND_net), .O(n28485));   // verilog/coms.v(127[12] 300[6])
    defparam i15426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21484_3_lut (.I0(n639), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n34533));
    defparam i21484_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15427_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n27753), .I3(GND_net), .O(n28486));   // verilog/coms.v(127[12] 300[6])
    defparam i15427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15428_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n27753), .I3(GND_net), .O(n28487));   // verilog/coms.v(127[12] 300[6])
    defparam i15428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15429_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n27753), .I3(GND_net), .O(n28488));   // verilog/coms.v(127[12] 300[6])
    defparam i15429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15430_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n27753), .I3(GND_net), .O(n28489));   // verilog/coms.v(127[12] 300[6])
    defparam i15430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15431_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n27753), .I3(GND_net), .O(n28490));   // verilog/coms.v(127[12] 300[6])
    defparam i15431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15432_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n27753), .I3(GND_net), .O(n28491));   // verilog/coms.v(127[12] 300[6])
    defparam i15432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15433_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n27753), .I3(GND_net), .O(n28492));   // verilog/coms.v(127[12] 300[6])
    defparam i15433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15434_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n27753), .I3(GND_net), .O(n28493));   // verilog/coms.v(127[12] 300[6])
    defparam i15434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15435_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n23943), .I3(GND_net), .O(n28494));   // verilog/coms.v(127[12] 300[6])
    defparam i15435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n1927), .I1(n1926), .I2(n1925), .I3(n1928), 
            .O(n45082));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1817 (.I0(n2026), .I1(n2027), .I2(GND_net), .I3(GND_net), 
            .O(n45392));
    defparam i1_2_lut_adj_1817.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n2025), .I1(n45392), .I2(n2024), .I3(n2028), 
            .O(n45396));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hfffe;
    SB_LUT4 i15436_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n23943), .I3(GND_net), .O(n28495));   // verilog/coms.v(127[12] 300[6])
    defparam i15436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15437_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n23943), .I3(GND_net), .O(n28496));   // verilog/coms.v(127[12] 300[6])
    defparam i15437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15438_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n23943), .I3(GND_net), .O(n28497));   // verilog/coms.v(127[12] 300[6])
    defparam i15438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15439_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n23943), .I3(GND_net), .O(n28498));   // verilog/coms.v(127[12] 300[6])
    defparam i15439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15440_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n23943), .I3(GND_net), .O(n28499));   // verilog/coms.v(127[12] 300[6])
    defparam i15440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15441_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n23943), .I3(GND_net), .O(n28500));   // verilog/coms.v(127[12] 300[6])
    defparam i15441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15442_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n23943), .I3(GND_net), .O(n28501));   // verilog/coms.v(127[12] 300[6])
    defparam i15442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15443_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n23943), .I3(GND_net), .O(n28502));   // verilog/coms.v(127[12] 300[6])
    defparam i15443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15444_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n23943), .I3(GND_net), .O(n28503));   // verilog/coms.v(127[12] 300[6])
    defparam i15444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15445_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n23943), .I3(GND_net), .O(n28504));   // verilog/coms.v(127[12] 300[6])
    defparam i15445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15446_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n23943), .I3(GND_net), .O(n28505));   // verilog/coms.v(127[12] 300[6])
    defparam i15446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15447_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n23943), .I3(GND_net), .O(n28506));   // verilog/coms.v(127[12] 300[6])
    defparam i15447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15104_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n2380), .I3(GND_net), .O(n28163));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15105_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n27752), .I3(GND_net), .O(n28164));   // verilog/coms.v(127[12] 300[6])
    defparam i15105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15106_4_lut (.I0(state_7__N_4003[3]), .I1(data[7]), .I2(n33700), 
            .I3(n26657), .O(n28165));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15106_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15107_4_lut (.I0(state_7__N_4003[3]), .I1(data[6]), .I2(n33700), 
            .I3(n26652), .O(n28166));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15107_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15108_4_lut (.I0(state_7__N_4003[3]), .I1(data[5]), .I2(n4_adj_4981), 
            .I3(n26657), .O(n28167));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15108_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15109_4_lut (.I0(state_7__N_4003[3]), .I1(data[4]), .I2(n4_adj_4981), 
            .I3(n26652), .O(n28168));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15109_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15110_4_lut (.I0(state_7__N_4003[3]), .I1(data[3]), .I2(n4_adj_4980), 
            .I3(n26657), .O(n28169));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15110_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15111_4_lut (.I0(state_7__N_4003[3]), .I1(data[2]), .I2(n4_adj_4980), 
            .I3(n26652), .O(n28170));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15111_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15448_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n23943), .I3(GND_net), .O(n28507));   // verilog/coms.v(127[12] 300[6])
    defparam i15448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15449_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n23943), .I3(GND_net), .O(n28508));   // verilog/coms.v(127[12] 300[6])
    defparam i15449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15450_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n23943), .I3(GND_net), .O(n28509));   // verilog/coms.v(127[12] 300[6])
    defparam i15450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15451_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n23943), .I3(GND_net), .O(n28510));   // verilog/coms.v(127[12] 300[6])
    defparam i15451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15452_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n23943), .I3(GND_net), .O(n28511));   // verilog/coms.v(127[12] 300[6])
    defparam i15452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15453_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n23943), .I3(GND_net), .O(n28512));   // verilog/coms.v(127[12] 300[6])
    defparam i15453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15454_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n23943), .I3(GND_net), .O(n28513));   // verilog/coms.v(127[12] 300[6])
    defparam i15454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15115_4_lut (.I0(state_7__N_4003[3]), .I1(data[1]), .I2(n10_adj_5097), 
            .I3(n26657), .O(n28174));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15115_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15117_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5009), 
            .I3(n26628), .O(n28176));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15117_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15118_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4984), 
            .I3(n26633), .O(n28177));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15118_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15455_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n23943), .I3(GND_net), .O(n28514));   // verilog/coms.v(127[12] 300[6])
    defparam i15455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15456_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n23943), .I3(GND_net), .O(n28515));   // verilog/coms.v(127[12] 300[6])
    defparam i15456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15457_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n23943), .I3(GND_net), .O(n28516));   // verilog/coms.v(127[12] 300[6])
    defparam i15457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15458_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n23943), .I3(GND_net), .O(n28517));   // verilog/coms.v(127[12] 300[6])
    defparam i15458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15459_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n23943), .I3(GND_net), .O(n28518));   // verilog/coms.v(127[12] 300[6])
    defparam i15459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15460_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n23943), .I3(GND_net), .O(n28519));   // verilog/coms.v(127[12] 300[6])
    defparam i15460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15461_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n23943), .I3(GND_net), .O(n28520));   // verilog/coms.v(127[12] 300[6])
    defparam i15461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21318_3_lut (.I0(n638), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n34363));
    defparam i21318_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15462_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n23943), .I3(GND_net), .O(n28521));   // verilog/coms.v(127[12] 300[6])
    defparam i15462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15463_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n23943), .I3(GND_net), .O(n28522));   // verilog/coms.v(127[12] 300[6])
    defparam i15463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15464_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n23943), .I3(GND_net), .O(n28523));   // verilog/coms.v(127[12] 300[6])
    defparam i15464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(n1922), .I1(n1923), .I2(n45082), .I3(n1924), 
            .O(n45088));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 i15465_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n23943), .I3(GND_net), .O(n28524));   // verilog/coms.v(127[12] 300[6])
    defparam i15465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1820 (.I0(n1929), .I1(n34363), .I2(n1930), .I3(n1931), 
            .O(n43181));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'ha080;
    SB_LUT4 i17137_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n23943), .I3(GND_net), .O(n28525));
    defparam i17137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15467_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n23943), .I3(GND_net), .O(n28526));   // verilog/coms.v(127[12] 300[6])
    defparam i15467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15468_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n23943), .I3(GND_net), .O(n28527));   // verilog/coms.v(127[12] 300[6])
    defparam i15468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15469_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n23943), .I3(GND_net), .O(n28528));   // verilog/coms.v(127[12] 300[6])
    defparam i15469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15470_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n23943), .I3(GND_net), .O(n28529));   // verilog/coms.v(127[12] 300[6])
    defparam i15470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15471_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n23943), .I3(GND_net), .O(n28530));   // verilog/coms.v(127[12] 300[6])
    defparam i15471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15472_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n23943), .I3(GND_net), .O(n28531));   // verilog/coms.v(127[12] 300[6])
    defparam i15472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15473_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n23943), .I3(GND_net), .O(n28532));   // verilog/coms.v(127[12] 300[6])
    defparam i15473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15474_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n23943), .I3(GND_net), .O(n28533));   // verilog/coms.v(127[12] 300[6])
    defparam i15474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15475_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n23943), .I3(GND_net), .O(n28534));   // verilog/coms.v(127[12] 300[6])
    defparam i15475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15476_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n23943), .I3(GND_net), .O(n28535));   // verilog/coms.v(127[12] 300[6])
    defparam i15476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15477_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n23943), .I3(GND_net), .O(n28536));   // verilog/coms.v(127[12] 300[6])
    defparam i15477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15478_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n23943), .I3(GND_net), .O(n28537));   // verilog/coms.v(127[12] 300[6])
    defparam i15478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15479_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n23943), .I3(GND_net), .O(n28538));   // verilog/coms.v(127[12] 300[6])
    defparam i15479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15480_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n23943), .I3(GND_net), .O(n28539));   // verilog/coms.v(127[12] 300[6])
    defparam i15480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15482_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n23943), .I3(GND_net), .O(n28541));   // verilog/coms.v(127[12] 300[6])
    defparam i15482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15483_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n23943), 
            .I3(GND_net), .O(n28542));   // verilog/coms.v(127[12] 300[6])
    defparam i15483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15484_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n23943), 
            .I3(GND_net), .O(n28543));   // verilog/coms.v(127[12] 300[6])
    defparam i15484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15485_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n23943), 
            .I3(GND_net), .O(n28544));   // verilog/coms.v(127[12] 300[6])
    defparam i15485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15486_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n23943), 
            .I3(GND_net), .O(n28545));   // verilog/coms.v(127[12] 300[6])
    defparam i15486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15487_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n23943), 
            .I3(GND_net), .O(n28546));   // verilog/coms.v(127[12] 300[6])
    defparam i15487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15488_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n23943), 
            .I3(GND_net), .O(n28547));   // verilog/coms.v(127[12] 300[6])
    defparam i15488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15489_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n23943), 
            .I3(GND_net), .O(n28548));   // verilog/coms.v(127[12] 300[6])
    defparam i15489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15490_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n23943), 
            .I3(GND_net), .O(n28549));   // verilog/coms.v(127[12] 300[6])
    defparam i15490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17127_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n23943), 
            .I3(GND_net), .O(n28550));
    defparam i17127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15492_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n23943), 
            .I3(GND_net), .O(n28551));   // verilog/coms.v(127[12] 300[6])
    defparam i15492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15493_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n23943), 
            .I3(GND_net), .O(n28552));   // verilog/coms.v(127[12] 300[6])
    defparam i15493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15494_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n23943), 
            .I3(GND_net), .O(n28553));   // verilog/coms.v(127[12] 300[6])
    defparam i15494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15495_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n23943), 
            .I3(GND_net), .O(n28554));   // verilog/coms.v(127[12] 300[6])
    defparam i15495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15496_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n23943), 
            .I3(GND_net), .O(n28555));   // verilog/coms.v(127[12] 300[6])
    defparam i15496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1821 (.I0(n2029), .I1(n34533), .I2(n2030), .I3(n2031), 
            .O(n43217));
    defparam i1_4_lut_adj_1821.LUT_INIT = 16'ha080;
    SB_LUT4 i15497_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n23943), 
            .I3(GND_net), .O(n28556));   // verilog/coms.v(127[12] 300[6])
    defparam i15497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1822 (.I0(n1920), .I1(n43181), .I2(n1921), .I3(n45088), 
            .O(n45094));
    defparam i1_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_LUT4 i15498_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n23943), 
            .I3(GND_net), .O(n28557));   // verilog/coms.v(127[12] 300[6])
    defparam i15498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34149_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n45094), 
            .O(n1950));
    defparam i34149_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15499_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n23943), 
            .I3(GND_net), .O(n28558));   // verilog/coms.v(127[12] 300[6])
    defparam i15499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15500_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n23943), 
            .I3(GND_net), .O(n28559));   // verilog/coms.v(127[12] 300[6])
    defparam i15500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15501_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n23943), 
            .I3(GND_net), .O(n28560));   // verilog/coms.v(127[12] 300[6])
    defparam i15501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15502_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n23943), 
            .I3(GND_net), .O(n28561));   // verilog/coms.v(127[12] 300[6])
    defparam i15502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15503_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n23943), 
            .I3(GND_net), .O(n28562));   // verilog/coms.v(127[12] 300[6])
    defparam i15503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15504_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n23943), 
            .I3(GND_net), .O(n28563));   // verilog/coms.v(127[12] 300[6])
    defparam i15504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15505_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n23943), 
            .I3(GND_net), .O(n28564));   // verilog/coms.v(127[12] 300[6])
    defparam i15505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15506_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n23943), 
            .I3(GND_net), .O(n28565));   // verilog/coms.v(127[12] 300[6])
    defparam i15506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15507_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n23943), .I3(GND_net), .O(n28566));   // verilog/coms.v(127[12] 300[6])
    defparam i15507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15508_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n23943), .I3(GND_net), .O(n28567));   // verilog/coms.v(127[12] 300[6])
    defparam i15508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15509_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n23943), .I3(GND_net), .O(n28568));   // verilog/coms.v(127[12] 300[6])
    defparam i15509_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.\a_new[1] (a_new[1]), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1188(CLK_c), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .b_prev(b_prev), .n28221(n28221), .n1152(n1152), .direction_N_3807(direction_N_3807), 
            .encoder0_position({encoder0_position}), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(187[57] 194[6])
    SB_LUT4 i15510_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n23943), .I3(GND_net), .O(n28569));   // verilog/coms.v(127[12] 300[6])
    defparam i15510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15511_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n23943), .I3(GND_net), .O(n28570));   // verilog/coms.v(127[12] 300[6])
    defparam i15511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n45396), 
            .O(n45402));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 i15512_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n23943), .I3(GND_net), .O(n28571));   // verilog/coms.v(127[12] 300[6])
    defparam i15512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15513_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n23943), .I3(GND_net), .O(n28572));   // verilog/coms.v(127[12] 300[6])
    defparam i15513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15514_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n23943), .I3(GND_net), .O(n28573));   // verilog/coms.v(127[12] 300[6])
    defparam i15514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15515_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n23943), .I3(GND_net), .O(n28574));   // verilog/coms.v(127[12] 300[6])
    defparam i15515_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 i15516_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n23943), .I3(GND_net), .O(n28575));   // verilog/coms.v(127[12] 300[6])
    defparam i15516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15517_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n23943), .I3(GND_net), .O(n28576));   // verilog/coms.v(127[12] 300[6])
    defparam i15517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1383_rep_34_3_lut (.I0(n2095), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n46578));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1383_rep_34_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15518_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n23943), .I3(GND_net), .O(n28577));   // verilog/coms.v(127[12] 300[6])
    defparam i15518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15519_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n23943), .I3(GND_net), .O(n28578));   // verilog/coms.v(127[12] 300[6])
    defparam i15519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15520_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n23943), .I3(GND_net), .O(n28579));   // verilog/coms.v(127[12] 300[6])
    defparam i15520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15165_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5009), 
            .I3(n26633), .O(n28224));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15165_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i274_2_lut (.I0(n777), .I1(n26487), .I2(GND_net), .I3(GND_net), 
            .O(n1419));   // verilog/TinyFPGA_B.v(278[9] 284[12])
    defparam i274_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4948));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15521_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n23943), .I3(GND_net), .O(n28580));   // verilog/coms.v(127[12] 300[6])
    defparam i15521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32795_4_lut (.I0(n5_adj_5017), .I1(n6_adj_5030), .I2(n5855), 
            .I3(n1419), .O(n47573));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i32795_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 i49_4_lut (.I0(n47573), .I1(data_ready), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n5855), .O(n41391));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i49_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_1824 (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_4977), .I3(control_mode[2]), .O(n26489));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam i1_2_lut_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26487), .I3(GND_net), .O(n5722));
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1825 (.I0(n2019), .I1(n2020), .I2(n45402), .I3(n43217), 
            .O(n45408));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32775_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n47518));
    defparam i32775_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26487), .I3(GND_net), .O(n26488));   // verilog/TinyFPGA_B.v(277[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5161[1]), .I1(r_SM_Main_adj_5161[0]), 
            .I2(r_SM_Main_adj_5161[2]), .I3(r_SM_Main_2__N_3513[1]), .O(n49552));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15173_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n2380), .I3(GND_net), .O(n28232));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15174_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n2380), .I3(GND_net), .O(n28233));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15175_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n2380), .I3(GND_net), .O(n28234));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15176_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n2380), .I3(GND_net), .O(n28235));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15177_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n2380), .I3(GND_net), .O(n28236));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15178_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n2380), .I3(GND_net), .O(n28237));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15179_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n2380), .I3(GND_net), .O(n28238));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15180_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n2380), .I3(GND_net), .O(n28239));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15181_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n2380), .I3(GND_net), .O(n28240));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15182_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n2380), .I3(GND_net), .O(n28241));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15183_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n2380), .I3(GND_net), .O(n28242));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15522_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n23943), .I3(GND_net), .O(n28581));   // verilog/coms.v(127[12] 300[6])
    defparam i15522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15184_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n2380), .I3(GND_net), .O(n28243));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15185_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n2380), .I3(GND_net), .O(n28244));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15186_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n2380), .I3(GND_net), .O(n28245));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4973));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4972));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4971));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4970));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4969));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4968));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4967));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4966));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4965));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4964));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4963));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4962));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4961));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15187_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n2380), .I3(GND_net), .O(n28246));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4960));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4959));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4958));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4957));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4956));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4955));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4954));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4953));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder0_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5005));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5004));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder0_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder1_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15119_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4984), 
            .I3(n26628), .O(n28178));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15119_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15188_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n2380), .I3(GND_net), .O(n28247));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34179_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n45408), 
            .O(n2049));
    defparam i34179_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_3_lut_adj_1826 (.I0(n2125), .I1(n2124), .I2(n2127), .I3(GND_net), 
            .O(n45240));
    defparam i1_3_lut_adj_1826.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1827 (.I0(n2123), .I1(n2128), .I2(n2126), .I3(GND_net), 
            .O(n45242));
    defparam i1_3_lut_adj_1827.LUT_INIT = 16'hfefe;
    SB_LUT4 i21584_4_lut (.I0(n640), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n34637));
    defparam i21584_4_lut.LUT_INIT = 16'hfcec;
    motorControl control (.PWMLimit({PWMLimit}), .GND_net(GND_net), .\Ki[8] (Ki[8]), 
            .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), 
            .\Kp[2] (Kp[2]), .\Ki[4] (Ki[4]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), 
            .\Ki[5] (Ki[5]), .\Kp[6] (Kp[6]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), 
            .\Ki[9] (Ki[9]), .\Kp[7] (Kp[7]), .\Kp[3] (Kp[3]), .\Kp[8] (Kp[8]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[9] (Kp[9]), .\Ki[10] (Ki[10]), 
            .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .setpoint({setpoint}), .motor_state({motor_state}), 
            .\Kp[15] (Kp[15]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), 
            .duty({duty}), .clk32MHz(clk32MHz), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), 
            .IntegralLimit({IntegralLimit}), .VCC_net(VCC_net), .n49248(n49248)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(173[16] 185[4])
    SB_LUT4 i1_4_lut_adj_1828 (.I0(n2121), .I1(n2122), .I2(n45242), .I3(n45240), 
            .O(n45248));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n2129), .I1(n45248), .I2(n34637), .I3(n2130), 
            .O(n45250));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'heccc;
    \quadrature_decoder(1,500000)  quad_counter1 (.\a_new[1] (a_new_adj_5130[1]), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1188(CLK_c), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .b_prev(b_prev_adj_5011), .n28216(n28216), .n1193(n1193), 
            .direction_N_3807(direction_N_3807_adj_5012), .encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(196[57] 203[6])
    coms neopxl_color_23__I_0 (.CLK_c(CLK_c), .n28292(n28292), .control_mode({control_mode}), 
         .n28291(n28291), .n28290(n28290), .n28289(n28289), .n28288(n28288), 
         .GND_net(GND_net), .\data_in_frame[3] ({\data_in_frame[3] }), .n28287(n28287), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .n28286(n28286), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .n28285(n28285), .PWMLimit({PWMLimit}), .n28284(n28284), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .n23943(n23943), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .byte_transmit_counter({Open_0, Open_1, Open_2, Open_3, Open_4, 
         byte_transmit_counter[2:1], Open_5}), .n28283(n28283), .n28282(n28282), 
         .n28281(n28281), .n28280(n28280), .\data_in_frame[0] ({\data_in_frame[0] }), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n28279(n28279), .n28278(n28278), .n28277(n28277), .n28276(n28276), 
         .rx_data_ready(rx_data_ready), .setpoint({setpoint}), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n28275(n28275), .n28274(n28274), .\data_in[3] ({\data_in[3] }), 
         .\data_in[1] ({\data_in[1] }), .\data_in[0] ({\data_in[0] }), .\data_in[2] ({\data_in[2] }), 
         .n28273(n28273), .n28272(n28272), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .\byte_transmit_counter[0] (byte_transmit_counter[0]), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .n28271(n28271), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n28270(n28270), 
         .n28269(n28269), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n28268(n28268), 
         .n28267(n28267), .n28266(n28266), .n28265(n28265), .n28264(n28264), 
         .n28263(n28263), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] [7], 
         Open_6, \data_out_frame[18] [5:2], Open_7, \data_out_frame[18] [0]}), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .DE_c(DE_c), .tx_active(tx_active), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .n49368(n49368), .n46660(n46660), .ID({ID}), .n43603(n43603), 
         .n42551(n42551), .n27752(n27752), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n47614(n47614), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .n42541(n42541), .n42790(n42790), .LED_c(LED_c), .n49422(n49422), 
         .n28189(n28189), .n43610(n43610), .n27554(n27554), .n28188(n28188), 
         .n42897(n42897), .\data_out_frame[18][6] (\data_out_frame[18] [6]), 
         .n40598(n40598), .n28187(n28187), .n28186(n28186), .neopxl_color({neopxl_color}), 
         .n28185(n28185), .\Ki[0] (Ki[0]), .n28184(n28184), .\Kp[0] (Kp[0]), 
         .n28183(n28183), .n28738(n28738), .IntegralLimit({IntegralLimit}), 
         .n28737(n28737), .n28736(n28736), .n28735(n28735), .n28734(n28734), 
         .n28733(n28733), .n28732(n28732), .n28731(n28731), .n28730(n28730), 
         .n28729(n28729), .n28728(n28728), .n28727(n28727), .n28726(n28726), 
         .n28725(n28725), .n28724(n28724), .n28723(n28723), .n28722(n28722), 
         .n28721(n28721), .n28720(n28720), .n28719(n28719), .n28718(n28718), 
         .n28717(n28717), .n28716(n28716), .n28715(n28715), .n28714(n28714), 
         .n28713(n28713), .n28712(n28712), .n28711(n28711), .n28710(n28710), 
         .n28709(n28709), .n28708(n28708), .n28707(n28707), .n28706(n28706), 
         .n28705(n28705), .n28704(n28704), .n28703(n28703), .n28702(n28702), 
         .n28701(n28701), .n28700(n28700), .n28698(n28698), .n28697(n28697), 
         .n28696(n28696), .n28695(n28695), .n28694(n28694), .n28693(n28693), 
         .n28692(n28692), .n28691(n28691), .n28690(n28690), .n28689(n28689), 
         .n28688(n28688), .n28687(n28687), .n28686(n28686), .n28685(n28685), 
         .n28684(n28684), .n28683(n28683), .\Kp[1] (Kp[1]), .n28682(n28682), 
         .\Kp[2] (Kp[2]), .n28681(n28681), .\Kp[3] (Kp[3]), .n28680(n28680), 
         .\Kp[4] (Kp[4]), .n28679(n28679), .\Kp[5] (Kp[5]), .n28678(n28678), 
         .\Kp[6] (Kp[6]), .n28677(n28677), .\Kp[7] (Kp[7]), .n28676(n28676), 
         .\Kp[8] (Kp[8]), .n28675(n28675), .\Kp[9] (Kp[9]), .n28674(n28674), 
         .\Kp[10] (Kp[10]), .n28673(n28673), .\Kp[11] (Kp[11]), .n28672(n28672), 
         .\Kp[12] (Kp[12]), .n28671(n28671), .\Kp[13] (Kp[13]), .n28670(n28670), 
         .\Kp[14] (Kp[14]), .n28669(n28669), .\Kp[15] (Kp[15]), .n28668(n28668), 
         .\Ki[1] (Ki[1]), .n28667(n28667), .\Ki[2] (Ki[2]), .n28666(n28666), 
         .\Ki[3] (Ki[3]), .n28665(n28665), .\Ki[4] (Ki[4]), .n28664(n28664), 
         .\Ki[5] (Ki[5]), .n28663(n28663), .\Ki[6] (Ki[6]), .n28662(n28662), 
         .\Ki[7] (Ki[7]), .n28661(n28661), .\Ki[8] (Ki[8]), .n28660(n28660), 
         .\Ki[9] (Ki[9]), .n28659(n28659), .\Ki[10] (Ki[10]), .n28658(n28658), 
         .\Ki[11] (Ki[11]), .n28657(n28657), .\Ki[12] (Ki[12]), .n28656(n28656), 
         .\Ki[13] (Ki[13]), .n28655(n28655), .\Ki[14] (Ki[14]), .n28654(n28654), 
         .\Ki[15] (Ki[15]), .n28653(n28653), .n28652(n28652), .n28651(n28651), 
         .n28650(n28650), .n28649(n28649), .n28648(n28648), .n28647(n28647), 
         .n28646(n28646), .n28645(n28645), .n28644(n28644), .n28643(n28643), 
         .n28642(n28642), .n28641(n28641), .n28640(n28640), .n28639(n28639), 
         .n28638(n28638), .n28637(n28637), .n28636(n28636), .n28635(n28635), 
         .n28634(n28634), .n28633(n28633), .n28632(n28632), .n28631(n28631), 
         .n28630(n28630), .n28629(n28629), .n28628(n28628), .n28627(n28627), 
         .n28626(n28626), .n28625(n28625), .n28624(n28624), .n28623(n28623), 
         .n28622(n28622), .n28621(n28621), .n28620(n28620), .n28619(n28619), 
         .n28618(n28618), .n28617(n28617), .n28616(n28616), .n28615(n28615), 
         .n28614(n28614), .n28613(n28613), .n28612(n28612), .n28611(n28611), 
         .n28610(n28610), .n28609(n28609), .n28608(n28608), .n28607(n28607), 
         .n28606(n28606), .n28605(n28605), .n28604(n28604), .n28603(n28603), 
         .n28602(n28602), .n28601(n28601), .n28600(n28600), .n28599(n28599), 
         .n28598(n28598), .n28597(n28597), .n28596(n28596), .n28595(n28595), 
         .n28594(n28594), .n28593(n28593), .n28592(n28592), .n28591(n28591), 
         .n28590(n28590), .n28589(n28589), .n28588(n28588), .n28587(n28587), 
         .n28586(n28586), .n28585(n28585), .n28584(n28584), .n28583(n28583), 
         .n28582(n28582), .rx_data({rx_data}), .n28581(n28581), .n28580(n28580), 
         .n28579(n28579), .n28578(n28578), .n28577(n28577), .n28576(n28576), 
         .n28575(n28575), .n28574(n28574), .n28573(n28573), .n28572(n28572), 
         .n28571(n28571), .n28570(n28570), .n28569(n28569), .n28568(n28568), 
         .n28567(n28567), .n28566(n28566), .n28565(n28565), .n28564(n28564), 
         .n28563(n28563), .n28562(n28562), .n28561(n28561), .n28560(n28560), 
         .n28559(n28559), .n28558(n28558), .n28557(n28557), .n28556(n28556), 
         .n28555(n28555), .n28554(n28554), .n28553(n28553), .n28552(n28552), 
         .n28551(n28551), .n28550(n28550), .n28549(n28549), .n28548(n28548), 
         .n28547(n28547), .n28546(n28546), .n28545(n28545), .n28544(n28544), 
         .n28543(n28543), .n28542(n28542), .n28541(n28541), .n28539(n28539), 
         .n28538(n28538), .n28537(n28537), .n28536(n28536), .n28535(n28535), 
         .n28534(n28534), .n28533(n28533), .n28532(n28532), .n28531(n28531), 
         .n28530(n28530), .n28529(n28529), .n28528(n28528), .n28527(n28527), 
         .n28526(n28526), .n28525(n28525), .n28524(n28524), .n28523(n28523), 
         .n28522(n28522), .n28521(n28521), .n28520(n28520), .n28519(n28519), 
         .n28518(n28518), .n28517(n28517), .n28516(n28516), .n28515(n28515), 
         .n28514(n28514), .n28513(n28513), .n28512(n28512), .n28511(n28511), 
         .n28510(n28510), .n28509(n28509), .n28508(n28508), .n28507(n28507), 
         .n28164(n28164), .n28506(n28506), .n28505(n28505), .n28504(n28504), 
         .n28503(n28503), .n28502(n28502), .n28501(n28501), .n28500(n28500), 
         .n28499(n28499), .n28498(n28498), .n28497(n28497), .n28496(n28496), 
         .n28495(n28495), .n28494(n28494), .n28493(n28493), .n28492(n28492), 
         .n28491(n28491), .n28490(n28490), .n28489(n28489), .n28488(n28488), 
         .n28487(n28487), .n28486(n28486), .n28485(n28485), .n28484(n28484), 
         .n28483(n28483), .n28482(n28482), .n28481(n28481), .n28480(n28480), 
         .n28479(n28479), .n28478(n28478), .n28477(n28477), .n28476(n28476), 
         .n28475(n28475), .n28474(n28474), .n28473(n28473), .n28472(n28472), 
         .n28471(n28471), .n28470(n28470), .n28469(n28469), .n28468(n28468), 
         .n28467(n28467), .n28466(n28466), .n28465(n28465), .n28464(n28464), 
         .n28405(n28405), .n28403(n28403), .n28402(n28402), .n28401(n28401), 
         .n28400(n28400), .n28399(n28399), .n28398(n28398), .n28397(n28397), 
         .n4(n4_adj_5028), .\state[0] (state_adj_5170[0]), .\state[2] (state_adj_5170[2]), 
         .\state[3] (state_adj_5170[3]), .n6014(n6014), .\displacement[17] (displacement[17]), 
         .n27753(n27753), .n42230(n42230), .n42229(n42229), .\r_SM_Main_2__N_3513[1] (r_SM_Main_2__N_3513[1]), 
         .r_SM_Main({r_SM_Main_adj_5161}), .\r_Bit_Index[0] (r_Bit_Index_adj_5163[0]), 
         .n42123(n42123), .n27820(n27820), .tx_o(tx_o), .n19247(n19247), 
         .n49552(n49552), .n28192(n28192), .n4_adj_6(n4_adj_5007), .n28212(n28212), 
         .VCC_net(VCC_net), .tx_enable(tx_enable), .n4_adj_7(n4_adj_5013), 
         .r_SM_Main_adj_14({r_SM_Main}), .r_Rx_Data(r_Rx_Data), .\r_SM_Main_2__N_3442[2] (r_SM_Main_2__N_3442[2]), 
         .n27824(n27824), .\r_Bit_Index[0]_adj_11 (r_Bit_Index[0]), .n26628(n26628), 
         .n33696(n33696), .RX_N_10(RX_N_10), .n42126(n42126), .n41813(n41813), 
         .n28224(n28224), .n28182(n28182), .n28181(n28181), .n28180(n28180), 
         .n27784(n27784), .n28179(n28179), .n28178(n28178), .n28177(n28177), 
         .n28176(n28176), .n42185(n42185), .n28215(n28215), .n26633(n26633), 
         .n4_adj_12(n4_adj_5009), .n4_adj_13(n4_adj_4984)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(140[8] 163[4])
    SB_LUT4 i1_4_lut_adj_1830 (.I0(n2118), .I1(n2119), .I2(n45250), .I3(n2120), 
            .O(n45256));
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'hfffe;
    EEPROM eeprom (.CLK_c(CLK_c), .\state[3] (state_adj_5170[3]), .n6(n6_adj_5032), 
           .GND_net(GND_net), .read(read), .\state[0] (state_adj_5154[0]), 
           .enable_slow_N_4090(enable_slow_N_4090), .n4226({n4227}), .\state[1] (state_adj_5154[1]), 
           .\state[2] (state_adj_5170[2]), .n7(n7_adj_5098), .n28191(n28191), 
           .rw(rw), .n41955(n41955), .data_ready(data_ready), .n41845(n41845), 
           .n41841(n41841), .n43002(n43002), .n43073(n43073), .n34306(n34306), 
           .\state_7__N_3987[0] (state_7__N_3987[0]), .\state_7__N_4003[3] (state_7__N_4003[3]), 
           .\saved_addr[0] (saved_addr[0]), .\state[0]_adj_2 (state_adj_5170[0]), 
           .n5538(n5538), .n33499(n33499), .sda_enable(sda_enable), .scl_enable(scl_enable), 
           .n10(n10_adj_5097), .n6014(n6014), .n8(n8_adj_5089), .VCC_net(VCC_net), 
           .n28202(n28202), .data({data}), .sda_out(sda_out), .n28194(n28194), 
           .n47597(n47597), .scl(scl), .n26652(n26652), .n28174(n28174), 
           .n28170(n28170), .n28169(n28169), .n28168(n28168), .n28167(n28167), 
           .n28166(n28166), .n28165(n28165), .n33700(n33700), .n4(n4_adj_4981), 
           .n4_adj_3(n4_adj_4980), .n26657(n26657)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(289[10] 300[6])
    pwm PWM (.n48297(n48297), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n26499(n26499), .pwm_counter({pwm_counter}), .GND_net(GND_net), 
        .n26497(n26497)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (\neo_pixel_transmitter.done , 
            CLK_c, n34515, \state[1] , \state[0] , GND_net, n2380, 
            n30301, \neo_pixel_transmitter.t0 , n28262, neopxl_color, 
            n28261, n28260, n28259, n28258, n28257, n28256, n28255, 
            n28254, n47523, n28253, n28252, n28251, n28250, n28249, 
            n28248, timer, VCC_net, n28247, n28246, n28245, n28244, 
            n28243, n28242, n28241, n28240, n28239, n28238, n28237, 
            n28236, n28235, n28234, n28233, n28232, n12, NEOPXL_c, 
            n28163, LED_c) /* synthesis syn_module_defined=1 */ ;
    output \neo_pixel_transmitter.done ;
    input CLK_c;
    output n34515;
    output \state[1] ;
    output \state[0] ;
    input GND_net;
    output n2380;
    output n30301;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input n28262;
    input [23:0]neopxl_color;
    input n28261;
    input n28260;
    input n28259;
    input n28258;
    input n28257;
    input n28256;
    input n28255;
    input n28254;
    output n47523;
    input n28253;
    input n28252;
    input n28251;
    input n28250;
    input n28249;
    input n28248;
    output [31:0]timer;
    input VCC_net;
    input n28247;
    input n28246;
    input n28245;
    input n28244;
    input n28243;
    input n28242;
    input n28241;
    input n28240;
    input n28239;
    input n28238;
    input n28237;
    input n28236;
    input n28235;
    input n28234;
    input n28233;
    input n28232;
    input n12;
    output NEOPXL_c;
    input n28163;
    input LED_c;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire \neo_pixel_transmitter.done_N_636 , n42167, n30298, start, 
        n43053, n45, n43000, n48266, n42927, n4, n48267, \neo_pixel_transmitter.done_N_642 ;
    wire [31:0]n255;
    
    wire n27723;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n28057, n4_adj_4823, n113, n167, n147, n47535, n47534, 
        n156, n41189, n3017, n49247, n2903;
    wire [31:0]n2951;
    
    wire n2918, n3002, n2889, n2988, n2892, n2991, n2887, n2986, 
        n30674, n2899, n2998, n2908, n3007, n2900, n2999, n2886, 
        n2985, n2909, n3008, n2890, n2989, n2901, n3000, n2888, 
        n2987, n2904, n3003, n2896, n2995, n2894, n2993, n2905, 
        n3004, n2891, n2990, n2893, n2992, n2907, n3006, n2895, 
        n2994, n2898, n2997, n2902, n3001, n2906, n3005, n2897, 
        n2996, n2984, n44, n42, n43, n41, n40, n39, n50, n45_adj_4824, 
        n32, n42_adj_4825, n2885, n38, n43_adj_4826, n40_adj_4827, 
        n46, n39_adj_4828, n47, n2819, n49246;
    wire [31:0]n3149;
    
    wire n3116, n3209, n3104, n3103, n3106, n3098, n46_adj_4829, 
        n3096, n3109, n35, n3085, n3087, n3086, n3088, n42_adj_4830, 
        n3091, n3092, n32_adj_4831, n3093, n3095, n3094, n3101, 
        n44_adj_4832, n3108, n3102, n50_adj_4833, n3100, n3084, 
        n3083, n48, n3089, n3090, n49, n3107, n3105, n3099, 
        n3097, n47_adj_4834, n39_adj_4835, n35_adj_4836, n33, n45686, 
        n41_adj_4837, n45688, n45690, n11, n23, n45684, n45692, 
        n45700, n43_adj_4838, n45704, n45706, n45708, n13, n46104, 
        n19, n46106, n46108, n46112, n46114, n45710, n44606, n55, 
        n57, n45716, n59, n61, n46490, n39350, n30278, n60, 
        n20, n46404, n28098, n27897, n49883, n49350, n49344, n46770;
    wire [4:0]color_bit_N_622;
    
    wire n49296, n49524, n47580, n49254, n48438;
    wire [3:0]state_3__N_428;
    
    wire n2696;
    wire [31:0]n2753;
    
    wire n2720, n2795, n2691, n2790, n2707, n2806, n2700, n2799, 
        n2709, n2808, n2703, n2802, n2708, n2807, n2688, n2787, 
        n2701, n2800, n2694, n2793, n2695, n2794, n2690, n2789, 
        n2692, n2791, n2702, n2801, n2699, n2798, n2693, n2792, 
        n2705, n2804, n2706, n2805, n2697, n2796, n2704, n2803, 
        n2689, n2788, n2809, n2698, n2797, n30, n40_adj_4839, 
        n26, n37245, n38_adj_4840, n2786, n44_adj_4841, n42_adj_4842, 
        n43_adj_4843, n41_adj_4844, n2589;
    wire [31:0]n2654;
    
    wire n2621, n2604, n2603, n2600, n2606, n2608, n2607, n2602, 
        n2609, n2605, n37244, n2601, n2599, n2593, n2591, n2592, 
        n2590, n2597, n2595, n2596, n2594, n37243, n2598, n29, 
        n37, n36, n42_adj_4845, n40_adj_4846, n2687, n41_adj_4847, 
        n39_adj_4848, n37242, n37241;
    wire [31:0]n1;
    
    wire n37240, n37239, n37238, n2508;
    wire [31:0]n2555;
    
    wire n2522, n2502, n2506, n2497, n2501, n2509, n2504, n2498, 
        n2500, n2505, n2503, n2499, n2492, n2491, n2490, n2496, 
        n2494, n2495, n2493, n2507, n28_adj_4854, n35_adj_4855, 
        n2588, n34, n40_adj_4856, n38_adj_4857, n39_adj_4858, n37_adj_4859, 
        n37237, n37236, n37235, n46743, n46744, n46747, n46746, 
        n40382, n2405;
    wire [31:0]n2456;
    
    wire n2423, n2403, n37234, n2406, n2409, n2407, n2395, n2393, 
        n2394, n2392, n2399, n2397, n2398, n2396, n2400, n2401, 
        n2402, n2404, n2408, n2391, n2489, n22, n36_adj_4861, 
        n27_adj_4862, n34_adj_4863, n33_adj_4864, n37_adj_4865, n39_adj_4866, 
        n37233, n160, n37380, n46398, n37379, n46396, n37378, 
        n46394, n37377, n46392, n1499, n1400, n37835, n1433;
    wire [31:0]n1466;
    
    wire n1401, n37834, n1402, n37833, n1403, n37832, n1404, n37831, 
        n37232, n1405, n37830, n1406, n37829, n1407, n37828, n1408, 
        n37827, n1409, n37826, n37376, n46390, n2307;
    wire [31:0]n2357;
    
    wire n2324, n2301, n2299, n2303, n2300, n37231, n2302, n2294, 
        n2293, n2292, n2297, n2296, n37375, n46388, n2298, n2295, 
        n37374, n46386, n2305, n2304, n37373, n46384, n37230, 
        n2308, n2306, n37372, n46382, n2309, n34_adj_4869, n25_adj_4870, 
        n32_adj_4871, n2390, n31_adj_4872, n35_adj_4873, n37_adj_4874, 
        n1301, n38307, n1334;
    wire [31:0]n1367;
    
    wire n1302, n38306, n37371, n46380, n46_adj_4876, n44_adj_4877, 
        n45_adj_4878, n43_adj_4879, n42_adj_4880, n1303, n38305, n41_adj_4881, 
        n52, n47_adj_4882, n11_adj_4883, n37370, n46378, n1304, 
        n38304, n47529, n47530, n12_adj_4884, n1235, n49249, n14, 
        n1204, n1209, n12_adj_4885, n1205, n1208, n1207, n1206, 
        n13_adj_4886, n1203, n1202, n2196;
    wire [31:0]n2258;
    
    wire n2225, n2200, n2194, n2195, n2197, n2198, n2201, n2202, 
        n2208, n2207, n2209, n2204, n2205, n2199, n2206, n1305, 
        n38303, n2193, n2203, n30_adj_4887, n34405, n2291, n34_adj_4888, 
        n32_adj_4889, n33_adj_4890, n31_adj_4891, n37369, n46376;
    wire [31:0]one_wire_N_579;
    
    wire n4_adj_4893, n46352, n46354, n29_adj_4894, n37229, n1306, 
        n38302, n37368, n46374, n1103, n48865, n1037, n39004, 
        n37367, n46372, n1104, n48792, n39003, n1307, n38301, 
        n1105, n1006, n39002, n48737, n1308, n38300, n1106, n1007, 
        n39001, n48738, n1107, n1008, n39000, n1108, n1009, n49244, 
        n38999, n1309, n38299, n37228, n1109, n1136, n38998, n38997, 
        n38996, n38995, n38994, n38993, n49245, n38992, n1697, 
        n1598, n38991, n1631;
    wire [31:0]n1664;
    
    wire n1599, n38990, n1600, n38989, n1601, n38988, n1602, n38987, 
        n1603, n38986, n1604, n38985, n1605, n38984, n37366, n46370, 
        n1606, n38983, n1607, n38982, n1608, n38981, n1609, n38980, 
        n1796, n38979, n1730;
    wire [31:0]n1763;
    
    wire n1698, n38978, n1699, n38977, n1700, n38976, n1701, n38975, 
        n1702, n38974, n1703, n38973, n1704, n38972, n1705, n38971, 
        n1706, n38970, n1707, n38969, n37365, n46368, n1708, n38968, 
        n1709, n38967, n1895, n38966, n1829;
    wire [31:0]n1862;
    
    wire n1797, n38965, n1798, n38964, n1799, n38963, n1800, n38962, 
        n1801, n38961, n1802, n38960, n1803, n38959, n1804, n38958, 
        n1805, n38957, n1806, n38956, n1807, n38955, n1808, n38954, 
        n1809, n38953, n1994, n38952, n1928;
    wire [31:0]n1961;
    
    wire n1896, n38951, n1897, n38950, n1898, n38949, n1899, n38948, 
        n1900, n38947, n1901, n38946, n1902, n38945, n1903, n38944, 
        n1904, n38943, n1905, n38942, n1906, n38941, n1907, n38940, 
        n1908, n38939, n1909, n38938, n2093, n38937, n2027;
    wire [31:0]n2060;
    
    wire n1995, n38936, n1996, n38935, n1997, n38934, n1998, n38933, 
        n1999, n38932, n2000, n38931, n2001, n38930, n2002, n38929, 
        n2003, n38928, n2004, n38927, n2005, n38926, n2006, n38925, 
        n2007, n38924, n2008, n38923, n2009, n38922, n2192, n38921, 
        n2126;
    wire [31:0]n2159;
    
    wire n2094, n38920, n37364, n46366, n2095, n38919, n2096, 
        n38918, n2097, n38917, n2098, n38916, n2099, n38915, n2100, 
        n38914, n2101, n38913, n2102, n38912, n2103, n38911, n2104, 
        n38910, n2105, n38909, n2106, n38908, n2107, n38907, n2108, 
        n38906, n2109, n38905, n38904, n38903, n38902, n38901, 
        n38900, n38899, n38898, n37363, n46364, n38897, n37362, 
        n46362;
    wire [31:0]n133;
    
    wire n38896, n49521, n38895, n38894, n38893, n38892, n38891, 
        n38890, n38889, n38888, n38887, n38886, n38885, n38884, 
        n37227, n38883, n38882, n38881, n38880, n38879, n38878, 
        n38877, n38876, n38875, n38874, n38873, n38872, n38871, 
        n38870, n38869, n38868, n38867, n38866, n38865, n38864, 
        n38863, n38862, n38861, n38860, n38859, n38858, n38857, 
        n38856, n38855, n38854, n37361, n38853, n37360, n38852, 
        n38851, n38850, n38849, n38848, n38847, n38846, n38845, 
        n38844, n38843, n38842, n38841, n38840, n38839, n38838, 
        n38837, n38836, n38835, n38834, n38833, n38832, n38831, 
        n38830, n38829, n37359, n38828, n38827, n38826, n38825, 
        n38824, n37358, n38823, n37226, n38822, n38821, n49347, 
        n49341, n38820, n38819, n38818, n37357, n38817, n38816, 
        n37225, n37356, n46350, n37355, n46348, n37354, n38815, 
        n38814, n37353, n37352, n37351, n37224, n38813, n38812, 
        n37223, n38811, n38810, n38809, n38808, n37350, n38807, 
        n38806, n37222, n38805, n38804, n38803, n38802, n38801, 
        n38800, n37609, n1532;
    wire [31:0]n1565;
    
    wire n1500, n37608, n1501, n37607, n38799, n38798, n1502, 
        n37606, n38797, n1503, n37605, n38796, n1504, n37604, 
        n38795, n37221, n38794, n38793, n38792, n38791, n1505, 
        n37603, n1506, n37602, n1507, n37601, n38790, n1508, n37600, 
        n38789, n1509, n37599, n38788, n37220, n38787, n38786, 
        n38785, n38784, n38783, n38782, n28_adj_4899, n31_adj_4900, 
        n22_adj_4901, n38781, n30_adj_4902, n34_adj_4903, n21_adj_4904, 
        n38780, n38779, n38778, n38777, n38776, n38775, n38774, 
        n38773, n38772, n38771, n38770, n38769, n38768, n38767, 
        n38766, n38765, n38764, n38763, n38762, n38761, n37219, 
        n38760, n38759, n38758, n37218, n38757, n38756, n38755, 
        n38754, n38753, n38752, n38751, n38750, n38749, n38748, 
        n38747, n38746, n38745, n37217, n38744, n38743, n38742, 
        n38741, n38740, n38739, n38738, n38737, n38736, n38735, 
        n38734, n38733, n38732, n38731, n38730, n38729, n38728, 
        n38727, n38726, n38725, n38724, n38723, n38722, n38721, 
        n38720, n38719, n38718, n38717, n38716, n38715, n38714, 
        n37216, n38713, n38712, n38711, n38710, n38709, n38708, 
        n38707, n38706, n38705, n38704, n38703, n38702, n38701, 
        n38700, n38699, n38698, n38697, n38696, n38695, n38694, 
        n38693, n38692, n37215, n38691, n38690, n38689, n38688, 
        n38687, n38686, n38685, n38684, n38683, n38682, n38681, 
        n38680;
    wire [31:0]n971;
    
    wire n37334, n37333, n27993, n37332, n27950, n37331, n25171, 
        n37330, n25173, n27956, n44951, n56, n2_adj_4905, n8_adj_4906, 
        n49293, n18_adj_4907, n34401, n30_adj_4908, n28_adj_4909, 
        n29_adj_4910, n27_adj_4911, n34399, n28_adj_4915, n26_adj_4916, 
        n27_adj_4917, n25_adj_4918, n20_adj_4919, n26_adj_4920, n16_adj_4921, 
        n24_adj_4922, n28_adj_4923, n38535, n38534, n38533, n38532, 
        n38531, n38530, n38529, n38528, n38527, n38526, n38525, 
        n38524, n38523, n38522, n38521, n38520, n38519, n38518, 
        n38517, n38516, n38515, n38514, n38513, n38512, n38511, 
        n38510, n38509, n38508, n38507, n38506, n38505, n38504, 
        n38503, n38502, n38501, n38500, n38499, n38498, n38497, 
        n24_adj_4924, n17_adj_4925, n22_adj_4926, n26_adj_4927, n18_adj_4928, 
        n21_adj_4929, n20_adj_4930, n24_adj_4931, n18_adj_4932, n20_adj_4933, 
        n15_adj_4934, n14_adj_4935, n20_adj_4936, n18_adj_4937, n22_adj_4938, 
        n34387, n12_adj_4939, n7_adj_4940, n14_adj_4941, n12_adj_4942, 
        n16_adj_4943, n12_adj_4944, n16_adj_4945, n17_adj_4946, n49251;
    
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n42167), .D(\neo_pixel_transmitter.done_N_636 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i48_4_lut (.I0(n30298), .I1(n34515), .I2(\state[1] ), .I3(start), 
            .O(n43053));
    defparam i48_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i33313_4_lut (.I0(n43053), .I1(n45), .I2(\neo_pixel_transmitter.done ), 
            .I3(n43000), .O(n48266));
    defparam i33313_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i33314_4_lut (.I0(n48266), .I1(n42927), .I2(\state[0] ), .I3(n4), 
            .O(n48267));
    defparam i33314_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 i117_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_642 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i117_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n27723), .D(n255[1]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n27723), .D(n255[2]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n27723), .D(n255[3]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n27723), .D(n255[4]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n27723), .D(n255[5]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n27723), .D(n255[6]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n27723), .D(n255[7]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n27723), .D(n255[8]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n27723), .D(n255[9]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n27723), 
            .D(n255[10]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n27723), 
            .D(n255[11]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n27723), 
            .D(n255[12]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n27723), 
            .D(n255[13]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n27723), 
            .D(n255[14]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n27723), 
            .D(n255[15]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n27723), 
            .D(n255[16]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n27723), 
            .D(n255[17]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n27723), 
            .D(n255[18]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n27723), 
            .D(n255[19]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n27723), 
            .D(n255[20]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n27723), 
            .D(n255[21]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n27723), 
            .D(n255[22]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n27723), 
            .D(n255[23]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n27723), 
            .D(n255[24]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n27723), 
            .D(n255[25]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n27723), 
            .D(n255[26]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i17240_4_lut (.I0(n4_adj_4823), .I1(n113), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n167));   // verilog/neopixel.v(16[20:25])
    defparam i17240_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n147), .I2(n167), .I3(start), 
            .O(n2380));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_4_lut.LUT_INIT = 16'h5554;
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n27723), 
            .D(n255[27]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n27723), 
            .D(n255[28]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n27723), 
            .D(n255[29]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n27723), 
            .D(n255[30]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n27723), 
            .D(n255[31]), .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i32726_4_lut (.I0(n113), .I1(n147), .I2(n4_adj_4823), .I3(\state[0] ), 
            .O(n47535));   // verilog/neopixel.v(16[20:25])
    defparam i32726_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i18_4_lut (.I0(n47535), .I1(n47534), .I2(\state[1] ), .I3(n156), 
            .O(n41189));   // verilog/neopixel.v(16[20:25])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i34294_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49247));
    defparam i34294_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i2029_3_lut (.I0(n2903), .I1(n2951[13]), .I2(n2918), 
            .I3(GND_net), .O(n3002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2015_3_lut (.I0(n2889), .I1(n2951[27]), .I2(n2918), 
            .I3(GND_net), .O(n2988));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2018_3_lut (.I0(n2892), .I1(n2951[24]), .I2(n2918), 
            .I3(GND_net), .O(n2991));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2013_3_lut (.I0(n2887), .I1(n2951[29]), .I2(n2918), 
            .I3(GND_net), .O(n2986));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17624_3_lut (.I0(bit_ctr[6]), .I1(n2951[6]), .I2(n2918), 
            .I3(GND_net), .O(n30674));
    defparam i17624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2025_3_lut (.I0(n2899), .I1(n2951[17]), .I2(n2918), 
            .I3(GND_net), .O(n2998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2034_3_lut (.I0(n2908), .I1(n2951[8]), .I2(n2918), 
            .I3(GND_net), .O(n3007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2026_3_lut (.I0(n2900), .I1(n2951[16]), .I2(n2918), 
            .I3(GND_net), .O(n2999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2012_3_lut (.I0(n2886), .I1(n2951[30]), .I2(n2918), 
            .I3(GND_net), .O(n2985));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2035_3_lut (.I0(n2909), .I1(n2951[7]), .I2(n2918), 
            .I3(GND_net), .O(n3008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2016_3_lut (.I0(n2890), .I1(n2951[26]), .I2(n2918), 
            .I3(GND_net), .O(n2989));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2027_3_lut (.I0(n2901), .I1(n2951[15]), .I2(n2918), 
            .I3(GND_net), .O(n3000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2014_3_lut (.I0(n2888), .I1(n2951[28]), .I2(n2918), 
            .I3(GND_net), .O(n2987));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2030_3_lut (.I0(n2904), .I1(n2951[12]), .I2(n2918), 
            .I3(GND_net), .O(n3003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2022_3_lut (.I0(n2896), .I1(n2951[20]), .I2(n2918), 
            .I3(GND_net), .O(n2995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2020_3_lut (.I0(n2894), .I1(n2951[22]), .I2(n2918), 
            .I3(GND_net), .O(n2993));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2031_3_lut (.I0(n2905), .I1(n2951[11]), .I2(n2918), 
            .I3(GND_net), .O(n3004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2017_3_lut (.I0(n2891), .I1(n2951[25]), .I2(n2918), 
            .I3(GND_net), .O(n2990));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2019_3_lut (.I0(n2893), .I1(n2951[23]), .I2(n2918), 
            .I3(GND_net), .O(n2992));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2033_3_lut (.I0(n2907), .I1(n2951[9]), .I2(n2918), 
            .I3(GND_net), .O(n3006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2021_3_lut (.I0(n2895), .I1(n2951[21]), .I2(n2918), 
            .I3(GND_net), .O(n2994));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2024_3_lut (.I0(n2898), .I1(n2951[18]), .I2(n2918), 
            .I3(GND_net), .O(n2997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2028_3_lut (.I0(n2902), .I1(n2951[14]), .I2(n2918), 
            .I3(GND_net), .O(n3001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2032_3_lut (.I0(n2906), .I1(n2951[10]), .I2(n2918), 
            .I3(GND_net), .O(n3005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2023_3_lut (.I0(n2897), .I1(n2951[19]), .I2(n2918), 
            .I3(GND_net), .O(n2996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1530 (.I0(n2984), .I1(n2996), .I2(n3005), .I3(n3001), 
            .O(n44));
    defparam i18_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2997), .I1(n2994), .I2(n3006), .I3(n2992), 
            .O(n42));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n2990), .I1(n3004), .I2(n2993), .I3(n2995), 
            .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n3003), .I1(n2987), .I2(n3000), .I3(n2989), 
            .O(n41));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n3008), .I1(n2985), .I2(n2999), .I3(n3007), 
            .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2998), .I1(bit_ctr[5]), .I2(n30674), .I3(GND_net), 
            .O(n39));
    defparam i13_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n2986), .I1(n2991), .I2(n2988), .I3(n3002), 
            .O(n45_adj_4824));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45_adj_4824), .I1(n50), .I2(n39), .I3(n40), 
            .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n2897), .I1(bit_ctr[6]), .I2(n2909), .I3(GND_net), 
            .O(n32));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i17_4_lut_adj_1531 (.I0(n2907), .I1(n2908), .I2(n2903), .I3(n2904), 
            .O(n42_adj_4825));
    defparam i17_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut_adj_1532 (.I0(n2899), .I1(n2886), .I2(n2885), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut_adj_1532.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1533 (.I0(n2902), .I1(n2898), .I2(n2906), .I3(n2905), 
            .O(n43_adj_4826));
    defparam i18_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1534 (.I0(n2891), .I1(n2893), .I2(n2892), .I3(n2894), 
            .O(n40_adj_4827));
    defparam i15_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n2895), .I1(n42_adj_4825), .I2(n32), .I3(n2896), 
            .O(n46));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1535 (.I0(n2887), .I1(n2889), .I2(n2888), .I3(n2890), 
            .O(n39_adj_4828));
    defparam i14_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43_adj_4826), .I1(n2901), .I2(n38), .I3(n2900), 
            .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1536 (.I0(n47), .I1(n39_adj_4828), .I2(n46), 
            .I3(n40_adj_4827), .O(n2918));
    defparam i24_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i34293_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49246));
    defparam i34293_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i2172_3_lut (.I0(bit_ctr[4]), .I1(n3149[4]), .I2(n3116), 
            .I3(GND_net), .O(n3209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_4_lut_adj_1537 (.I0(n3104), .I1(n3103), .I2(n3106), .I3(n3098), 
            .O(n46_adj_4829));
    defparam i19_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[4]), .I1(n3096), .I2(n3109), .I3(GND_net), 
            .O(n35));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1538 (.I0(n3085), .I1(n3087), .I2(n3086), .I3(n3088), 
            .O(n42_adj_4830));
    defparam i15_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n3091), .I1(n3092), .I2(GND_net), .I3(GND_net), 
            .O(n32_adj_4831));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1539 (.I0(n3093), .I1(n3095), .I2(n3094), .I3(n3101), 
            .O(n44_adj_4832));
    defparam i17_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n35), .I1(n46_adj_4829), .I2(n3108), .I3(n3102), 
            .O(n50_adj_4833));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1540 (.I0(n3100), .I1(n42_adj_4830), .I2(n3084), 
            .I3(n3083), .O(n48));
    defparam i21_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1541 (.I0(n3089), .I1(n44_adj_4832), .I2(n32_adj_4831), 
            .I3(n3090), .O(n49));
    defparam i22_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n3107), .I1(n3105), .I2(n3099), .I3(n3097), 
            .O(n47_adj_4834));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n47_adj_4834), .I1(n49), .I2(n48), .I3(n50_adj_4833), 
            .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2157_3_lut (.I0(n3095), .I1(n3149[19]), .I2(n3116), 
            .I3(GND_net), .O(n39_adj_4835));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2159_3_lut (.I0(n3097), .I1(n3149[17]), .I2(n3116), 
            .I3(GND_net), .O(n35_adj_4836));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2160_3_lut (.I0(n3098), .I1(n3149[16]), .I2(n3116), 
            .I3(GND_net), .O(n33));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1542 (.I0(n3100), .I1(n39_adj_4835), .I2(n3149[14]), 
            .I3(n3116), .O(n45686));
    defparam i1_4_lut_adj_1542.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2156_3_lut (.I0(n3094), .I1(n3149[20]), .I2(n3116), 
            .I3(GND_net), .O(n41_adj_4837));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1543 (.I0(n3101), .I1(n35_adj_4836), .I2(n3149[13]), 
            .I3(n3116), .O(n45688));
    defparam i1_4_lut_adj_1543.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1544 (.I0(n3102), .I1(n33), .I2(n3149[12]), .I3(n3116), 
            .O(n45690));
    defparam i1_4_lut_adj_1544.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2171_3_lut (.I0(n3109), .I1(n3149[5]), .I2(n3116), 
            .I3(GND_net), .O(n11));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2165_3_lut (.I0(n3103), .I1(n3149[11]), .I2(n3116), 
            .I3(GND_net), .O(n23));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1545 (.I0(n3099), .I1(n23), .I2(n3149[15]), .I3(n3116), 
            .O(n45684));
    defparam i1_4_lut_adj_1545.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1546 (.I0(n3107), .I1(n11), .I2(n3149[7]), .I3(n3116), 
            .O(n45692));
    defparam i1_4_lut_adj_1546.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1547 (.I0(n45690), .I1(n45688), .I2(n41_adj_4837), 
            .I3(n45686), .O(n45700));
    defparam i1_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2155_3_lut (.I0(n3093), .I1(n3149[21]), .I2(n3116), 
            .I3(GND_net), .O(n43_adj_4838));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1548 (.I0(n43_adj_4838), .I1(n45700), .I2(n45692), 
            .I3(n45684), .O(n45704));
    defparam i1_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1549 (.I0(n3091), .I1(n45704), .I2(n3149[23]), 
            .I3(n3116), .O(n45706));
    defparam i1_4_lut_adj_1549.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1550 (.I0(n3090), .I1(n45706), .I2(n3149[24]), 
            .I3(n3116), .O(n45708));
    defparam i1_4_lut_adj_1550.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2170_3_lut (.I0(n3108), .I1(n3149[6]), .I2(n3116), 
            .I3(GND_net), .O(n13));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1551 (.I0(n3104), .I1(n13), .I2(n3149[10]), .I3(n3116), 
            .O(n46104));
    defparam i1_4_lut_adj_1551.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2167_3_lut (.I0(n3105), .I1(n3149[9]), .I2(n3116), 
            .I3(GND_net), .O(n19));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1552 (.I0(n3106), .I1(n19), .I2(n3149[8]), .I3(n3116), 
            .O(n46106));
    defparam i1_4_lut_adj_1552.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1553 (.I0(n46104), .I1(n3096), .I2(n3149[18]), 
            .I3(n3116), .O(n46108));
    defparam i1_4_lut_adj_1553.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1554 (.I0(n46108), .I1(bit_ctr[3]), .I2(n46106), 
            .I3(n3209), .O(n46112));
    defparam i1_4_lut_adj_1554.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1555 (.I0(n3092), .I1(n46112), .I2(n3149[22]), 
            .I3(n3116), .O(n46114));
    defparam i1_4_lut_adj_1555.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1556 (.I0(n3089), .I1(n45708), .I2(n3149[25]), 
            .I3(n3116), .O(n45710));
    defparam i1_4_lut_adj_1556.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1557 (.I0(n46114), .I1(n3088), .I2(n3149[26]), 
            .I3(n3116), .O(n44606));
    defparam i1_4_lut_adj_1557.LUT_INIT = 16'hfaee;
    SB_LUT4 mod_5_i2149_3_lut (.I0(n3087), .I1(n3149[27]), .I2(n3116), 
            .I3(GND_net), .O(n55));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2148_3_lut (.I0(n3086), .I1(n3149[28]), .I2(n3116), 
            .I3(GND_net), .O(n57));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1558 (.I0(n57), .I1(n55), .I2(n44606), .I3(n45710), 
            .O(n45716));
    defparam i1_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2147_3_lut (.I0(n3085), .I1(n3149[29]), .I2(n3116), 
            .I3(GND_net), .O(n59));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2146_3_lut (.I0(n3084), .I1(n3149[30]), .I2(n3116), 
            .I3(GND_net), .O(n61));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1559 (.I0(n61), .I1(n46490), .I2(n59), .I3(n45716), 
            .O(n39350));
    defparam i1_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_3_lut (.I0(n30278), .I1(n60), .I2(\state[1] ), .I3(GND_net), 
            .O(n20));   // verilog/neopixel.v(35[12] 117[6])
    defparam i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_4_lut_adj_1560 (.I0(n20), .I1(n46404), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n28098));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_4_lut_adj_1560.LUT_INIT = 16'h05c5;
    SB_LUT4 i1_4_lut_adj_1561 (.I0(\state[1] ), .I1(n30301), .I2(n60), 
            .I3(\state[0] ), .O(n27897));
    defparam i1_4_lut_adj_1561.LUT_INIT = 16'hee4e;
    SB_LUT4 i1_rep_341_2_lut (.I0(bit_ctr[3]), .I1(n39350), .I2(GND_net), 
            .I3(GND_net), .O(n49883));
    defparam i1_rep_341_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31817_3_lut (.I0(n49350), .I1(n49344), .I2(bit_ctr[2]), .I3(GND_net), 
            .O(n46770));
    defparam i31817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32949_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n39350), .I3(GND_net), 
            .O(color_bit_N_622[4]));
    defparam i32949_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i33026_4_lut (.I0(n49296), .I1(n49883), .I2(n49524), .I3(bit_ctr[2]), 
            .O(n47580));
    defparam i33026_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i33485_4_lut (.I0(n49254), .I1(n46770), .I2(bit_ctr[3]), .I3(n39350), 
            .O(n48438));   // verilog/neopixel.v(22[26:36])
    defparam i33485_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i20507_4_lut (.I0(n48438), .I1(state_3__N_428[1]), .I2(n47580), 
            .I3(color_bit_N_622[4]), .O(state_3__N_428[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i20507_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mod_5_i1886_3_lut (.I0(n2696), .I1(n2753[22]), .I2(n2720), 
            .I3(GND_net), .O(n2795));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1881_3_lut (.I0(n2691), .I1(n2753[27]), .I2(n2720), 
            .I3(GND_net), .O(n2790));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1897_3_lut (.I0(n2707), .I1(n2753[11]), .I2(n2720), 
            .I3(GND_net), .O(n2806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1890_3_lut (.I0(n2700), .I1(n2753[18]), .I2(n2720), 
            .I3(GND_net), .O(n2799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1899_3_lut (.I0(n2709), .I1(n2753[9]), .I2(n2720), 
            .I3(GND_net), .O(n2808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1893_3_lut (.I0(n2703), .I1(n2753[15]), .I2(n2720), 
            .I3(GND_net), .O(n2802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1898_3_lut (.I0(n2708), .I1(n2753[10]), .I2(n2720), 
            .I3(GND_net), .O(n2807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1878_3_lut (.I0(n2688), .I1(n2753[30]), .I2(n2720), 
            .I3(GND_net), .O(n2787));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1891_3_lut (.I0(n2701), .I1(n2753[17]), .I2(n2720), 
            .I3(GND_net), .O(n2800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1884_3_lut (.I0(n2694), .I1(n2753[24]), .I2(n2720), 
            .I3(GND_net), .O(n2793));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1885_3_lut (.I0(n2695), .I1(n2753[23]), .I2(n2720), 
            .I3(GND_net), .O(n2794));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1880_3_lut (.I0(n2690), .I1(n2753[28]), .I2(n2720), 
            .I3(GND_net), .O(n2789));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1882_3_lut (.I0(n2692), .I1(n2753[26]), .I2(n2720), 
            .I3(GND_net), .O(n2791));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1892_3_lut (.I0(n2702), .I1(n2753[16]), .I2(n2720), 
            .I3(GND_net), .O(n2801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1889_3_lut (.I0(n2699), .I1(n2753[19]), .I2(n2720), 
            .I3(GND_net), .O(n2798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1883_3_lut (.I0(n2693), .I1(n2753[25]), .I2(n2720), 
            .I3(GND_net), .O(n2792));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1895_3_lut (.I0(n2705), .I1(n2753[13]), .I2(n2720), 
            .I3(GND_net), .O(n2804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1896_3_lut (.I0(n2706), .I1(n2753[12]), .I2(n2720), 
            .I3(GND_net), .O(n2805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1887_3_lut (.I0(n2697), .I1(n2753[21]), .I2(n2720), 
            .I3(GND_net), .O(n2796));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1894_3_lut (.I0(n2704), .I1(n2753[14]), .I2(n2720), 
            .I3(GND_net), .O(n2803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1879_3_lut (.I0(n2689), .I1(n2753[29]), .I2(n2720), 
            .I3(GND_net), .O(n2788));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1900_3_lut (.I0(bit_ctr[8]), .I1(n2753[8]), .I2(n2720), 
            .I3(GND_net), .O(n2809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1888_3_lut (.I0(n2698), .I1(n2753[20]), .I2(n2720), 
            .I3(GND_net), .O(n2797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(bit_ctr[7]), .I1(n2797), .I2(n2809), .I3(GND_net), 
            .O(n30));
    defparam i6_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1562 (.I0(n2796), .I1(n2805), .I2(n2804), .I3(n2792), 
            .O(n40_adj_4839));
    defparam i16_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(n2788), .I1(n2803), .I2(GND_net), .I3(GND_net), 
            .O(n26));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n37245), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_1563 (.I0(n2801), .I1(n2791), .I2(n2789), .I3(n2794), 
            .O(n38_adj_4840));
    defparam i14_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1564 (.I0(n2786), .I1(n40_adj_4839), .I2(n30), 
            .I3(n2798), .O(n44_adj_4841));
    defparam i20_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1565 (.I0(n2802), .I1(n2808), .I2(n2799), .I3(n2806), 
            .O(n42_adj_4842));
    defparam i18_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1566 (.I0(n2790), .I1(n38_adj_4840), .I2(n26), 
            .I3(n2795), .O(n43_adj_4843));
    defparam i19_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1567 (.I0(n2793), .I1(n2800), .I2(n2787), .I3(n2807), 
            .O(n41_adj_4844));
    defparam i17_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1568 (.I0(n41_adj_4844), .I1(n43_adj_4843), .I2(n42_adj_4842), 
            .I3(n44_adj_4841), .O(n2819));
    defparam i23_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1811_3_lut (.I0(n2589), .I1(n2654[30]), .I2(n2621), 
            .I3(GND_net), .O(n2688));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1826_3_lut (.I0(n2604), .I1(n2654[15]), .I2(n2621), 
            .I3(GND_net), .O(n2703));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1825_3_lut (.I0(n2603), .I1(n2654[16]), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1822_3_lut (.I0(n2600), .I1(n2654[19]), .I2(n2621), 
            .I3(GND_net), .O(n2699));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1828_3_lut (.I0(n2606), .I1(n2654[13]), .I2(n2621), 
            .I3(GND_net), .O(n2705));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1830_3_lut (.I0(n2608), .I1(n2654[11]), .I2(n2621), 
            .I3(GND_net), .O(n2707));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1829_3_lut (.I0(n2607), .I1(n2654[12]), .I2(n2621), 
            .I3(GND_net), .O(n2706));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1824_3_lut (.I0(n2602), .I1(n2654[17]), .I2(n2621), 
            .I3(GND_net), .O(n2701));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1831_3_lut (.I0(n2609), .I1(n2654[10]), .I2(n2621), 
            .I3(GND_net), .O(n2708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1827_3_lut (.I0(n2605), .I1(n2654[14]), .I2(n2621), 
            .I3(GND_net), .O(n2704));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n37244), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1823_3_lut (.I0(n2601), .I1(n2654[18]), .I2(n2621), 
            .I3(GND_net), .O(n2700));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1821_3_lut (.I0(n2599), .I1(n2654[20]), .I2(n2621), 
            .I3(GND_net), .O(n2698));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1815_3_lut (.I0(n2593), .I1(n2654[26]), .I2(n2621), 
            .I3(GND_net), .O(n2692));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1813_3_lut (.I0(n2591), .I1(n2654[28]), .I2(n2621), 
            .I3(GND_net), .O(n2690));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1814_3_lut (.I0(n2592), .I1(n2654[27]), .I2(n2621), 
            .I3(GND_net), .O(n2691));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1812_3_lut (.I0(n2590), .I1(n2654[29]), .I2(n2621), 
            .I3(GND_net), .O(n2689));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1819_3_lut (.I0(n2597), .I1(n2654[22]), .I2(n2621), 
            .I3(GND_net), .O(n2696));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1817_3_lut (.I0(n2595), .I1(n2654[24]), .I2(n2621), 
            .I3(GND_net), .O(n2694));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1818_3_lut (.I0(n2596), .I1(n2654[23]), .I2(n2621), 
            .I3(GND_net), .O(n2695));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1816_3_lut (.I0(n2594), .I1(n2654[25]), .I2(n2621), 
            .I3(GND_net), .O(n2693));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1832_3_lut (.I0(bit_ctr[9]), .I1(n2654[9]), .I2(n2621), 
            .I3(GND_net), .O(n2709));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_32 (.CI(n37244), .I0(bit_ctr[30]), .I1(GND_net), .CO(n37245));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n37243), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1820_3_lut (.I0(n2598), .I1(n2654[21]), .I2(n2621), 
            .I3(GND_net), .O(n2697));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut_adj_1569 (.I0(n2697), .I1(bit_ctr[8]), .I2(n2709), 
            .I3(GND_net), .O(n29));
    defparam i6_3_lut_adj_1569.LUT_INIT = 16'heaea;
    SB_LUT4 i14_4_lut_adj_1570 (.I0(n2693), .I1(n2695), .I2(n2694), .I3(n2696), 
            .O(n37));
    defparam i14_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2689), .I1(n2691), .I2(n2690), .I3(n2692), 
            .O(n36));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1571 (.I0(n37), .I1(n29), .I2(n2698), .I3(n2700), 
            .O(n42_adj_4845));
    defparam i19_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1572 (.I0(n2704), .I1(n2708), .I2(n2701), .I3(n2706), 
            .O(n40_adj_4846));
    defparam i17_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1573 (.I0(n2703), .I1(n36), .I2(n2688), .I3(n2687), 
            .O(n41_adj_4847));
    defparam i18_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1574 (.I0(n2707), .I1(n2705), .I2(n2699), .I3(n2702), 
            .O(n39_adj_4848));
    defparam i16_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1575 (.I0(n39_adj_4848), .I1(n41_adj_4847), .I2(n40_adj_4846), 
            .I3(n42_adj_4845), .O(n2720));
    defparam i22_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_31 (.CI(n37243), .I0(bit_ctr[29]), .I1(GND_net), .CO(n37244));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n37242), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n37242), .I0(bit_ctr[28]), .I1(GND_net), .CO(n37243));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n37241), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_29 (.CI(n37241), .I0(bit_ctr[27]), .I1(GND_net), .CO(n37242));
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n37240), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_28 (.CI(n37240), .I0(bit_ctr[26]), .I1(GND_net), .CO(n37241));
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n37239), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_27 (.CI(n37239), .I0(bit_ctr[25]), .I1(GND_net), .CO(n37240));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n37238), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1762_3_lut (.I0(n2508), .I1(n2555[12]), .I2(n2522), 
            .I3(GND_net), .O(n2607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1756_3_lut (.I0(n2502), .I1(n2555[18]), .I2(n2522), 
            .I3(GND_net), .O(n2601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1760_3_lut (.I0(n2506), .I1(n2555[14]), .I2(n2522), 
            .I3(GND_net), .O(n2605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1751_3_lut (.I0(n2497), .I1(n2555[23]), .I2(n2522), 
            .I3(GND_net), .O(n2596));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1755_3_lut (.I0(n2501), .I1(n2555[19]), .I2(n2522), 
            .I3(GND_net), .O(n2600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1763_3_lut (.I0(n2509), .I1(n2555[11]), .I2(n2522), 
            .I3(GND_net), .O(n2608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1758_3_lut (.I0(n2504), .I1(n2555[16]), .I2(n2522), 
            .I3(GND_net), .O(n2603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1752_3_lut (.I0(n2498), .I1(n2555[22]), .I2(n2522), 
            .I3(GND_net), .O(n2597));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1754_3_lut (.I0(n2500), .I1(n2555[20]), .I2(n2522), 
            .I3(GND_net), .O(n2599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1759_3_lut (.I0(n2505), .I1(n2555[15]), .I2(n2522), 
            .I3(GND_net), .O(n2604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1757_3_lut (.I0(n2503), .I1(n2555[17]), .I2(n2522), 
            .I3(GND_net), .O(n2602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1753_3_lut (.I0(n2499), .I1(n2555[21]), .I2(n2522), 
            .I3(GND_net), .O(n2598));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1746_3_lut (.I0(n2492), .I1(n2555[28]), .I2(n2522), 
            .I3(GND_net), .O(n2591));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1745_3_lut (.I0(n2491), .I1(n2555[29]), .I2(n2522), 
            .I3(GND_net), .O(n2590));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1744_3_lut (.I0(n2490), .I1(n2555[30]), .I2(n2522), 
            .I3(GND_net), .O(n2589));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1750_3_lut (.I0(n2496), .I1(n2555[24]), .I2(n2522), 
            .I3(GND_net), .O(n2595));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1748_3_lut (.I0(n2494), .I1(n2555[26]), .I2(n2522), 
            .I3(GND_net), .O(n2593));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1749_3_lut (.I0(n2495), .I1(n2555[25]), .I2(n2522), 
            .I3(GND_net), .O(n2594));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1747_3_lut (.I0(n2493), .I1(n2555[27]), .I2(n2522), 
            .I3(GND_net), .O(n2592));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1764_3_lut (.I0(bit_ctr[10]), .I1(n2555[10]), .I2(n2522), 
            .I3(GND_net), .O(n2609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1761_3_lut (.I0(n2507), .I1(n2555[13]), .I2(n2522), 
            .I3(GND_net), .O(n2606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut_adj_1576 (.I0(bit_ctr[9]), .I1(n2606), .I2(n2609), 
            .I3(GND_net), .O(n28_adj_4854));   // verilog/neopixel.v(22[26:36])
    defparam i6_3_lut_adj_1576.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1577 (.I0(n2592), .I1(n2594), .I2(n2593), .I3(n2595), 
            .O(n35_adj_4855));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2589), .I1(n2590), .I2(n2588), .I3(n2591), 
            .O(n34));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1578 (.I0(n35_adj_4855), .I1(n2598), .I2(n28_adj_4854), 
            .I3(n2602), .O(n40_adj_4856));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1579 (.I0(n2604), .I1(n2599), .I2(n2597), .I3(n2603), 
            .O(n38_adj_4857));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2608), .I1(n34), .I2(n2600), .I3(GND_net), 
            .O(n39_adj_4858));   // verilog/neopixel.v(22[26:36])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1580 (.I0(n2596), .I1(n2605), .I2(n2601), .I3(n2607), 
            .O(n37_adj_4859));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1581 (.I0(n37_adj_4859), .I1(n39_adj_4858), .I2(n38_adj_4857), 
            .I3(n40_adj_4856), .O(n2621));   // verilog/neopixel.v(22[26:36])
    defparam i21_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_26 (.CI(n37238), .I0(bit_ctr[24]), .I1(GND_net), .CO(n37239));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n37237), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_25 (.CI(n37237), .I0(bit_ctr[23]), .I1(GND_net), .CO(n37238));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n37236), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_24 (.CI(n37236), .I0(bit_ctr[22]), .I1(GND_net), .CO(n37237));
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n28262));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n37235), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n37235), .I0(bit_ctr[21]), .I1(GND_net), .CO(n37236));
    SB_LUT4 i31790_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46743));
    defparam i31790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31791_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46744));
    defparam i31791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31794_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46747));
    defparam i31794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31793_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46746));
    defparam i31793_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n28261));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n28260));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n28259));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n28258));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n28257));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n28256));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n28255));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n28254));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i32673_3_lut_4_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(\state[0] ), 
            .I3(n40382), .O(n47523));
    defparam i32673_3_lut_4_lut.LUT_INIT = 16'h0070;
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n28253));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n28252));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n28251));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n28250));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n28249));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n28248));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1691_3_lut (.I0(n2405), .I1(n2456[16]), .I2(n2423), 
            .I3(GND_net), .O(n2504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1689_3_lut (.I0(n2403), .I1(n2456[18]), .I2(n2423), 
            .I3(GND_net), .O(n2502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n37234), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1692_3_lut (.I0(n2406), .I1(n2456[15]), .I2(n2423), 
            .I3(GND_net), .O(n2505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1695_3_lut (.I0(n2409), .I1(n2456[12]), .I2(n2423), 
            .I3(GND_net), .O(n2508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1693_3_lut (.I0(n2407), .I1(n2456[14]), .I2(n2423), 
            .I3(GND_net), .O(n2506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(n40382), 
            .I3(GND_net), .O(state_3__N_428[1]));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 mod_5_i1681_3_lut (.I0(n2395), .I1(n2456[26]), .I2(n2423), 
            .I3(GND_net), .O(n2494));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1679_3_lut (.I0(n2393), .I1(n2456[28]), .I2(n2423), 
            .I3(GND_net), .O(n2492));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1680_3_lut (.I0(n2394), .I1(n2456[27]), .I2(n2423), 
            .I3(GND_net), .O(n2493));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1678_3_lut (.I0(n2392), .I1(n2456[29]), .I2(n2423), 
            .I3(GND_net), .O(n2491));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1685_3_lut (.I0(n2399), .I1(n2456[22]), .I2(n2423), 
            .I3(GND_net), .O(n2498));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1683_3_lut (.I0(n2397), .I1(n2456[24]), .I2(n2423), 
            .I3(GND_net), .O(n2496));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1684_3_lut (.I0(n2398), .I1(n2456[23]), .I2(n2423), 
            .I3(GND_net), .O(n2497));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1682_3_lut (.I0(n2396), .I1(n2456[25]), .I2(n2423), 
            .I3(GND_net), .O(n2495));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1696_3_lut (.I0(bit_ctr[11]), .I1(n2456[11]), .I2(n2423), 
            .I3(GND_net), .O(n2509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1686_3_lut (.I0(n2400), .I1(n2456[21]), .I2(n2423), 
            .I3(GND_net), .O(n2499));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1687_3_lut (.I0(n2401), .I1(n2456[20]), .I2(n2423), 
            .I3(GND_net), .O(n2500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1688_3_lut (.I0(n2402), .I1(n2456[19]), .I2(n2423), 
            .I3(GND_net), .O(n2501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1690_3_lut (.I0(n2404), .I1(n2456[17]), .I2(n2423), 
            .I3(GND_net), .O(n2503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1694_3_lut (.I0(n2408), .I1(n2456[13]), .I2(n2423), 
            .I3(GND_net), .O(n2507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1677_3_lut (.I0(n2391), .I1(n2456[30]), .I2(n2423), 
            .I3(GND_net), .O(n2490));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n2490), .I1(n2489), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_21_22 (.CI(n37234), .I0(bit_ctr[20]), .I1(GND_net), .CO(n37235));
    SB_LUT4 i15_4_lut_adj_1582 (.I0(n2507), .I1(n2503), .I2(n2501), .I3(n2500), 
            .O(n36_adj_4861));
    defparam i15_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_3_lut_adj_1583 (.I0(bit_ctr[10]), .I1(n2499), .I2(n2509), 
            .I3(GND_net), .O(n27_adj_4862));
    defparam i6_3_lut_adj_1583.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1584 (.I0(n2495), .I1(n2497), .I2(n2496), .I3(n2498), 
            .O(n34_adj_4863));
    defparam i13_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1585 (.I0(n2491), .I1(n2493), .I2(n2492), .I3(n2494), 
            .O(n33_adj_4864));
    defparam i12_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1586 (.I0(n2506), .I1(n2508), .I2(n2505), .I3(n22), 
            .O(n37_adj_4865));
    defparam i16_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1587 (.I0(n27_adj_4862), .I1(n36_adj_4861), .I2(n2502), 
            .I3(n2504), .O(n39_adj_4866));
    defparam i18_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n37233), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20_4_lut_adj_1588 (.I0(n39_adj_4866), .I1(n37_adj_4865), .I2(n33_adj_4864), 
            .I3(n34_adj_4863), .O(n2522));
    defparam i20_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_33_lut (.I0(n46398), .I1(timer[31]), .I2(n1[31]), 
            .I3(n37380), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n46396), .I1(timer[30]), .I2(n1[30]), 
            .I3(n37379), .O(n46398)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n37379), .I0(timer[30]), .I1(n1[30]), 
            .CO(n37380));
    SB_LUT4 sub_14_add_2_31_lut (.I0(n46394), .I1(timer[29]), .I2(n1[29]), 
            .I3(n37378), .O(n46396)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n37378), .I0(timer[29]), .I1(n1[29]), 
            .CO(n37379));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n46392), .I1(timer[28]), .I2(n1[28]), 
            .I3(n37377), .O(n46394)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1433), .I1(n1400), .I2(VCC_net), 
            .I3(n37835), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_30 (.CI(n37377), .I0(timer[28]), .I1(n1[28]), 
            .CO(n37378));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(GND_net), .I1(n1401), .I2(VCC_net), 
            .I3(n37834), .O(n1466[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_11 (.CI(n37834), .I0(n1401), .I1(VCC_net), 
            .CO(n37835));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(GND_net), .I1(n1402), .I2(VCC_net), 
            .I3(n37833), .O(n1466[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_21 (.CI(n37233), .I0(bit_ctr[19]), .I1(GND_net), .CO(n37234));
    SB_CARRY mod_5_add_1004_10 (.CI(n37833), .I0(n1402), .I1(VCC_net), 
            .CO(n37834));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(GND_net), .I1(n1403), .I2(VCC_net), 
            .I3(n37832), .O(n1466[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_9 (.CI(n37832), .I0(n1403), .I1(VCC_net), 
            .CO(n37833));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(GND_net), .I1(n1404), .I2(VCC_net), 
            .I3(n37831), .O(n1466[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n37232), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_8 (.CI(n37831), .I0(n1404), .I1(VCC_net), 
            .CO(n37832));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(GND_net), .I1(n1405), .I2(VCC_net), 
            .I3(n37830), .O(n1466[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_7 (.CI(n37830), .I0(n1405), .I1(VCC_net), 
            .CO(n37831));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(GND_net), .I1(n1406), .I2(VCC_net), 
            .I3(n37829), .O(n1466[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1004_6 (.CI(n37829), .I0(n1406), .I1(VCC_net), 
            .CO(n37830));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(GND_net), .I1(n1407), .I2(VCC_net), 
            .I3(n37828), .O(n1466[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1004_5 (.CI(n37828), .I0(n1407), .I1(VCC_net), 
            .CO(n37829));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(GND_net), .I1(n1408), .I2(VCC_net), 
            .I3(n37827), .O(n1466[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_4 (.CI(n37827), .I0(n1408), .I1(VCC_net), 
            .CO(n37828));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(GND_net), .I1(n1409), .I2(GND_net), 
            .I3(n37826), .O(n1466[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_3 (.CI(n37826), .I0(n1409), .I1(GND_net), 
            .CO(n37827));
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n28247));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_29_lut (.I0(n46390), .I1(timer[27]), .I2(n1[27]), 
            .I3(n37376), .O(n46392)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(VCC_net), .O(n1466[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(GND_net), 
            .CO(n37826));
    SB_CARRY add_21_20 (.CI(n37232), .I0(bit_ctr[18]), .I1(GND_net), .CO(n37233));
    SB_LUT4 mod_5_i1625_3_lut (.I0(n2307), .I1(n2357[15]), .I2(n2324), 
            .I3(GND_net), .O(n2406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1619_3_lut (.I0(n2301), .I1(n2357[21]), .I2(n2324), 
            .I3(GND_net), .O(n2400));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1617_3_lut (.I0(n2299), .I1(n2357[23]), .I2(n2324), 
            .I3(GND_net), .O(n2398));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1621_3_lut (.I0(n2303), .I1(n2357[19]), .I2(n2324), 
            .I3(GND_net), .O(n2402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1618_3_lut (.I0(n2300), .I1(n2357[22]), .I2(n2324), 
            .I3(GND_net), .O(n2399));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n37231), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1620_3_lut (.I0(n2302), .I1(n2357[20]), .I2(n2324), 
            .I3(GND_net), .O(n2401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1620_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_19 (.CI(n37231), .I0(bit_ctr[17]), .I1(GND_net), .CO(n37232));
    SB_LUT4 mod_5_i1612_3_lut (.I0(n2294), .I1(n2357[28]), .I2(n2324), 
            .I3(GND_net), .O(n2393));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1611_3_lut (.I0(n2293), .I1(n2357[29]), .I2(n2324), 
            .I3(GND_net), .O(n2392));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1610_3_lut (.I0(n2292), .I1(n2357[30]), .I2(n2324), 
            .I3(GND_net), .O(n2391));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1615_3_lut (.I0(n2297), .I1(n2357[25]), .I2(n2324), 
            .I3(GND_net), .O(n2396));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1614_3_lut (.I0(n2296), .I1(n2357[26]), .I2(n2324), 
            .I3(GND_net), .O(n2395));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1614_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_29 (.CI(n37376), .I0(timer[27]), .I1(n1[27]), 
            .CO(n37377));
    SB_LUT4 sub_14_add_2_28_lut (.I0(n46388), .I1(timer[26]), .I2(n1[26]), 
            .I3(n37375), .O(n46390)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_i1616_3_lut (.I0(n2298), .I1(n2357[24]), .I2(n2324), 
            .I3(GND_net), .O(n2397));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1613_3_lut (.I0(n2295), .I1(n2357[27]), .I2(n2324), 
            .I3(GND_net), .O(n2394));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1613_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_28 (.CI(n37375), .I0(timer[26]), .I1(n1[26]), 
            .CO(n37376));
    SB_LUT4 mod_5_i1628_3_lut (.I0(bit_ctr[12]), .I1(n2357[12]), .I2(n2324), 
            .I3(GND_net), .O(n2409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_27_lut (.I0(n46386), .I1(timer[25]), .I2(n1[25]), 
            .I3(n37374), .O(n46388)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_27 (.CI(n37374), .I0(timer[25]), .I1(n1[25]), 
            .CO(n37375));
    SB_LUT4 mod_5_i1623_3_lut (.I0(n2305), .I1(n2357[17]), .I2(n2324), 
            .I3(GND_net), .O(n2404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1622_3_lut (.I0(n2304), .I1(n2357[18]), .I2(n2324), 
            .I3(GND_net), .O(n2403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_26_lut (.I0(n46384), .I1(timer[24]), .I2(n1[24]), 
            .I3(n37373), .O(n46386)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n37230), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1626_3_lut (.I0(n2308), .I1(n2357[14]), .I2(n2324), 
            .I3(GND_net), .O(n2407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1626_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_26 (.CI(n37373), .I0(timer[24]), .I1(n1[24]), 
            .CO(n37374));
    SB_LUT4 mod_5_i1624_3_lut (.I0(n2306), .I1(n2357[16]), .I2(n2324), 
            .I3(GND_net), .O(n2405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_25_lut (.I0(n46382), .I1(timer[23]), .I2(n1[23]), 
            .I3(n37372), .O(n46384)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_i1627_3_lut (.I0(n2309), .I1(n2357[13]), .I2(n2324), 
            .I3(GND_net), .O(n2408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_1589 (.I0(n2408), .I1(n2405), .I2(n2407), .I3(n2403), 
            .O(n34_adj_4869));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(n2404), .I1(bit_ctr[11]), .I2(n2409), .I3(GND_net), 
            .O(n25_adj_4870));   // verilog/neopixel.v(22[26:36])
    defparam i5_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1590 (.I0(n2394), .I1(n2397), .I2(n2395), .I3(n2396), 
            .O(n32_adj_4871));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2391), .I1(n2392), .I2(n2390), .I3(n2393), 
            .O(n31_adj_4872));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1591 (.I0(n2401), .I1(n2399), .I2(n2402), .I3(n2398), 
            .O(n35_adj_4873));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1592 (.I0(n25_adj_4870), .I1(n34_adj_4869), .I2(n2400), 
            .I3(n2406), .O(n37_adj_4874));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1593 (.I0(n37_adj_4874), .I1(n35_adj_4873), .I2(n31_adj_4872), 
            .I3(n32_adj_4871), .O(n2423));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n28246));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_25 (.CI(n37372), .I0(timer[23]), .I1(n1[23]), 
            .CO(n37373));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1334), .I1(n1301), .I2(VCC_net), 
            .I3(n38307), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_10_lut (.I0(GND_net), .I1(n1302), .I2(VCC_net), 
            .I3(n38306), .O(n1367[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_10 (.CI(n38306), .I0(n1302), .I1(VCC_net), 
            .CO(n38307));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n46380), .I1(timer[22]), .I2(n1[22]), 
            .I3(n37371), .O(n46382)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i19_4_lut_adj_1594 (.I0(bit_ctr[16]), .I1(bit_ctr[24]), .I2(bit_ctr[8]), 
            .I3(bit_ctr[18]), .O(n46_adj_4876));
    defparam i19_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1595 (.I0(bit_ctr[22]), .I1(bit_ctr[6]), .I2(bit_ctr[26]), 
            .I3(bit_ctr[28]), .O(n44_adj_4877));
    defparam i17_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1596 (.I0(bit_ctr[19]), .I1(bit_ctr[23]), .I2(bit_ctr[13]), 
            .I3(bit_ctr[20]), .O(n45_adj_4878));
    defparam i18_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1597 (.I0(bit_ctr[29]), .I1(bit_ctr[21]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[14]), .O(n43_adj_4879));
    defparam i16_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1598 (.I0(bit_ctr[25]), .I1(bit_ctr[17]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[7]), .O(n42_adj_4880));
    defparam i15_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_9_lut (.I0(GND_net), .I1(n1303), .I2(VCC_net), 
            .I3(n38305), .O(n1367[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_3_lut (.I0(bit_ctr[5]), .I1(bit_ctr[12]), .I2(bit_ctr[30]), 
            .I3(GND_net), .O(n41_adj_4881));
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i25_4_lut_adj_1599 (.I0(n43_adj_4879), .I1(n45_adj_4878), .I2(n44_adj_4877), 
            .I3(n46_adj_4876), .O(n52));
    defparam i25_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1600 (.I0(bit_ctr[9]), .I1(bit_ctr[10]), .I2(bit_ctr[27]), 
            .I3(bit_ctr[31]), .O(n47_adj_4882));
    defparam i20_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_24 (.CI(n37371), .I0(timer[22]), .I1(n1[22]), 
            .CO(n37372));
    SB_LUT4 i26_4_lut_adj_1601 (.I0(n47_adj_4882), .I1(n52), .I2(n41_adj_4881), 
            .I3(n42_adj_4880), .O(n40382));
    defparam i26_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1602 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_adj_1602.LUT_INIT = 16'h4444;
    SB_LUT4 i15027_3_lut (.I0(n27723), .I1(n46404), .I2(n11_adj_4883), 
            .I3(GND_net), .O(n28057));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15027_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 sub_14_add_2_23_lut (.I0(n46378), .I1(timer[21]), .I2(n1[21]), 
            .I3(n37370), .O(n46380)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n37370), .I0(timer[21]), .I1(n1[21]), 
            .CO(n37371));
    SB_CARRY mod_5_add_937_9 (.CI(n38305), .I0(n1303), .I1(VCC_net), .CO(n38306));
    SB_LUT4 mod_5_add_937_8_lut (.I0(GND_net), .I1(n1304), .I2(VCC_net), 
            .I3(n38304), .O(n1367[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1603 (.I0(\state[0] ), .I1(n47529), .I2(n47530), 
            .I3(\state[1] ), .O(n12_adj_4884));
    defparam i1_4_lut_adj_1603.LUT_INIT = 16'ha088;
    SB_LUT4 i34296_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49249));
    defparam i34296_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1604 (.I0(n12_adj_4884), .I1(n156), .I2(n14), 
            .I3(\state[1] ), .O(n27723));
    defparam i1_4_lut_adj_1604.LUT_INIT = 16'haaea;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[23]), .I1(n1204), .I2(n1209), .I3(GND_net), 
            .O(n12_adj_4885));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i5_4_lut (.I0(n1205), .I1(n1208), .I2(n1207), .I3(n1206), 
            .O(n13_adj_4886));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n13_adj_4886), .I1(n1203), .I2(n12_adj_4885), 
            .I3(n1202), .O(n1235));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_937_8 (.CI(n38304), .I0(n1304), .I1(VCC_net), .CO(n38305));
    SB_LUT4 mod_5_i1546_3_lut (.I0(n2196), .I1(n2258[27]), .I2(n2225), 
            .I3(GND_net), .O(n2295));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1550_3_lut (.I0(n2200), .I1(n2258[23]), .I2(n2225), 
            .I3(GND_net), .O(n2299));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1550_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n28245));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n28244));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n28243));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n28242));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n28241));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n28240));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n28239));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n28238));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n28237));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n28236));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n28235));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n28234));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n28233));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n28232));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1544_3_lut (.I0(n2194), .I1(n2258[29]), .I2(n2225), 
            .I3(GND_net), .O(n2293));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1545_3_lut (.I0(n2195), .I1(n2258[28]), .I2(n2225), 
            .I3(GND_net), .O(n2294));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1547_3_lut (.I0(n2197), .I1(n2258[26]), .I2(n2225), 
            .I3(GND_net), .O(n2296));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1548_3_lut (.I0(n2198), .I1(n2258[25]), .I2(n2225), 
            .I3(GND_net), .O(n2297));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1551_3_lut (.I0(n2201), .I1(n2258[22]), .I2(n2225), 
            .I3(GND_net), .O(n2300));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1552_3_lut (.I0(n2202), .I1(n2258[21]), .I2(n2225), 
            .I3(GND_net), .O(n2301));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1558_3_lut (.I0(n2208), .I1(n2258[15]), .I2(n2225), 
            .I3(GND_net), .O(n2307));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1557_3_lut (.I0(n2207), .I1(n2258[16]), .I2(n2225), 
            .I3(GND_net), .O(n2306));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1559_3_lut (.I0(n2209), .I1(n2258[14]), .I2(n2225), 
            .I3(GND_net), .O(n2308));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1554_3_lut (.I0(n2204), .I1(n2258[19]), .I2(n2225), 
            .I3(GND_net), .O(n2303));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1555_3_lut (.I0(n2205), .I1(n2258[18]), .I2(n2225), 
            .I3(GND_net), .O(n2304));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1549_3_lut (.I0(n2199), .I1(n2258[24]), .I2(n2225), 
            .I3(GND_net), .O(n2298));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1556_3_lut (.I0(n2206), .I1(n2258[17]), .I2(n2225), 
            .I3(GND_net), .O(n2305));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_937_7_lut (.I0(GND_net), .I1(n1305), .I2(VCC_net), 
            .I3(n38303), .O(n1367[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1543_3_lut (.I0(n2193), .I1(n2258[30]), .I2(n2225), 
            .I3(GND_net), .O(n2292));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1553_3_lut (.I0(n2203), .I1(n2258[20]), .I2(n2225), 
            .I3(GND_net), .O(n2302));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1560_3_lut (.I0(bit_ctr[13]), .I1(n2258[13]), .I2(n2225), 
            .I3(GND_net), .O(n2309));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1605 (.I0(n2294), .I1(n2293), .I2(n2299), .I3(n2295), 
            .O(n30_adj_4887));
    defparam i11_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 i21359_2_lut (.I0(bit_ctr[12]), .I1(n2309), .I2(GND_net), 
            .I3(GND_net), .O(n34405));
    defparam i21359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15_4_lut_adj_1606 (.I0(n2302), .I1(n30_adj_4887), .I2(n2292), 
            .I3(n2291), .O(n34_adj_4888));
    defparam i15_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1607 (.I0(n2305), .I1(n2298), .I2(n2304), .I3(n2303), 
            .O(n32_adj_4889));
    defparam i13_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1608 (.I0(n2308), .I1(n34405), .I2(n2306), .I3(n2307), 
            .O(n33_adj_4890));
    defparam i14_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1609 (.I0(n2301), .I1(n2300), .I2(n2297), .I3(n2296), 
            .O(n31_adj_4891));
    defparam i12_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1610 (.I0(n31_adj_4891), .I1(n33_adj_4890), .I2(n32_adj_4889), 
            .I3(n34_adj_4888), .O(n2324));
    defparam i18_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_18 (.CI(n37230), .I0(bit_ctr[16]), .I1(GND_net), .CO(n37231));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n46376), .I1(timer[20]), .I2(n1[20]), 
            .I3(n37369), .O(n46378)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i2_2_lut_adj_1611 (.I0(one_wire_N_579[3]), .I1(n4_adj_4893), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/neopixel.v(6[16:24])
    defparam i2_2_lut_adj_1611.LUT_INIT = 16'h8888;
    SB_LUT4 i28128_2_lut (.I0(\state[1] ), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n43000));
    defparam i28128_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1612 (.I0(one_wire_N_579[3]), .I1(one_wire_N_579[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4823));
    defparam i1_2_lut_adj_1612.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1613 (.I0(one_wire_N_579[8]), .I1(n46352), .I2(GND_net), 
            .I3(GND_net), .O(n46354));
    defparam i1_2_lut_adj_1613.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(one_wire_N_579[10]), .I1(n160), .I2(one_wire_N_579[9]), 
            .I3(n46354), .O(n147));
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1615 (.I0(n45), .I1(n30298), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n29_adj_4894));
    defparam i1_4_lut_adj_1615.LUT_INIT = 16'h3553;
    SB_LUT4 i33565_2_lut (.I0(n29_adj_4894), .I1(n43000), .I2(GND_net), 
            .I3(GND_net), .O(n42167));
    defparam i33565_2_lut.LUT_INIT = 16'hdddd;
    SB_CARRY sub_14_add_2_22 (.CI(n37369), .I0(timer[20]), .I1(n1[20]), 
            .CO(n37370));
    SB_LUT4 i17276_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_636 ));   // verilog/neopixel.v(16[20:25])
    defparam i17276_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n37229), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_17 (.CI(n37229), .I0(bit_ctr[15]), .I1(GND_net), .CO(n37230));
    SB_CARRY mod_5_add_937_7 (.CI(n38303), .I0(n1305), .I1(VCC_net), .CO(n38304));
    SB_LUT4 mod_5_add_937_6_lut (.I0(GND_net), .I1(n1306), .I2(VCC_net), 
            .I3(n38302), .O(n1367[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_21_lut (.I0(n46374), .I1(timer[19]), .I2(n1[19]), 
            .I3(n37368), .O(n46376)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_21 (.CI(n37368), .I0(timer[19]), .I1(n1[19]), 
            .CO(n37369));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n48865), .I1(n48865), .I2(n1037), 
            .I3(n39004), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_20_lut (.I0(n46372), .I1(timer[18]), .I2(n1[18]), 
            .I3(n37367), .O(n46374)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n48792), .I1(n48792), .I2(n1037), 
            .I3(n39003), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n38302), .I0(n1306), .I1(VCC_net), .CO(n38303));
    SB_LUT4 mod_5_add_937_5_lut (.I0(GND_net), .I1(n1307), .I2(VCC_net), 
            .I3(n38301), .O(n1367[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_5 (.CI(n38301), .I0(n1307), .I1(VCC_net), .CO(n38302));
    SB_CARRY sub_14_add_2_20 (.CI(n37367), .I0(timer[18]), .I1(n1[18]), 
            .CO(n37368));
    SB_CARRY mod_5_add_736_7 (.CI(n39003), .I0(n48792), .I1(n1037), .CO(n39004));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n48737), .I1(n1006), .I2(n1037), 
            .I3(n39002), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n39002), .I0(n1006), .I1(n1037), .CO(n39003));
    SB_LUT4 mod_5_add_937_4_lut (.I0(GND_net), .I1(n1308), .I2(VCC_net), 
            .I3(n38300), .O(n1367[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_736_5_lut (.I0(n48738), .I1(n1007), .I2(n1037), 
            .I3(n39001), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n38300), .I0(n1308), .I1(VCC_net), .CO(n38301));
    SB_CARRY mod_5_add_736_5 (.CI(n39001), .I0(n1007), .I1(n1037), .CO(n39002));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n39000), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n39000), .I0(n1008), .I1(n1037), .CO(n39001));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n49244), 
            .I3(n38999), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n38999), .I0(n1009), .I1(n49244), .CO(n39000));
    SB_LUT4 mod_5_add_937_3_lut (.I0(GND_net), .I1(n1309), .I2(GND_net), 
            .I3(n38299), .O(n1367[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n37228), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n49244), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n49244), 
            .CO(n38999));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n38998), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n38997), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n38997), .I0(n1104), .I1(n1136), .CO(n38998));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n38996), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n38996), .I0(n1105), .I1(n1136), .CO(n38997));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n38995), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n38995), .I0(n1106), .I1(n1136), .CO(n38996));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n38994), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n38994), .I0(n1107), .I1(n1136), .CO(n38995));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n38993), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n38993), .I0(n1108), .I1(n1136), .CO(n38994));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n49245), 
            .I3(n38992), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n38992), .I0(n1109), .I1(n49245), .CO(n38993));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n49245), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n49245), 
            .CO(n38992));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1631), .I1(n1598), .I2(VCC_net), 
            .I3(n38991), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(GND_net), .I1(n1599), .I2(VCC_net), 
            .I3(n38990), .O(n1664[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_13 (.CI(n38990), .I0(n1599), .I1(VCC_net), 
            .CO(n38991));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(GND_net), .I1(n1600), .I2(VCC_net), 
            .I3(n38989), .O(n1664[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_12 (.CI(n38989), .I0(n1600), .I1(VCC_net), 
            .CO(n38990));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(GND_net), .I1(n1601), .I2(VCC_net), 
            .I3(n38988), .O(n1664[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_11 (.CI(n38988), .I0(n1601), .I1(VCC_net), 
            .CO(n38989));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(GND_net), .I1(n1602), .I2(VCC_net), 
            .I3(n38987), .O(n1664[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_3 (.CI(n38299), .I0(n1309), .I1(GND_net), .CO(n38300));
    SB_CARRY mod_5_add_1138_10 (.CI(n38987), .I0(n1602), .I1(VCC_net), 
            .CO(n38988));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(GND_net), .I1(n1603), .I2(VCC_net), 
            .I3(n38986), .O(n1664[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_9 (.CI(n38986), .I0(n1603), .I1(VCC_net), 
            .CO(n38987));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(GND_net), .I1(n1604), .I2(VCC_net), 
            .I3(n38985), .O(n1664[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_8 (.CI(n38985), .I0(n1604), .I1(VCC_net), 
            .CO(n38986));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(GND_net), .I1(n1605), .I2(VCC_net), 
            .I3(n38984), .O(n1664[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_19_lut (.I0(n46370), .I1(timer[17]), .I2(n1[17]), 
            .I3(n37366), .O(n46372)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1138_7 (.CI(n38984), .I0(n1605), .I1(VCC_net), 
            .CO(n38985));
    SB_LUT4 mod_5_add_937_2_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(VCC_net), .O(n1367[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(GND_net), 
            .CO(n38299));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(GND_net), .I1(n1606), .I2(VCC_net), 
            .I3(n38983), .O(n1664[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_6 (.CI(n38983), .I0(n1606), .I1(VCC_net), 
            .CO(n38984));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(GND_net), .I1(n1607), .I2(VCC_net), 
            .I3(n38982), .O(n1664[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_5 (.CI(n38982), .I0(n1607), .I1(VCC_net), 
            .CO(n38983));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(GND_net), .I1(n1608), .I2(VCC_net), 
            .I3(n38981), .O(n1664[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_4 (.CI(n38981), .I0(n1608), .I1(VCC_net), 
            .CO(n38982));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(GND_net), .I1(n1609), .I2(GND_net), 
            .I3(n38980), .O(n1664[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_3 (.CI(n38980), .I0(n1609), .I1(GND_net), 
            .CO(n38981));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(VCC_net), .O(n1664[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(GND_net), 
            .CO(n38980));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1730), .I1(n1697), .I2(VCC_net), 
            .I3(n38979), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(GND_net), .I1(n1698), .I2(VCC_net), 
            .I3(n38978), .O(n1763[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_14 (.CI(n38978), .I0(n1698), .I1(VCC_net), 
            .CO(n38979));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(GND_net), .I1(n1699), .I2(VCC_net), 
            .I3(n38977), .O(n1763[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_13 (.CI(n38977), .I0(n1699), .I1(VCC_net), 
            .CO(n38978));
    SB_CARRY sub_14_add_2_19 (.CI(n37366), .I0(timer[17]), .I1(n1[17]), 
            .CO(n37367));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(GND_net), .I1(n1700), .I2(VCC_net), 
            .I3(n38976), .O(n1763[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_12 (.CI(n38976), .I0(n1700), .I1(VCC_net), 
            .CO(n38977));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(GND_net), .I1(n1701), .I2(VCC_net), 
            .I3(n38975), .O(n1763[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_11 (.CI(n38975), .I0(n1701), .I1(VCC_net), 
            .CO(n38976));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(GND_net), .I1(n1702), .I2(VCC_net), 
            .I3(n38974), .O(n1763[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_10 (.CI(n38974), .I0(n1702), .I1(VCC_net), 
            .CO(n38975));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(GND_net), .I1(n1703), .I2(VCC_net), 
            .I3(n38973), .O(n1763[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_9 (.CI(n38973), .I0(n1703), .I1(VCC_net), 
            .CO(n38974));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(GND_net), .I1(n1704), .I2(VCC_net), 
            .I3(n38972), .O(n1763[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_8 (.CI(n38972), .I0(n1704), .I1(VCC_net), 
            .CO(n38973));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(GND_net), .I1(n1705), .I2(VCC_net), 
            .I3(n38971), .O(n1763[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_7 (.CI(n38971), .I0(n1705), .I1(VCC_net), 
            .CO(n38972));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(GND_net), .I1(n1706), .I2(VCC_net), 
            .I3(n38970), .O(n1763[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_6 (.CI(n38970), .I0(n1706), .I1(VCC_net), 
            .CO(n38971));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(GND_net), .I1(n1707), .I2(VCC_net), 
            .I3(n38969), .O(n1763[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_5 (.CI(n38969), .I0(n1707), .I1(VCC_net), 
            .CO(n38970));
    SB_LUT4 sub_14_add_2_18_lut (.I0(n46368), .I1(timer[16]), .I2(n1[16]), 
            .I3(n37365), .O(n46370)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(GND_net), .I1(n1708), .I2(VCC_net), 
            .I3(n38968), .O(n1763[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_4 (.CI(n38968), .I0(n1708), .I1(VCC_net), 
            .CO(n38969));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(GND_net), .I1(n1709), .I2(GND_net), 
            .I3(n38967), .O(n1763[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_3 (.CI(n38967), .I0(n1709), .I1(GND_net), 
            .CO(n38968));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(VCC_net), .O(n1763[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(GND_net), 
            .CO(n38967));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1829), .I1(n1796), .I2(VCC_net), 
            .I3(n38966), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(GND_net), .I1(n1797), .I2(VCC_net), 
            .I3(n38965), .O(n1862[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_15 (.CI(n38965), .I0(n1797), .I1(VCC_net), 
            .CO(n38966));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(GND_net), .I1(n1798), .I2(VCC_net), 
            .I3(n38964), .O(n1862[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_14 (.CI(n38964), .I0(n1798), .I1(VCC_net), 
            .CO(n38965));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(GND_net), .I1(n1799), .I2(VCC_net), 
            .I3(n38963), .O(n1862[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_13 (.CI(n38963), .I0(n1799), .I1(VCC_net), 
            .CO(n38964));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(GND_net), .I1(n1800), .I2(VCC_net), 
            .I3(n38962), .O(n1862[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_12 (.CI(n38962), .I0(n1800), .I1(VCC_net), 
            .CO(n38963));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(GND_net), .I1(n1801), .I2(VCC_net), 
            .I3(n38961), .O(n1862[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_11 (.CI(n38961), .I0(n1801), .I1(VCC_net), 
            .CO(n38962));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(GND_net), .I1(n1802), .I2(VCC_net), 
            .I3(n38960), .O(n1862[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_10 (.CI(n38960), .I0(n1802), .I1(VCC_net), 
            .CO(n38961));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(GND_net), .I1(n1803), .I2(VCC_net), 
            .I3(n38959), .O(n1862[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_9 (.CI(n38959), .I0(n1803), .I1(VCC_net), 
            .CO(n38960));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(GND_net), .I1(n1804), .I2(VCC_net), 
            .I3(n38958), .O(n1862[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_8 (.CI(n38958), .I0(n1804), .I1(VCC_net), 
            .CO(n38959));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(GND_net), .I1(n1805), .I2(VCC_net), 
            .I3(n38957), .O(n1862[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_7 (.CI(n38957), .I0(n1805), .I1(VCC_net), 
            .CO(n38958));
    SB_CARRY add_21_16 (.CI(n37228), .I0(bit_ctr[14]), .I1(GND_net), .CO(n37229));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(GND_net), .I1(n1806), .I2(VCC_net), 
            .I3(n38956), .O(n1862[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_6 (.CI(n38956), .I0(n1806), .I1(VCC_net), 
            .CO(n38957));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(GND_net), .I1(n1807), .I2(VCC_net), 
            .I3(n38955), .O(n1862[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_5 (.CI(n38955), .I0(n1807), .I1(VCC_net), 
            .CO(n38956));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(GND_net), .I1(n1808), .I2(VCC_net), 
            .I3(n38954), .O(n1862[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_4 (.CI(n38954), .I0(n1808), .I1(VCC_net), 
            .CO(n38955));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(GND_net), .I1(n1809), .I2(GND_net), 
            .I3(n38953), .O(n1862[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_3 (.CI(n38953), .I0(n1809), .I1(GND_net), 
            .CO(n38954));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(VCC_net), .O(n1862[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(GND_net), 
            .CO(n38953));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1928), .I1(n1895), .I2(VCC_net), 
            .I3(n38952), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(GND_net), .I1(n1896), .I2(VCC_net), 
            .I3(n38951), .O(n1961[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_16 (.CI(n38951), .I0(n1896), .I1(VCC_net), 
            .CO(n38952));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(GND_net), .I1(n1897), .I2(VCC_net), 
            .I3(n38950), .O(n1961[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_15 (.CI(n38950), .I0(n1897), .I1(VCC_net), 
            .CO(n38951));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(GND_net), .I1(n1898), .I2(VCC_net), 
            .I3(n38949), .O(n1961[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_14 (.CI(n38949), .I0(n1898), .I1(VCC_net), 
            .CO(n38950));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(GND_net), .I1(n1899), .I2(VCC_net), 
            .I3(n38948), .O(n1961[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_13 (.CI(n38948), .I0(n1899), .I1(VCC_net), 
            .CO(n38949));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(GND_net), .I1(n1900), .I2(VCC_net), 
            .I3(n38947), .O(n1961[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_12 (.CI(n38947), .I0(n1900), .I1(VCC_net), 
            .CO(n38948));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(GND_net), .I1(n1901), .I2(VCC_net), 
            .I3(n38946), .O(n1961[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_11 (.CI(n38946), .I0(n1901), .I1(VCC_net), 
            .CO(n38947));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(GND_net), .I1(n1902), .I2(VCC_net), 
            .I3(n38945), .O(n1961[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_10 (.CI(n38945), .I0(n1902), .I1(VCC_net), 
            .CO(n38946));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(GND_net), .I1(n1903), .I2(VCC_net), 
            .I3(n38944), .O(n1961[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_9 (.CI(n38944), .I0(n1903), .I1(VCC_net), 
            .CO(n38945));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(GND_net), .I1(n1904), .I2(VCC_net), 
            .I3(n38943), .O(n1961[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_8 (.CI(n38943), .I0(n1904), .I1(VCC_net), 
            .CO(n38944));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(GND_net), .I1(n1905), .I2(VCC_net), 
            .I3(n38942), .O(n1961[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_7 (.CI(n38942), .I0(n1905), .I1(VCC_net), 
            .CO(n38943));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(GND_net), .I1(n1906), .I2(VCC_net), 
            .I3(n38941), .O(n1961[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_6 (.CI(n38941), .I0(n1906), .I1(VCC_net), 
            .CO(n38942));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(GND_net), .I1(n1907), .I2(VCC_net), 
            .I3(n38940), .O(n1961[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_5 (.CI(n38940), .I0(n1907), .I1(VCC_net), 
            .CO(n38941));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(GND_net), .I1(n1908), .I2(VCC_net), 
            .I3(n38939), .O(n1961[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_4 (.CI(n38939), .I0(n1908), .I1(VCC_net), 
            .CO(n38940));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(GND_net), .I1(n1909), .I2(GND_net), 
            .I3(n38938), .O(n1961[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_3 (.CI(n38938), .I0(n1909), .I1(GND_net), 
            .CO(n38939));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(VCC_net), .O(n1961[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(GND_net), 
            .CO(n38938));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n2027), .I1(n1994), .I2(VCC_net), 
            .I3(n38937), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(GND_net), .I1(n1995), .I2(VCC_net), 
            .I3(n38936), .O(n2060[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_17 (.CI(n38936), .I0(n1995), .I1(VCC_net), 
            .CO(n38937));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(GND_net), .I1(n1996), .I2(VCC_net), 
            .I3(n38935), .O(n2060[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n37365), .I0(timer[16]), .I1(n1[16]), 
            .CO(n37366));
    SB_CARRY mod_5_add_1406_16 (.CI(n38935), .I0(n1996), .I1(VCC_net), 
            .CO(n38936));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(GND_net), .I1(n1997), .I2(VCC_net), 
            .I3(n38934), .O(n2060[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_15 (.CI(n38934), .I0(n1997), .I1(VCC_net), 
            .CO(n38935));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(GND_net), .I1(n1998), .I2(VCC_net), 
            .I3(n38933), .O(n2060[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_14 (.CI(n38933), .I0(n1998), .I1(VCC_net), 
            .CO(n38934));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(GND_net), .I1(n1999), .I2(VCC_net), 
            .I3(n38932), .O(n2060[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_13 (.CI(n38932), .I0(n1999), .I1(VCC_net), 
            .CO(n38933));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(GND_net), .I1(n2000), .I2(VCC_net), 
            .I3(n38931), .O(n2060[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_12 (.CI(n38931), .I0(n2000), .I1(VCC_net), 
            .CO(n38932));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(GND_net), .I1(n2001), .I2(VCC_net), 
            .I3(n38930), .O(n2060[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_11 (.CI(n38930), .I0(n2001), .I1(VCC_net), 
            .CO(n38931));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(GND_net), .I1(n2002), .I2(VCC_net), 
            .I3(n38929), .O(n2060[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_10 (.CI(n38929), .I0(n2002), .I1(VCC_net), 
            .CO(n38930));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(GND_net), .I1(n2003), .I2(VCC_net), 
            .I3(n38928), .O(n2060[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_9 (.CI(n38928), .I0(n2003), .I1(VCC_net), 
            .CO(n38929));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(GND_net), .I1(n2004), .I2(VCC_net), 
            .I3(n38927), .O(n2060[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_8 (.CI(n38927), .I0(n2004), .I1(VCC_net), 
            .CO(n38928));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(GND_net), .I1(n2005), .I2(VCC_net), 
            .I3(n38926), .O(n2060[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_7 (.CI(n38926), .I0(n2005), .I1(VCC_net), 
            .CO(n38927));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(GND_net), .I1(n2006), .I2(VCC_net), 
            .I3(n38925), .O(n2060[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_6 (.CI(n38925), .I0(n2006), .I1(VCC_net), 
            .CO(n38926));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(GND_net), .I1(n2007), .I2(VCC_net), 
            .I3(n38924), .O(n2060[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_5 (.CI(n38924), .I0(n2007), .I1(VCC_net), 
            .CO(n38925));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(GND_net), .I1(n2008), .I2(VCC_net), 
            .I3(n38923), .O(n2060[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_4 (.CI(n38923), .I0(n2008), .I1(VCC_net), 
            .CO(n38924));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(GND_net), .I1(n2009), .I2(GND_net), 
            .I3(n38922), .O(n2060[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_3 (.CI(n38922), .I0(n2009), .I1(GND_net), 
            .CO(n38923));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(VCC_net), .O(n2060[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(GND_net), 
            .CO(n38922));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2126), .I1(n2093), .I2(VCC_net), 
            .I3(n38921), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(GND_net), .I1(n2094), .I2(VCC_net), 
            .I3(n38920), .O(n2159[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_17_lut (.I0(n46366), .I1(timer[15]), .I2(n1[15]), 
            .I3(n37364), .O(n46368)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_17 (.CI(n37364), .I0(timer[15]), .I1(n1[15]), 
            .CO(n37365));
    SB_CARRY mod_5_add_1473_18 (.CI(n38920), .I0(n2094), .I1(VCC_net), 
            .CO(n38921));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(GND_net), .I1(n2095), .I2(VCC_net), 
            .I3(n38919), .O(n2159[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_17 (.CI(n38919), .I0(n2095), .I1(VCC_net), 
            .CO(n38920));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(GND_net), .I1(n2096), .I2(VCC_net), 
            .I3(n38918), .O(n2159[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_16 (.CI(n38918), .I0(n2096), .I1(VCC_net), 
            .CO(n38919));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(GND_net), .I1(n2097), .I2(VCC_net), 
            .I3(n38917), .O(n2159[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_15 (.CI(n38917), .I0(n2097), .I1(VCC_net), 
            .CO(n38918));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(GND_net), .I1(n2098), .I2(VCC_net), 
            .I3(n38916), .O(n2159[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_14 (.CI(n38916), .I0(n2098), .I1(VCC_net), 
            .CO(n38917));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(GND_net), .I1(n2099), .I2(VCC_net), 
            .I3(n38915), .O(n2159[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_13 (.CI(n38915), .I0(n2099), .I1(VCC_net), 
            .CO(n38916));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(GND_net), .I1(n2100), .I2(VCC_net), 
            .I3(n38914), .O(n2159[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_12 (.CI(n38914), .I0(n2100), .I1(VCC_net), 
            .CO(n38915));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(GND_net), .I1(n2101), .I2(VCC_net), 
            .I3(n38913), .O(n2159[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_11 (.CI(n38913), .I0(n2101), .I1(VCC_net), 
            .CO(n38914));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(GND_net), .I1(n2102), .I2(VCC_net), 
            .I3(n38912), .O(n2159[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_10 (.CI(n38912), .I0(n2102), .I1(VCC_net), 
            .CO(n38913));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(GND_net), .I1(n2103), .I2(VCC_net), 
            .I3(n38911), .O(n2159[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_9 (.CI(n38911), .I0(n2103), .I1(VCC_net), 
            .CO(n38912));
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(GND_net), .I1(n2104), .I2(VCC_net), 
            .I3(n38910), .O(n2159[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_8 (.CI(n38910), .I0(n2104), .I1(VCC_net), 
            .CO(n38911));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(GND_net), .I1(n2105), .I2(VCC_net), 
            .I3(n38909), .O(n2159[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_7 (.CI(n38909), .I0(n2105), .I1(VCC_net), 
            .CO(n38910));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(GND_net), .I1(n2106), .I2(VCC_net), 
            .I3(n38908), .O(n2159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(CLK_c), .E(VCC_net), .D(n12));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1473_6 (.CI(n38908), .I0(n2106), .I1(VCC_net), 
            .CO(n38909));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(GND_net), .I1(n2107), .I2(VCC_net), 
            .I3(n38907), .O(n2159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_5 (.CI(n38907), .I0(n2107), .I1(VCC_net), 
            .CO(n38908));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(GND_net), .I1(n2108), .I2(VCC_net), 
            .I3(n38906), .O(n2159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_4 (.CI(n38906), .I0(n2108), .I1(VCC_net), 
            .CO(n38907));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(GND_net), .I1(n2109), .I2(GND_net), 
            .I3(n38905), .O(n2159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_3 (.CI(n38905), .I0(n2109), .I1(GND_net), 
            .CO(n38906));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(VCC_net), .O(n2159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(GND_net), 
            .CO(n38905));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2225), .I1(n2192), .I2(VCC_net), 
            .I3(n38904), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(GND_net), .I1(n2193), .I2(VCC_net), 
            .I3(n38903), .O(n2258[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_19 (.CI(n38903), .I0(n2193), .I1(VCC_net), 
            .CO(n38904));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(GND_net), .I1(n2194), .I2(VCC_net), 
            .I3(n38902), .O(n2258[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_18 (.CI(n38902), .I0(n2194), .I1(VCC_net), 
            .CO(n38903));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(GND_net), .I1(n2195), .I2(VCC_net), 
            .I3(n38901), .O(n2258[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_17 (.CI(n38901), .I0(n2195), .I1(VCC_net), 
            .CO(n38902));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(GND_net), .I1(n2196), .I2(VCC_net), 
            .I3(n38900), .O(n2258[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_16 (.CI(n38900), .I0(n2196), .I1(VCC_net), 
            .CO(n38901));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(GND_net), .I1(n2197), .I2(VCC_net), 
            .I3(n38899), .O(n2258[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_15 (.CI(n38899), .I0(n2197), .I1(VCC_net), 
            .CO(n38900));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(GND_net), .I1(n2198), .I2(VCC_net), 
            .I3(n38898), .O(n2258[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_16_lut (.I0(n46364), .I1(timer[14]), .I2(n1[14]), 
            .I3(n37363), .O(n46366)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n37363), .I0(timer[14]), .I1(n1[14]), 
            .CO(n37364));
    SB_CARRY mod_5_add_1540_14 (.CI(n38898), .I0(n2198), .I1(VCC_net), 
            .CO(n38899));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(GND_net), .I1(n2199), .I2(VCC_net), 
            .I3(n38897), .O(n2258[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_15_lut (.I0(n46362), .I1(timer[13]), .I2(n1[13]), 
            .I3(n37362), .O(n46364)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1540_13 (.CI(n38897), .I0(n2199), .I1(VCC_net), 
            .CO(n38898));
    SB_DFF timer_1547__i0 (.Q(timer[0]), .C(CLK_c), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1540_12_lut (.I0(GND_net), .I1(n2200), .I2(VCC_net), 
            .I3(n38896), .O(n2258[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_12 (.CI(n38896), .I0(n2200), .I1(VCC_net), 
            .CO(n38897));
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n49521));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49521_bdd_4_lut (.I0(n49521), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n49524));
    defparam n49521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1540_11_lut (.I0(GND_net), .I1(n2201), .I2(VCC_net), 
            .I3(n38895), .O(n2258[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_11 (.CI(n38895), .I0(n2201), .I1(VCC_net), 
            .CO(n38896));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(GND_net), .I1(n2202), .I2(VCC_net), 
            .I3(n38894), .O(n2258[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_10 (.CI(n38894), .I0(n2202), .I1(VCC_net), 
            .CO(n38895));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(GND_net), .I1(n2203), .I2(VCC_net), 
            .I3(n38893), .O(n2258[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_9 (.CI(n38893), .I0(n2203), .I1(VCC_net), 
            .CO(n38894));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(GND_net), .I1(n2204), .I2(VCC_net), 
            .I3(n38892), .O(n2258[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_8 (.CI(n38892), .I0(n2204), .I1(VCC_net), 
            .CO(n38893));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(GND_net), .I1(n2205), .I2(VCC_net), 
            .I3(n38891), .O(n2258[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_7 (.CI(n38891), .I0(n2205), .I1(VCC_net), 
            .CO(n38892));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(GND_net), .I1(n2206), .I2(VCC_net), 
            .I3(n38890), .O(n2258[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_6 (.CI(n38890), .I0(n2206), .I1(VCC_net), 
            .CO(n38891));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(GND_net), .I1(n2207), .I2(VCC_net), 
            .I3(n38889), .O(n2258[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_5 (.CI(n38889), .I0(n2207), .I1(VCC_net), 
            .CO(n38890));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(GND_net), .I1(n2208), .I2(VCC_net), 
            .I3(n38888), .O(n2258[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_4 (.CI(n38888), .I0(n2208), .I1(VCC_net), 
            .CO(n38889));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(GND_net), .I1(n2209), .I2(GND_net), 
            .I3(n38887), .O(n2258[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_3 (.CI(n38887), .I0(n2209), .I1(GND_net), 
            .CO(n38888));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(VCC_net), .O(n2258[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(GND_net), 
            .CO(n38887));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2324), .I1(n2291), .I2(VCC_net), 
            .I3(n38886), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(GND_net), .I1(n2292), .I2(VCC_net), 
            .I3(n38885), .O(n2357[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_20 (.CI(n38885), .I0(n2292), .I1(VCC_net), 
            .CO(n38886));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(GND_net), .I1(n2293), .I2(VCC_net), 
            .I3(n38884), .O(n2357[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n37227), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_19 (.CI(n38884), .I0(n2293), .I1(VCC_net), 
            .CO(n38885));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(GND_net), .I1(n2294), .I2(VCC_net), 
            .I3(n38883), .O(n2357[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_18 (.CI(n38883), .I0(n2294), .I1(VCC_net), 
            .CO(n38884));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(GND_net), .I1(n2295), .I2(VCC_net), 
            .I3(n38882), .O(n2357[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_17 (.CI(n38882), .I0(n2295), .I1(VCC_net), 
            .CO(n38883));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(GND_net), .I1(n2296), .I2(VCC_net), 
            .I3(n38881), .O(n2357[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_16 (.CI(n38881), .I0(n2296), .I1(VCC_net), 
            .CO(n38882));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(GND_net), .I1(n2297), .I2(VCC_net), 
            .I3(n38880), .O(n2357[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_15 (.CI(n38880), .I0(n2297), .I1(VCC_net), 
            .CO(n38881));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(GND_net), .I1(n2298), .I2(VCC_net), 
            .I3(n38879), .O(n2357[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_14 (.CI(n38879), .I0(n2298), .I1(VCC_net), 
            .CO(n38880));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(GND_net), .I1(n2299), .I2(VCC_net), 
            .I3(n38878), .O(n2357[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_13 (.CI(n38878), .I0(n2299), .I1(VCC_net), 
            .CO(n38879));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(GND_net), .I1(n2300), .I2(VCC_net), 
            .I3(n38877), .O(n2357[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_12 (.CI(n38877), .I0(n2300), .I1(VCC_net), 
            .CO(n38878));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(GND_net), .I1(n2301), .I2(VCC_net), 
            .I3(n38876), .O(n2357[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_11 (.CI(n38876), .I0(n2301), .I1(VCC_net), 
            .CO(n38877));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(GND_net), .I1(n2302), .I2(VCC_net), 
            .I3(n38875), .O(n2357[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n38875), .I0(n2302), .I1(VCC_net), 
            .CO(n38876));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(GND_net), .I1(n2303), .I2(VCC_net), 
            .I3(n38874), .O(n2357[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_9 (.CI(n38874), .I0(n2303), .I1(VCC_net), 
            .CO(n38875));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(GND_net), .I1(n2304), .I2(VCC_net), 
            .I3(n38873), .O(n2357[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_8 (.CI(n38873), .I0(n2304), .I1(VCC_net), 
            .CO(n38874));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(GND_net), .I1(n2305), .I2(VCC_net), 
            .I3(n38872), .O(n2357[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_7 (.CI(n38872), .I0(n2305), .I1(VCC_net), 
            .CO(n38873));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(GND_net), .I1(n2306), .I2(VCC_net), 
            .I3(n38871), .O(n2357[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_6 (.CI(n38871), .I0(n2306), .I1(VCC_net), 
            .CO(n38872));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(GND_net), .I1(n2307), .I2(VCC_net), 
            .I3(n38870), .O(n2357[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_5 (.CI(n38870), .I0(n2307), .I1(VCC_net), 
            .CO(n38871));
    SB_CARRY sub_14_add_2_15 (.CI(n37362), .I0(timer[13]), .I1(n1[13]), 
            .CO(n37363));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(GND_net), .I1(n2308), .I2(VCC_net), 
            .I3(n38869), .O(n2357[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_4 (.CI(n38869), .I0(n2308), .I1(VCC_net), 
            .CO(n38870));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(GND_net), .I1(n2309), .I2(GND_net), 
            .I3(n38868), .O(n2357[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_3 (.CI(n38868), .I0(n2309), .I1(GND_net), 
            .CO(n38869));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(VCC_net), .O(n2357[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(GND_net), 
            .CO(n38868));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2423), .I1(n2390), .I2(VCC_net), 
            .I3(n38867), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(GND_net), .I1(n2391), .I2(VCC_net), 
            .I3(n38866), .O(n2456[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_21 (.CI(n38866), .I0(n2391), .I1(VCC_net), 
            .CO(n38867));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(GND_net), .I1(n2392), .I2(VCC_net), 
            .I3(n38865), .O(n2456[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_20 (.CI(n38865), .I0(n2392), .I1(VCC_net), 
            .CO(n38866));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(GND_net), .I1(n2393), .I2(VCC_net), 
            .I3(n38864), .O(n2456[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_19 (.CI(n38864), .I0(n2393), .I1(VCC_net), 
            .CO(n38865));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(GND_net), .I1(n2394), .I2(VCC_net), 
            .I3(n38863), .O(n2456[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_18 (.CI(n38863), .I0(n2394), .I1(VCC_net), 
            .CO(n38864));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(GND_net), .I1(n2395), .I2(VCC_net), 
            .I3(n38862), .O(n2456[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_17 (.CI(n38862), .I0(n2395), .I1(VCC_net), 
            .CO(n38863));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(GND_net), .I1(n2396), .I2(VCC_net), 
            .I3(n38861), .O(n2456[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_16 (.CI(n38861), .I0(n2396), .I1(VCC_net), 
            .CO(n38862));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(GND_net), .I1(n2397), .I2(VCC_net), 
            .I3(n38860), .O(n2456[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_15 (.CI(n38860), .I0(n2397), .I1(VCC_net), 
            .CO(n38861));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(GND_net), .I1(n2398), .I2(VCC_net), 
            .I3(n38859), .O(n2456[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_14 (.CI(n38859), .I0(n2398), .I1(VCC_net), 
            .CO(n38860));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(GND_net), .I1(n2399), .I2(VCC_net), 
            .I3(n38858), .O(n2456[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_13 (.CI(n38858), .I0(n2399), .I1(VCC_net), 
            .CO(n38859));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(GND_net), .I1(n2400), .I2(VCC_net), 
            .I3(n38857), .O(n2456[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_12 (.CI(n38857), .I0(n2400), .I1(VCC_net), 
            .CO(n38858));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(GND_net), .I1(n2401), .I2(VCC_net), 
            .I3(n38856), .O(n2456[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_11 (.CI(n38856), .I0(n2401), .I1(VCC_net), 
            .CO(n38857));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(GND_net), .I1(n2402), .I2(VCC_net), 
            .I3(n38855), .O(n2456[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_10 (.CI(n38855), .I0(n2402), .I1(VCC_net), 
            .CO(n38856));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(GND_net), .I1(n2403), .I2(VCC_net), 
            .I3(n38854), .O(n2456[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n38854), .I0(n2403), .I1(VCC_net), 
            .CO(n38855));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_579[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n37361), .O(n46362)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_14 (.CI(n37361), .I0(timer[12]), .I1(n1[12]), 
            .CO(n37362));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(GND_net), .I1(n2404), .I2(VCC_net), 
            .I3(n38853), .O(n2456[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_8 (.CI(n38853), .I0(n2404), .I1(VCC_net), 
            .CO(n38854));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n37360), .O(one_wire_N_579[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_15 (.CI(n37227), .I0(bit_ctr[13]), .I1(GND_net), .CO(n37228));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(GND_net), .I1(n2405), .I2(VCC_net), 
            .I3(n38852), .O(n2456[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_7 (.CI(n38852), .I0(n2405), .I1(VCC_net), 
            .CO(n38853));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(GND_net), .I1(n2406), .I2(VCC_net), 
            .I3(n38851), .O(n2456[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_6 (.CI(n38851), .I0(n2406), .I1(VCC_net), 
            .CO(n38852));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(GND_net), .I1(n2407), .I2(VCC_net), 
            .I3(n38850), .O(n2456[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_5 (.CI(n38850), .I0(n2407), .I1(VCC_net), 
            .CO(n38851));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(GND_net), .I1(n2408), .I2(VCC_net), 
            .I3(n38849), .O(n2456[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_4 (.CI(n38849), .I0(n2408), .I1(VCC_net), 
            .CO(n38850));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(GND_net), .I1(n2409), .I2(GND_net), 
            .I3(n38848), .O(n2456[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_3 (.CI(n38848), .I0(n2409), .I1(GND_net), 
            .CO(n38849));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(VCC_net), .O(n2456[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(GND_net), 
            .CO(n38848));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2522), .I1(n2489), .I2(VCC_net), 
            .I3(n38847), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(GND_net), .I1(n2490), .I2(VCC_net), 
            .I3(n38846), .O(n2555[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_22 (.CI(n38846), .I0(n2490), .I1(VCC_net), 
            .CO(n38847));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(GND_net), .I1(n2491), .I2(VCC_net), 
            .I3(n38845), .O(n2555[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_21 (.CI(n38845), .I0(n2491), .I1(VCC_net), 
            .CO(n38846));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(GND_net), .I1(n2492), .I2(VCC_net), 
            .I3(n38844), .O(n2555[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_20 (.CI(n38844), .I0(n2492), .I1(VCC_net), 
            .CO(n38845));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(GND_net), .I1(n2493), .I2(VCC_net), 
            .I3(n38843), .O(n2555[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_19 (.CI(n38843), .I0(n2493), .I1(VCC_net), 
            .CO(n38844));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(GND_net), .I1(n2494), .I2(VCC_net), 
            .I3(n38842), .O(n2555[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_18 (.CI(n38842), .I0(n2494), .I1(VCC_net), 
            .CO(n38843));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(GND_net), .I1(n2495), .I2(VCC_net), 
            .I3(n38841), .O(n2555[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_17 (.CI(n38841), .I0(n2495), .I1(VCC_net), 
            .CO(n38842));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(GND_net), .I1(n2496), .I2(VCC_net), 
            .I3(n38840), .O(n2555[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_16 (.CI(n38840), .I0(n2496), .I1(VCC_net), 
            .CO(n38841));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(GND_net), .I1(n2497), .I2(VCC_net), 
            .I3(n38839), .O(n2555[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_15 (.CI(n38839), .I0(n2497), .I1(VCC_net), 
            .CO(n38840));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(GND_net), .I1(n2498), .I2(VCC_net), 
            .I3(n38838), .O(n2555[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_14 (.CI(n38838), .I0(n2498), .I1(VCC_net), 
            .CO(n38839));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(GND_net), .I1(n2499), .I2(VCC_net), 
            .I3(n38837), .O(n2555[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_13 (.CI(n38837), .I0(n2499), .I1(VCC_net), 
            .CO(n38838));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(GND_net), .I1(n2500), .I2(VCC_net), 
            .I3(n38836), .O(n2555[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_12 (.CI(n38836), .I0(n2500), .I1(VCC_net), 
            .CO(n38837));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(GND_net), .I1(n2501), .I2(VCC_net), 
            .I3(n38835), .O(n2555[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_11 (.CI(n38835), .I0(n2501), .I1(VCC_net), 
            .CO(n38836));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(GND_net), .I1(n2502), .I2(VCC_net), 
            .I3(n38834), .O(n2555[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_10 (.CI(n38834), .I0(n2502), .I1(VCC_net), 
            .CO(n38835));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(GND_net), .I1(n2503), .I2(VCC_net), 
            .I3(n38833), .O(n2555[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n37360), .I0(timer[11]), .I1(n1[11]), 
            .CO(n37361));
    SB_CARRY mod_5_add_1741_9 (.CI(n38833), .I0(n2503), .I1(VCC_net), 
            .CO(n38834));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(GND_net), .I1(n2504), .I2(VCC_net), 
            .I3(n38832), .O(n2555[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_8 (.CI(n38832), .I0(n2504), .I1(VCC_net), 
            .CO(n38833));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(GND_net), .I1(n2505), .I2(VCC_net), 
            .I3(n38831), .O(n2555[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_7 (.CI(n38831), .I0(n2505), .I1(VCC_net), 
            .CO(n38832));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(GND_net), .I1(n2506), .I2(VCC_net), 
            .I3(n38830), .O(n2555[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_6 (.CI(n38830), .I0(n2506), .I1(VCC_net), 
            .CO(n38831));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(GND_net), .I1(n2507), .I2(VCC_net), 
            .I3(n38829), .O(n2555[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_5 (.CI(n38829), .I0(n2507), .I1(VCC_net), 
            .CO(n38830));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n37359), .O(one_wire_N_579[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(GND_net), .I1(n2508), .I2(VCC_net), 
            .I3(n38828), .O(n2555[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_4 (.CI(n38828), .I0(n2508), .I1(VCC_net), 
            .CO(n38829));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(GND_net), .I1(n2509), .I2(GND_net), 
            .I3(n38827), .O(n2555[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_3 (.CI(n38827), .I0(n2509), .I1(GND_net), 
            .CO(n38828));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(VCC_net), .O(n2555[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(GND_net), 
            .CO(n38827));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2621), .I1(n2588), .I2(VCC_net), 
            .I3(n38826), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_12 (.CI(n37359), .I0(timer[10]), .I1(n1[10]), 
            .CO(n37360));
    SB_LUT4 mod_5_add_1808_23_lut (.I0(GND_net), .I1(n2589), .I2(VCC_net), 
            .I3(n38825), .O(n2654[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_23 (.CI(n38825), .I0(n2589), .I1(VCC_net), 
            .CO(n38826));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(GND_net), .I1(n2590), .I2(VCC_net), 
            .I3(n38824), .O(n2654[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_22 (.CI(n38824), .I0(n2590), .I1(VCC_net), 
            .CO(n38825));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n37358), .O(one_wire_N_579[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_21_lut (.I0(GND_net), .I1(n2591), .I2(VCC_net), 
            .I3(n38823), .O(n2654[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n37226), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_21 (.CI(n38823), .I0(n2591), .I1(VCC_net), 
            .CO(n38824));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(GND_net), .I1(n2592), .I2(VCC_net), 
            .I3(n38822), .O(n2654[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_20 (.CI(n38822), .I0(n2592), .I1(VCC_net), 
            .CO(n38823));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(GND_net), .I1(n2593), .I2(VCC_net), 
            .I3(n38821), .O(n2654[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_0__bdd_4_lut_34520 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n49347));
    defparam bit_ctr_0__bdd_4_lut_34520.LUT_INIT = 16'he4aa;
    SB_LUT4 n49347_bdd_4_lut (.I0(n49347), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n49350));
    defparam n49347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_34377 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n49341));
    defparam bit_ctr_0__bdd_4_lut_34377.LUT_INIT = 16'he4aa;
    SB_LUT4 n49341_bdd_4_lut (.I0(n49341), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n49344));
    defparam n49341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY mod_5_add_1808_19 (.CI(n38821), .I0(n2593), .I1(VCC_net), 
            .CO(n38822));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(GND_net), .I1(n2594), .I2(VCC_net), 
            .I3(n38820), .O(n2654[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_18 (.CI(n38820), .I0(n2594), .I1(VCC_net), 
            .CO(n38821));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(GND_net), .I1(n2595), .I2(VCC_net), 
            .I3(n38819), .O(n2654[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_17 (.CI(n38819), .I0(n2595), .I1(VCC_net), 
            .CO(n38820));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(GND_net), .I1(n2596), .I2(VCC_net), 
            .I3(n38818), .O(n2654[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n37358), .I0(timer[9]), .I1(n1[9]), 
            .CO(n37359));
    SB_CARRY add_21_14 (.CI(n37226), .I0(bit_ctr[12]), .I1(GND_net), .CO(n37227));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n37357), .O(one_wire_N_579[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_16 (.CI(n38818), .I0(n2596), .I1(VCC_net), 
            .CO(n38819));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(GND_net), .I1(n2597), .I2(VCC_net), 
            .I3(n38817), .O(n2654[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_15 (.CI(n38817), .I0(n2597), .I1(VCC_net), 
            .CO(n38818));
    SB_CARRY sub_14_add_2_10 (.CI(n37357), .I0(timer[8]), .I1(n1[8]), 
            .CO(n37358));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(GND_net), .I1(n2598), .I2(VCC_net), 
            .I3(n38816), .O(n2654[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_14 (.CI(n38816), .I0(n2598), .I1(VCC_net), 
            .CO(n38817));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n37225), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_9_lut (.I0(n46350), .I1(timer[7]), .I2(n1[7]), 
            .I3(n37356), .O(n46352)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_9 (.CI(n37356), .I0(timer[7]), .I1(n1[7]), .CO(n37357));
    SB_LUT4 sub_14_add_2_8_lut (.I0(n46348), .I1(timer[6]), .I2(n1[6]), 
            .I3(n37355), .O(n46350)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_8 (.CI(n37355), .I0(timer[6]), .I1(n1[6]), .CO(n37356));
    SB_LUT4 sub_14_add_2_7_lut (.I0(one_wire_N_579[4]), .I1(timer[5]), .I2(n1[5]), 
            .I3(n37354), .O(n46348)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1808_13_lut (.I0(GND_net), .I1(n2599), .I2(VCC_net), 
            .I3(n38815), .O(n2654[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_13 (.CI(n38815), .I0(n2599), .I1(VCC_net), 
            .CO(n38816));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(GND_net), .I1(n2600), .I2(VCC_net), 
            .I3(n38814), .O(n2654[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n37354), .I0(timer[5]), .I1(n1[5]), .CO(n37355));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n37353), .O(one_wire_N_579[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n37353), .I0(timer[4]), .I1(n1[4]), .CO(n37354));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n37352), .O(one_wire_N_579[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n37352), .I0(timer[3]), .I1(n1[3]), .CO(n37353));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n37351), .O(one_wire_N_579[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_13 (.CI(n37225), .I0(bit_ctr[11]), .I1(GND_net), .CO(n37226));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n37224), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_12 (.CI(n38814), .I0(n2600), .I1(VCC_net), 
            .CO(n38815));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(GND_net), .I1(n2601), .I2(VCC_net), 
            .I3(n38813), .O(n2654[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_11 (.CI(n38813), .I0(n2601), .I1(VCC_net), 
            .CO(n38814));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(GND_net), .I1(n2602), .I2(VCC_net), 
            .I3(n38812), .O(n2654[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_10 (.CI(n38812), .I0(n2602), .I1(VCC_net), 
            .CO(n38813));
    SB_CARRY add_21_12 (.CI(n37224), .I0(bit_ctr[10]), .I1(GND_net), .CO(n37225));
    SB_CARRY sub_14_add_2_4 (.CI(n37351), .I0(timer[2]), .I1(n1[2]), .CO(n37352));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n37223), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_9_lut (.I0(GND_net), .I1(n2603), .I2(VCC_net), 
            .I3(n38811), .O(n2654[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_9 (.CI(n38811), .I0(n2603), .I1(VCC_net), 
            .CO(n38812));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(GND_net), .I1(n2604), .I2(VCC_net), 
            .I3(n38810), .O(n2654[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_8 (.CI(n38810), .I0(n2604), .I1(VCC_net), 
            .CO(n38811));
    SB_CARRY add_21_11 (.CI(n37223), .I0(bit_ctr[9]), .I1(GND_net), .CO(n37224));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(GND_net), .I1(n2605), .I2(VCC_net), 
            .I3(n38809), .O(n2654[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_7 (.CI(n38809), .I0(n2605), .I1(VCC_net), 
            .CO(n38810));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(GND_net), .I1(n2606), .I2(VCC_net), 
            .I3(n38808), .O(n2654[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_579[2]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n37350), .O(n4_adj_4893)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1808_6 (.CI(n38808), .I0(n2606), .I1(VCC_net), 
            .CO(n38809));
    SB_CARRY sub_14_add_2_3 (.CI(n37350), .I0(timer[1]), .I1(n1[1]), .CO(n37351));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(GND_net), .I1(n2607), .I2(VCC_net), 
            .I3(n38807), .O(n2654[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_5 (.CI(n38807), .I0(n2607), .I1(VCC_net), 
            .CO(n38808));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n37350));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(GND_net), .I1(n2608), .I2(VCC_net), 
            .I3(n38806), .O(n2654[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n37222), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_4 (.CI(n38806), .I0(n2608), .I1(VCC_net), 
            .CO(n38807));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(GND_net), .I1(n2609), .I2(GND_net), 
            .I3(n38805), .O(n2654[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_3 (.CI(n38805), .I0(n2609), .I1(GND_net), 
            .CO(n38806));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(VCC_net), .O(n2654[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(GND_net), 
            .CO(n38805));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2720), .I1(n2687), .I2(VCC_net), 
            .I3(n38804), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(GND_net), .I1(n2688), .I2(VCC_net), 
            .I3(n38803), .O(n2753[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_24 (.CI(n38803), .I0(n2688), .I1(VCC_net), 
            .CO(n38804));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(GND_net), .I1(n2689), .I2(VCC_net), 
            .I3(n38802), .O(n2753[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_23 (.CI(n38802), .I0(n2689), .I1(VCC_net), 
            .CO(n38803));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(GND_net), .I1(n2690), .I2(VCC_net), 
            .I3(n38801), .O(n2753[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_22 (.CI(n38801), .I0(n2690), .I1(VCC_net), 
            .CO(n38802));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(GND_net), .I1(n2691), .I2(VCC_net), 
            .I3(n38800), .O(n2753[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1532), .I1(n1499), .I2(VCC_net), 
            .I3(n37609), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(GND_net), .I1(n1500), .I2(VCC_net), 
            .I3(n37608), .O(n1565[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_21 (.CI(n38800), .I0(n2691), .I1(VCC_net), 
            .CO(n38801));
    SB_CARRY mod_5_add_1071_12 (.CI(n37608), .I0(n1500), .I1(VCC_net), 
            .CO(n37609));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(GND_net), .I1(n1501), .I2(VCC_net), 
            .I3(n37607), .O(n1565[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_11 (.CI(n37607), .I0(n1501), .I1(VCC_net), 
            .CO(n37608));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(GND_net), .I1(n2692), .I2(VCC_net), 
            .I3(n38799), .O(n2753[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_20 (.CI(n38799), .I0(n2692), .I1(VCC_net), 
            .CO(n38800));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(GND_net), .I1(n2693), .I2(VCC_net), 
            .I3(n38798), .O(n2753[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_19 (.CI(n38798), .I0(n2693), .I1(VCC_net), 
            .CO(n38799));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(GND_net), .I1(n1502), .I2(VCC_net), 
            .I3(n37606), .O(n1565[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_18_lut (.I0(GND_net), .I1(n2694), .I2(VCC_net), 
            .I3(n38797), .O(n2753[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_10 (.CI(n37606), .I0(n1502), .I1(VCC_net), 
            .CO(n37607));
    SB_CARRY mod_5_add_1875_18 (.CI(n38797), .I0(n2694), .I1(VCC_net), 
            .CO(n38798));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(GND_net), .I1(n1503), .I2(VCC_net), 
            .I3(n37605), .O(n1565[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_9 (.CI(n37605), .I0(n1503), .I1(VCC_net), 
            .CO(n37606));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(GND_net), .I1(n2695), .I2(VCC_net), 
            .I3(n38796), .O(n2753[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_8_lut (.I0(GND_net), .I1(n1504), .I2(VCC_net), 
            .I3(n37604), .O(n1565[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_8 (.CI(n37604), .I0(n1504), .I1(VCC_net), 
            .CO(n37605));
    SB_CARRY mod_5_add_1875_17 (.CI(n38796), .I0(n2695), .I1(VCC_net), 
            .CO(n38797));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(GND_net), .I1(n2696), .I2(VCC_net), 
            .I3(n38795), .O(n2753[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_10 (.CI(n37222), .I0(bit_ctr[8]), .I1(GND_net), .CO(n37223));
    SB_CARRY mod_5_add_1875_16 (.CI(n38795), .I0(n2696), .I1(VCC_net), 
            .CO(n38796));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n37221), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_15_lut (.I0(GND_net), .I1(n2697), .I2(VCC_net), 
            .I3(n38794), .O(n2753[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_15 (.CI(n38794), .I0(n2697), .I1(VCC_net), 
            .CO(n38795));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(GND_net), .I1(n2698), .I2(VCC_net), 
            .I3(n38793), .O(n2753[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_14 (.CI(n38793), .I0(n2698), .I1(VCC_net), 
            .CO(n38794));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(GND_net), .I1(n2699), .I2(VCC_net), 
            .I3(n38792), .O(n2753[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_13 (.CI(n38792), .I0(n2699), .I1(VCC_net), 
            .CO(n38793));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(GND_net), .I1(n2700), .I2(VCC_net), 
            .I3(n38791), .O(n2753[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_12 (.CI(n38791), .I0(n2700), .I1(VCC_net), 
            .CO(n38792));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(GND_net), .I1(n1505), .I2(VCC_net), 
            .I3(n37603), .O(n1565[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_7 (.CI(n37603), .I0(n1505), .I1(VCC_net), 
            .CO(n37604));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(GND_net), .I1(n1506), .I2(VCC_net), 
            .I3(n37602), .O(n1565[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_6 (.CI(n37602), .I0(n1506), .I1(VCC_net), 
            .CO(n37603));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(GND_net), .I1(n1507), .I2(VCC_net), 
            .I3(n37601), .O(n1565[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_11_lut (.I0(GND_net), .I1(n2701), .I2(VCC_net), 
            .I3(n38790), .O(n2753[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_9 (.CI(n37221), .I0(bit_ctr[7]), .I1(GND_net), .CO(n37222));
    SB_CARRY mod_5_add_1071_5 (.CI(n37601), .I0(n1507), .I1(VCC_net), 
            .CO(n37602));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(GND_net), .I1(n1508), .I2(VCC_net), 
            .I3(n37600), .O(n1565[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_4 (.CI(n37600), .I0(n1508), .I1(VCC_net), 
            .CO(n37601));
    SB_CARRY mod_5_add_1875_11 (.CI(n38790), .I0(n2701), .I1(VCC_net), 
            .CO(n38791));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(GND_net), .I1(n2702), .I2(VCC_net), 
            .I3(n38789), .O(n2753[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_10 (.CI(n38789), .I0(n2702), .I1(VCC_net), 
            .CO(n38790));
    SB_LUT4 mod_5_i1488_3_lut (.I0(n2106), .I1(n2159[18]), .I2(n2126), 
            .I3(GND_net), .O(n2205));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1479_3_lut (.I0(n2097), .I1(n2159[27]), .I2(n2126), 
            .I3(GND_net), .O(n2196));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1482_3_lut (.I0(n2100), .I1(n2159[24]), .I2(n2126), 
            .I3(GND_net), .O(n2199));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1491_3_lut (.I0(n2109), .I1(n2159[15]), .I2(n2126), 
            .I3(GND_net), .O(n2208));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1484_3_lut (.I0(n2102), .I1(n2159[22]), .I2(n2126), 
            .I3(GND_net), .O(n2201));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1486_3_lut (.I0(n2104), .I1(n2159[20]), .I2(n2126), 
            .I3(GND_net), .O(n2203));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1485_3_lut (.I0(n2103), .I1(n2159[21]), .I2(n2126), 
            .I3(GND_net), .O(n2202));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1483_3_lut (.I0(n2101), .I1(n2159[23]), .I2(n2126), 
            .I3(GND_net), .O(n2200));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1489_3_lut (.I0(n2107), .I1(n2159[17]), .I2(n2126), 
            .I3(GND_net), .O(n2206));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1490_3_lut (.I0(n2108), .I1(n2159[16]), .I2(n2126), 
            .I3(GND_net), .O(n2207));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1071_3_lut (.I0(GND_net), .I1(n1509), .I2(GND_net), 
            .I3(n37599), .O(n1565[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_3 (.CI(n37599), .I0(n1509), .I1(GND_net), 
            .CO(n37600));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(VCC_net), .O(n1565[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(GND_net), 
            .CO(n37599));
    SB_LUT4 mod_5_i1481_3_lut (.I0(n2099), .I1(n2159[25]), .I2(n2126), 
            .I3(GND_net), .O(n2198));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(GND_net), .I1(n2703), .I2(VCC_net), 
            .I3(n38788), .O(n2753[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n37220), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_9 (.CI(n38788), .I0(n2703), .I1(VCC_net), 
            .CO(n38789));
    SB_LUT4 mod_5_i1487_3_lut (.I0(n2105), .I1(n2159[19]), .I2(n2126), 
            .I3(GND_net), .O(n2204));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1492_3_lut (.I0(bit_ctr[14]), .I1(n2159[14]), .I2(n2126), 
            .I3(GND_net), .O(n2209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_8_lut (.I0(GND_net), .I1(n2704), .I2(VCC_net), 
            .I3(n38787), .O(n2753[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_8 (.CI(n38787), .I0(n2704), .I1(VCC_net), 
            .CO(n38788));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(GND_net), .I1(n2705), .I2(VCC_net), 
            .I3(n38786), .O(n2753[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_7 (.CI(n38786), .I0(n2705), .I1(VCC_net), 
            .CO(n38787));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(GND_net), .I1(n2706), .I2(VCC_net), 
            .I3(n38785), .O(n2753[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1480_3_lut (.I0(n2098), .I1(n2159[26]), .I2(n2126), 
            .I3(GND_net), .O(n2197));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1478_3_lut (.I0(n2096), .I1(n2159[28]), .I2(n2126), 
            .I3(GND_net), .O(n2195));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1478_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_8 (.CI(n37220), .I0(bit_ctr[6]), .I1(GND_net), .CO(n37221));
    SB_CARRY mod_5_add_1875_6 (.CI(n38785), .I0(n2706), .I1(VCC_net), 
            .CO(n38786));
    SB_LUT4 mod_5_i1477_3_lut (.I0(n2095), .I1(n2159[29]), .I2(n2126), 
            .I3(GND_net), .O(n2194));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1476_3_lut (.I0(n2094), .I1(n2159[30]), .I2(n2126), 
            .I3(GND_net), .O(n2193));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_5_lut (.I0(GND_net), .I1(n2707), .I2(VCC_net), 
            .I3(n38784), .O(n2753[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_5 (.CI(n38784), .I0(n2707), .I1(VCC_net), 
            .CO(n38785));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(GND_net), .I1(n2708), .I2(VCC_net), 
            .I3(n38783), .O(n2753[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_4 (.CI(n38783), .I0(n2708), .I1(VCC_net), 
            .CO(n38784));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(GND_net), .I1(n2709), .I2(GND_net), 
            .I3(n38782), .O(n2753[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_3 (.CI(n38782), .I0(n2709), .I1(GND_net), 
            .CO(n38783));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(VCC_net), .O(n2753[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(GND_net), 
            .CO(n38782));
    SB_LUT4 i10_4_lut (.I0(n2193), .I1(n2194), .I2(n2192), .I3(n2195), 
            .O(n28_adj_4899));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1616 (.I0(n2204), .I1(n2198), .I2(n2207), .I3(n2206), 
            .O(n31_adj_4900));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1617 (.I0(bit_ctr[13]), .I1(n2197), .I2(n2209), 
            .I3(GND_net), .O(n22_adj_4901));   // verilog/neopixel.v(22[26:36])
    defparam i4_3_lut_adj_1617.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n38781), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_4_lut_adj_1618 (.I0(n2200), .I1(n2202), .I2(n2203), .I3(n2201), 
            .O(n30_adj_4902));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1619 (.I0(n31_adj_4900), .I1(n2208), .I2(n28_adj_4899), 
            .I3(n2199), .O(n34_adj_4903));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut (.I0(n2196), .I1(n2205), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_4904));   // verilog/neopixel.v(22[26:36])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(CLK_c), .E(n27897), .D(state_3__N_428[0]), 
            .S(n28098));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n38780), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n38780), .I0(n2787), .I1(n2819), .CO(n38781));
    SB_LUT4 i17_4_lut_adj_1620 (.I0(n21_adj_4904), .I1(n34_adj_4903), .I2(n30_adj_4902), 
            .I3(n22_adj_4901), .O(n2225));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n38779), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n38779), .I0(n2788), .I1(n2819), .CO(n38780));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n38778), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n38778), .I0(n2789), .I1(n2819), .CO(n38779));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n38777), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n38777), .I0(n2790), .I1(n2819), .CO(n38778));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n38776), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n38776), .I0(n2791), .I1(n2819), .CO(n38777));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n38775), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n38775), .I0(n2792), .I1(n2819), .CO(n38776));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n38774), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n38774), .I0(n2793), .I1(n2819), .CO(n38775));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n38773), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n38773), .I0(n2794), .I1(n2819), .CO(n38774));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n38772), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n38772), .I0(n2795), .I1(n2819), .CO(n38773));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n38771), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n38771), .I0(n2796), .I1(n2819), .CO(n38772));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n38770), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n38770), .I0(n2797), .I1(n2819), .CO(n38771));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n38769), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n38769), .I0(n2798), .I1(n2819), .CO(n38770));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n38768), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n38768), .I0(n2799), .I1(n2819), .CO(n38769));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n38767), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n38767), .I0(n2800), .I1(n2819), .CO(n38768));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n38766), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n38766), .I0(n2801), .I1(n2819), .CO(n38767));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n38765), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n38765), .I0(n2802), .I1(n2819), .CO(n38766));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n38764), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n38764), .I0(n2803), .I1(n2819), .CO(n38765));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n38763), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n38763), .I0(n2804), .I1(n2819), .CO(n38764));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n38762), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n38762), .I0(n2805), .I1(n2819), .CO(n38763));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n38761), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n37219), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_6 (.CI(n38761), .I0(n2806), .I1(n2819), .CO(n38762));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n38760), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n38760), .I0(n2807), .I1(n2819), .CO(n38761));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n38759), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n38759), .I0(n2808), .I1(n2819), .CO(n38760));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n49246), 
            .I3(n38758), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n38758), .I0(n2809), .I1(n49246), .CO(n38759));
    SB_CARRY add_21_7 (.CI(n37219), .I0(bit_ctr[5]), .I1(GND_net), .CO(n37220));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n49246), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n49246), 
            .CO(n38758));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n37218), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2918), .I1(n2885), .I2(VCC_net), 
            .I3(n38757), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(GND_net), .I1(n2886), .I2(VCC_net), 
            .I3(n38756), .O(n2951[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_26 (.CI(n38756), .I0(n2886), .I1(VCC_net), 
            .CO(n38757));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(GND_net), .I1(n2887), .I2(VCC_net), 
            .I3(n38755), .O(n2951[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_25 (.CI(n38755), .I0(n2887), .I1(VCC_net), 
            .CO(n38756));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(GND_net), .I1(n2888), .I2(VCC_net), 
            .I3(n38754), .O(n2951[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_24 (.CI(n38754), .I0(n2888), .I1(VCC_net), 
            .CO(n38755));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(GND_net), .I1(n2889), .I2(VCC_net), 
            .I3(n38753), .O(n2951[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_23 (.CI(n38753), .I0(n2889), .I1(VCC_net), 
            .CO(n38754));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(GND_net), .I1(n2890), .I2(VCC_net), 
            .I3(n38752), .O(n2951[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_22 (.CI(n38752), .I0(n2890), .I1(VCC_net), 
            .CO(n38753));
    SB_CARRY add_21_6 (.CI(n37218), .I0(bit_ctr[4]), .I1(GND_net), .CO(n37219));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(GND_net), .I1(n2891), .I2(VCC_net), 
            .I3(n38751), .O(n2951[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_21 (.CI(n38751), .I0(n2891), .I1(VCC_net), 
            .CO(n38752));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(GND_net), .I1(n2892), .I2(VCC_net), 
            .I3(n38750), .O(n2951[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_20 (.CI(n38750), .I0(n2892), .I1(VCC_net), 
            .CO(n38751));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(GND_net), .I1(n2893), .I2(VCC_net), 
            .I3(n38749), .O(n2951[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_19 (.CI(n38749), .I0(n2893), .I1(VCC_net), 
            .CO(n38750));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(GND_net), .I1(n2894), .I2(VCC_net), 
            .I3(n38748), .O(n2951[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_18 (.CI(n38748), .I0(n2894), .I1(VCC_net), 
            .CO(n38749));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(GND_net), .I1(n2895), .I2(VCC_net), 
            .I3(n38747), .O(n2951[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_17 (.CI(n38747), .I0(n2895), .I1(VCC_net), 
            .CO(n38748));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(GND_net), .I1(n2896), .I2(VCC_net), 
            .I3(n38746), .O(n2951[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_16 (.CI(n38746), .I0(n2896), .I1(VCC_net), 
            .CO(n38747));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(GND_net), .I1(n2897), .I2(VCC_net), 
            .I3(n38745), .O(n2951[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n37217), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_15 (.CI(n38745), .I0(n2897), .I1(VCC_net), 
            .CO(n38746));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(GND_net), .I1(n2898), .I2(VCC_net), 
            .I3(n38744), .O(n2951[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_14 (.CI(n38744), .I0(n2898), .I1(VCC_net), 
            .CO(n38745));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(GND_net), .I1(n2899), .I2(VCC_net), 
            .I3(n38743), .O(n2951[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_13 (.CI(n38743), .I0(n2899), .I1(VCC_net), 
            .CO(n38744));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(GND_net), .I1(n2900), .I2(VCC_net), 
            .I3(n38742), .O(n2951[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n38742), .I0(n2900), .I1(VCC_net), 
            .CO(n38743));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(GND_net), .I1(n2901), .I2(VCC_net), 
            .I3(n38741), .O(n2951[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_11 (.CI(n38741), .I0(n2901), .I1(VCC_net), 
            .CO(n38742));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(GND_net), .I1(n2902), .I2(VCC_net), 
            .I3(n38740), .O(n2951[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_10 (.CI(n38740), .I0(n2902), .I1(VCC_net), 
            .CO(n38741));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(GND_net), .I1(n2903), .I2(VCC_net), 
            .I3(n38739), .O(n2951[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_9 (.CI(n38739), .I0(n2903), .I1(VCC_net), 
            .CO(n38740));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(GND_net), .I1(n2904), .I2(VCC_net), 
            .I3(n38738), .O(n2951[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_8 (.CI(n38738), .I0(n2904), .I1(VCC_net), 
            .CO(n38739));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(GND_net), .I1(n2905), .I2(VCC_net), 
            .I3(n38737), .O(n2951[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_7 (.CI(n38737), .I0(n2905), .I1(VCC_net), 
            .CO(n38738));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(GND_net), .I1(n2906), .I2(VCC_net), 
            .I3(n38736), .O(n2951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_6 (.CI(n38736), .I0(n2906), .I1(VCC_net), 
            .CO(n38737));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(GND_net), .I1(n2907), .I2(VCC_net), 
            .I3(n38735), .O(n2951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_5 (.CI(n38735), .I0(n2907), .I1(VCC_net), 
            .CO(n38736));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(GND_net), .I1(n2908), .I2(VCC_net), 
            .I3(n38734), .O(n2951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n38734), .I0(n2908), .I1(VCC_net), 
            .CO(n38735));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(GND_net), .I1(n2909), .I2(GND_net), 
            .I3(n38733), .O(n2951[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_3 (.CI(n38733), .I0(n2909), .I1(GND_net), 
            .CO(n38734));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(VCC_net), .O(n2951[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(GND_net), 
            .CO(n38733));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n38732), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n38731), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n38731), .I0(n2985), .I1(n3017), .CO(n38732));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n38730), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n38730), .I0(n2986), .I1(n3017), .CO(n38731));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n38729), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n38729), .I0(n2987), .I1(n3017), .CO(n38730));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n38728), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n38728), .I0(n2988), .I1(n3017), .CO(n38729));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n38727), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n38727), .I0(n2989), .I1(n3017), .CO(n38728));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n38726), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n38726), .I0(n2990), .I1(n3017), .CO(n38727));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n38725), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n38725), .I0(n2991), .I1(n3017), .CO(n38726));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n38724), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n38724), .I0(n2992), .I1(n3017), .CO(n38725));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n38723), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n38723), .I0(n2993), .I1(n3017), .CO(n38724));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n38722), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n38722), .I0(n2994), .I1(n3017), .CO(n38723));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n38721), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n38721), .I0(n2995), .I1(n3017), .CO(n38722));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n38720), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n38720), .I0(n2996), .I1(n3017), .CO(n38721));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n38719), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n38719), .I0(n2997), .I1(n3017), .CO(n38720));
    SB_CARRY add_21_5 (.CI(n37217), .I0(bit_ctr[3]), .I1(GND_net), .CO(n37218));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n38718), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n38718), .I0(n2998), .I1(n3017), .CO(n38719));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n38717), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n38717), .I0(n2999), .I1(n3017), .CO(n38718));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n38716), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n38716), .I0(n3000), .I1(n3017), .CO(n38717));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n38715), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n38715), .I0(n3001), .I1(n3017), .CO(n38716));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n38714), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n38714), .I0(n3002), .I1(n3017), .CO(n38715));
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n37216), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n38713), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n38713), .I0(n3003), .I1(n3017), .CO(n38714));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n38712), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n38712), .I0(n3004), .I1(n3017), .CO(n38713));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n38711), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n38711), .I0(n3005), .I1(n3017), .CO(n38712));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n38710), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n38710), .I0(n3006), .I1(n3017), .CO(n38711));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n38709), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n38709), .I0(n3007), .I1(n3017), .CO(n38710));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n38708), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n38708), .I0(n3008), .I1(n3017), .CO(n38709));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n30674), .I1(n30674), .I2(n49247), 
            .I3(n38707), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n38707), .I0(n30674), .I1(n49247), 
            .CO(n38708));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n49247), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n49247), 
            .CO(n38707));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3116), .I1(n3083), .I2(VCC_net), 
            .I3(n38706), .O(n46490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(GND_net), .I1(n3084), .I2(VCC_net), 
            .I3(n38705), .O(n3149[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_28 (.CI(n38705), .I0(n3084), .I1(VCC_net), 
            .CO(n38706));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(GND_net), .I1(n3085), .I2(VCC_net), 
            .I3(n38704), .O(n3149[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_27 (.CI(n38704), .I0(n3085), .I1(VCC_net), 
            .CO(n38705));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(GND_net), .I1(n3086), .I2(VCC_net), 
            .I3(n38703), .O(n3149[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_26 (.CI(n38703), .I0(n3086), .I1(VCC_net), 
            .CO(n38704));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(GND_net), .I1(n3087), .I2(VCC_net), 
            .I3(n38702), .O(n3149[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_25 (.CI(n38702), .I0(n3087), .I1(VCC_net), 
            .CO(n38703));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(GND_net), .I1(n3088), .I2(VCC_net), 
            .I3(n38701), .O(n3149[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_24 (.CI(n38701), .I0(n3088), .I1(VCC_net), 
            .CO(n38702));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(GND_net), .I1(n3089), .I2(VCC_net), 
            .I3(n38700), .O(n3149[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_23 (.CI(n38700), .I0(n3089), .I1(VCC_net), 
            .CO(n38701));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(GND_net), .I1(n3090), .I2(VCC_net), 
            .I3(n38699), .O(n3149[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_22 (.CI(n38699), .I0(n3090), .I1(VCC_net), 
            .CO(n38700));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(GND_net), .I1(n3091), .I2(VCC_net), 
            .I3(n38698), .O(n3149[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_21 (.CI(n38698), .I0(n3091), .I1(VCC_net), 
            .CO(n38699));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(GND_net), .I1(n3092), .I2(VCC_net), 
            .I3(n38697), .O(n3149[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_20 (.CI(n38697), .I0(n3092), .I1(VCC_net), 
            .CO(n38698));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(GND_net), .I1(n3093), .I2(VCC_net), 
            .I3(n38696), .O(n3149[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_19 (.CI(n38696), .I0(n3093), .I1(VCC_net), 
            .CO(n38697));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(GND_net), .I1(n3094), .I2(VCC_net), 
            .I3(n38695), .O(n3149[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_18 (.CI(n38695), .I0(n3094), .I1(VCC_net), 
            .CO(n38696));
    SB_CARRY add_21_4 (.CI(n37216), .I0(bit_ctr[2]), .I1(GND_net), .CO(n37217));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(GND_net), .I1(n3095), .I2(VCC_net), 
            .I3(n38694), .O(n3149[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_17 (.CI(n38694), .I0(n3095), .I1(VCC_net), 
            .CO(n38695));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(GND_net), .I1(n3096), .I2(VCC_net), 
            .I3(n38693), .O(n3149[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_16 (.CI(n38693), .I0(n3096), .I1(VCC_net), 
            .CO(n38694));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(GND_net), .I1(n3097), .I2(VCC_net), 
            .I3(n38692), .O(n3149[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_15 (.CI(n38692), .I0(n3097), .I1(VCC_net), 
            .CO(n38693));
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n37215), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_14_lut (.I0(GND_net), .I1(n3098), .I2(VCC_net), 
            .I3(n38691), .O(n3149[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_14 (.CI(n38691), .I0(n3098), .I1(VCC_net), 
            .CO(n38692));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(GND_net), .I1(n3099), .I2(VCC_net), 
            .I3(n38690), .O(n3149[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_13 (.CI(n38690), .I0(n3099), .I1(VCC_net), 
            .CO(n38691));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(GND_net), .I1(n3100), .I2(VCC_net), 
            .I3(n38689), .O(n3149[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_12 (.CI(n38689), .I0(n3100), .I1(VCC_net), 
            .CO(n38690));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(GND_net), .I1(n3101), .I2(VCC_net), 
            .I3(n38688), .O(n3149[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_11 (.CI(n38688), .I0(n3101), .I1(VCC_net), 
            .CO(n38689));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(GND_net), .I1(n3102), .I2(VCC_net), 
            .I3(n38687), .O(n3149[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_10 (.CI(n38687), .I0(n3102), .I1(VCC_net), 
            .CO(n38688));
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n27723), .D(n255[0]), 
            .R(n28057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1547__i1 (.Q(timer[1]), .C(CLK_c), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_2143_9_lut (.I0(GND_net), .I1(n3103), .I2(VCC_net), 
            .I3(n38686), .O(n3149[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_9 (.CI(n38686), .I0(n3103), .I1(VCC_net), 
            .CO(n38687));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(GND_net), .I1(n3104), .I2(VCC_net), 
            .I3(n38685), .O(n3149[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_8 (.CI(n38685), .I0(n3104), .I1(VCC_net), 
            .CO(n38686));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(GND_net), .I1(n3105), .I2(VCC_net), 
            .I3(n38684), .O(n3149[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_7 (.CI(n38684), .I0(n3105), .I1(VCC_net), 
            .CO(n38685));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(GND_net), .I1(n3106), .I2(VCC_net), 
            .I3(n38683), .O(n3149[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_6 (.CI(n38683), .I0(n3106), .I1(VCC_net), 
            .CO(n38684));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(GND_net), .I1(n3107), .I2(VCC_net), 
            .I3(n38682), .O(n3149[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_5 (.CI(n38682), .I0(n3107), .I1(VCC_net), 
            .CO(n38683));
    SB_CARRY add_21_3 (.CI(n37215), .I0(bit_ctr[1]), .I1(GND_net), .CO(n37216));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(GND_net), .I1(n3108), .I2(VCC_net), 
            .I3(n38681), .O(n3149[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_4 (.CI(n38681), .I0(n3108), .I1(VCC_net), 
            .CO(n38682));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(GND_net), .I1(n3109), .I2(GND_net), 
            .I3(n38680), .O(n3149[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_3 (.CI(n38680), .I0(n3109), .I1(GND_net), 
            .CO(n38681));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(VCC_net), .O(n3149[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(GND_net), 
            .CO(n38680));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n37215));
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n37334), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n37333), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n37333), .I0(GND_net), .I1(VCC_net), 
            .CO(n37334));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n27993), .I2(VCC_net), 
            .I3(n37332), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n37332), .I0(n27993), .I1(VCC_net), 
            .CO(n37333));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n27950), .I2(VCC_net), 
            .I3(n37331), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n37331), .I0(n27950), .I1(VCC_net), 
            .CO(n37332));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n25171), .I2(GND_net), 
            .I3(n37330), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n37330), .I0(n25171), .I1(GND_net), 
            .CO(n37331));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n37330));
    SB_LUT4 i1_2_lut_3_lut_adj_1621 (.I0(bit_ctr[27]), .I1(n25173), .I2(n27956), 
            .I3(GND_net), .O(n25171));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_adj_1621.LUT_INIT = 16'h8585;
    SB_DFFE start_103 (.Q(start), .C(CLK_c), .E(VCC_net), .D(n41189));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n48267), .D(\neo_pixel_transmitter.done_N_642 ), 
            .R(n44951));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i21466_4_lut (.I0(one_wire_N_579[10]), .I1(n160), .I2(one_wire_N_579[8]), 
            .I3(one_wire_N_579[9]), .O(n34515));
    defparam i21466_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 i1_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n45), .I2(start), 
            .I3(GND_net), .O(n30278));
    defparam i1_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i17247_3_lut (.I0(n30278), .I1(n46404), .I2(\state[0] ), .I3(GND_net), 
            .O(n30301));   // verilog/neopixel.v(16[20:25])
    defparam i17247_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_2_lut_adj_1622 (.I0(\neo_pixel_transmitter.done ), .I1(n34515), 
            .I2(GND_net), .I3(GND_net), .O(n60));
    defparam i1_2_lut_adj_1622.LUT_INIT = 16'hbbbb;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1414_3_lut (.I0(n2000), .I1(n2060[25]), .I2(n2027), 
            .I3(GND_net), .O(n2099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21069_2_lut_3_lut_4_lut (.I0(bit_ctr[27]), .I1(n25173), .I2(n27956), 
            .I3(bit_ctr[26]), .O(n56));   // verilog/neopixel.v(22[26:36])
    defparam i21069_2_lut_3_lut_4_lut.LUT_INIT = 16'h7aff;
    SB_LUT4 mod_5_i1411_3_lut (.I0(n1997), .I1(n2060[28]), .I2(n2027), 
            .I3(GND_net), .O(n2096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1410_3_lut (.I0(n1996), .I1(n2060[29]), .I2(n2027), 
            .I3(GND_net), .O(n2095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut (.I0(n1007), .I1(n971[30]), .I2(n2_adj_4905), 
            .I3(GND_net), .O(n8_adj_4906));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 mod_5_i1412_3_lut (.I0(n1998), .I1(n2060[27]), .I2(n2027), 
            .I3(GND_net), .O(n2097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1423_3_lut (.I0(n2009), .I1(n2060[16]), .I2(n2027), 
            .I3(GND_net), .O(n2108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1418_3_lut (.I0(n2004), .I1(n2060[21]), .I2(n2027), 
            .I3(GND_net), .O(n2103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1417_3_lut (.I0(n2003), .I1(n2060[22]), .I2(n2027), 
            .I3(GND_net), .O(n2102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1413_3_lut (.I0(n1999), .I1(n2060[26]), .I2(n2027), 
            .I3(GND_net), .O(n2098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1421_3_lut (.I0(n2007), .I1(n2060[18]), .I2(n2027), 
            .I3(GND_net), .O(n2106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17641_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n27956));   // verilog/neopixel.v(18[12:19])
    defparam i17641_3_lut_4_lut.LUT_INIT = 16'hdb6d;
    SB_LUT4 bit_ctr_0__bdd_4_lut_34372 (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n49293));
    defparam bit_ctr_0__bdd_4_lut_34372.LUT_INIT = 16'he4aa;
    SB_LUT4 mod_5_i1415_3_lut (.I0(n2001), .I1(n2060[24]), .I2(n2027), 
            .I3(GND_net), .O(n2100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1416_3_lut (.I0(n2002), .I1(n2060[23]), .I2(n2027), 
            .I3(GND_net), .O(n2101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1419_3_lut (.I0(n2005), .I1(n2060[20]), .I2(n2027), 
            .I3(GND_net), .O(n2104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1422_3_lut (.I0(n2008), .I1(n2060[17]), .I2(n2027), 
            .I3(GND_net), .O(n2107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1420_3_lut (.I0(n2006), .I1(n2060[19]), .I2(n2027), 
            .I3(GND_net), .O(n2105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1424_3_lut (.I0(bit_ctr[15]), .I1(n2060[15]), .I2(n2027), 
            .I3(GND_net), .O(n2109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1409_3_lut (.I0(n1995), .I1(n2060[30]), .I2(n2027), 
            .I3(GND_net), .O(n2094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1623 (.I0(n2094), .I1(n2093), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4907));
    defparam i1_2_lut_adj_1623.LUT_INIT = 16'heeee;
    SB_LUT4 i21355_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n34401));
    defparam i21355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17643_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n25173));   // verilog/neopixel.v(18[12:19])
    defparam i17643_3_lut_4_lut.LUT_INIT = 16'hb6db;
    SB_LUT4 i13_4_lut_adj_1624 (.I0(n2105), .I1(n2107), .I2(n2104), .I3(n18_adj_4907), 
            .O(n30_adj_4908));
    defparam i13_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1625 (.I0(n2101), .I1(n2100), .I2(n2106), .I3(n2098), 
            .O(n28_adj_4909));
    defparam i11_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1626 (.I0(n2102), .I1(n2103), .I2(n34401), .I3(n2108), 
            .O(n29_adj_4910));
    defparam i12_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1627 (.I0(n2097), .I1(n2095), .I2(n2096), .I3(n2099), 
            .O(n27_adj_4911));
    defparam i10_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1628 (.I0(n27_adj_4911), .I1(n29_adj_4910), .I2(n28_adj_4909), 
            .I3(n30_adj_4908), .O(n2126));
    defparam i16_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 n49293_bdd_4_lut (.I0(n49293), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n49296));
    defparam n49293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF timer_1547__i2 (.Q(timer[2]), .C(CLK_c), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i3 (.Q(timer[3]), .C(CLK_c), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i4 (.Q(timer[4]), .C(CLK_c), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i5 (.Q(timer[5]), .C(CLK_c), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i6 (.Q(timer[6]), .C(CLK_c), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i7 (.Q(timer[7]), .C(CLK_c), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i8 (.Q(timer[8]), .C(CLK_c), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i9 (.Q(timer[9]), .C(CLK_c), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i10 (.Q(timer[10]), .C(CLK_c), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i11 (.Q(timer[11]), .C(CLK_c), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i12 (.Q(timer[12]), .C(CLK_c), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i13 (.Q(timer[13]), .C(CLK_c), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i14 (.Q(timer[14]), .C(CLK_c), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i15 (.Q(timer[15]), .C(CLK_c), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i16 (.Q(timer[16]), .C(CLK_c), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i17 (.Q(timer[17]), .C(CLK_c), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i18 (.Q(timer[18]), .C(CLK_c), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i19 (.Q(timer[19]), .C(CLK_c), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i20 (.Q(timer[20]), .C(CLK_c), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i21 (.Q(timer[21]), .C(CLK_c), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i22 (.Q(timer[22]), .C(CLK_c), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i23 (.Q(timer[23]), .C(CLK_c), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i24 (.Q(timer[24]), .C(CLK_c), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i25 (.Q(timer[25]), .C(CLK_c), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i26 (.Q(timer[26]), .C(CLK_c), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i27 (.Q(timer[27]), .C(CLK_c), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i28 (.Q(timer[28]), .C(CLK_c), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i29 (.Q(timer[29]), .C(CLK_c), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i30 (.Q(timer[30]), .C(CLK_c), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1547__i31 (.Q(timer[31]), .C(CLK_c), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n28163));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1344_3_lut (.I0(n1898), .I1(n1961[28]), .I2(n1928), 
            .I3(GND_net), .O(n1997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1343_3_lut (.I0(n1897), .I1(n1961[29]), .I2(n1928), 
            .I3(GND_net), .O(n1996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1342_3_lut (.I0(n1896), .I1(n1961[30]), .I2(n1928), 
            .I3(GND_net), .O(n1995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1346_3_lut (.I0(n1900), .I1(n1961[26]), .I2(n1928), 
            .I3(GND_net), .O(n1999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1350_3_lut (.I0(n1904), .I1(n1961[22]), .I2(n1928), 
            .I3(GND_net), .O(n2003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1347_3_lut (.I0(n1901), .I1(n1961[25]), .I2(n1928), 
            .I3(GND_net), .O(n2000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1355_3_lut (.I0(n1909), .I1(n1961[17]), .I2(n1928), 
            .I3(GND_net), .O(n2008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1349_3_lut (.I0(n1903), .I1(n1961[23]), .I2(n1928), 
            .I3(GND_net), .O(n2002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1345_3_lut (.I0(n1899), .I1(n1961[27]), .I2(n1928), 
            .I3(GND_net), .O(n1998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1352_3_lut (.I0(n1906), .I1(n1961[20]), .I2(n1928), 
            .I3(GND_net), .O(n2005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1348_3_lut (.I0(n1902), .I1(n1961[24]), .I2(n1928), 
            .I3(GND_net), .O(n2001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1353_3_lut (.I0(n1907), .I1(n1961[19]), .I2(n1928), 
            .I3(GND_net), .O(n2006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1354_3_lut (.I0(n1908), .I1(n1961[18]), .I2(n1928), 
            .I3(GND_net), .O(n2007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1351_3_lut (.I0(n1905), .I1(n1961[21]), .I2(n1928), 
            .I3(GND_net), .O(n2004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1356_3_lut (.I0(bit_ctr[16]), .I1(n1961[16]), .I2(n1928), 
            .I3(GND_net), .O(n2009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21353_2_lut (.I0(bit_ctr[15]), .I1(n2009), .I2(GND_net), 
            .I3(GND_net), .O(n34399));
    defparam i21353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1629 (.I0(n2004), .I1(n2007), .I2(n2006), .I3(n2001), 
            .O(n28_adj_4915));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1630 (.I0(n2005), .I1(n34399), .I2(n1998), .I3(n2002), 
            .O(n26_adj_4916));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1631 (.I0(n2008), .I1(n2000), .I2(n2003), .I3(n1999), 
            .O(n27_adj_4917));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1995), .I1(n1996), .I2(n1994), .I3(n1997), 
            .O(n25_adj_4918));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1632 (.I0(n25_adj_4918), .I1(n27_adj_4917), .I2(n26_adj_4916), 
            .I3(n28_adj_4915), .O(n2027));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1284_3_lut (.I0(n1806), .I1(n1862[21]), .I2(n1829), 
            .I3(GND_net), .O(n1905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1281_3_lut (.I0(n1803), .I1(n1862[24]), .I2(n1829), 
            .I3(GND_net), .O(n1902));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1280_3_lut (.I0(n1802), .I1(n1862[25]), .I2(n1829), 
            .I3(GND_net), .O(n1901));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1279_3_lut (.I0(n1801), .I1(n1862[26]), .I2(n1829), 
            .I3(GND_net), .O(n1900));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1277_3_lut (.I0(n1799), .I1(n1862[28]), .I2(n1829), 
            .I3(GND_net), .O(n1898));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1278_3_lut (.I0(n1800), .I1(n1862[27]), .I2(n1829), 
            .I3(GND_net), .O(n1899));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1276_3_lut (.I0(n1798), .I1(n1862[29]), .I2(n1829), 
            .I3(GND_net), .O(n1897));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1275_3_lut (.I0(n1797), .I1(n1862[30]), .I2(n1829), 
            .I3(GND_net), .O(n1896));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1287_3_lut (.I0(n1809), .I1(n1862[18]), .I2(n1829), 
            .I3(GND_net), .O(n1908));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1285_3_lut (.I0(n1807), .I1(n1862[20]), .I2(n1829), 
            .I3(GND_net), .O(n1906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1286_3_lut (.I0(n1808), .I1(n1862[19]), .I2(n1829), 
            .I3(GND_net), .O(n1907));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1282_3_lut (.I0(n1804), .I1(n1862[23]), .I2(n1829), 
            .I3(GND_net), .O(n1903));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1288_3_lut (.I0(bit_ctr[17]), .I1(n1862[17]), .I2(n1829), 
            .I3(GND_net), .O(n1909));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1283_3_lut (.I0(n1805), .I1(n1862[22]), .I2(n1829), 
            .I3(GND_net), .O(n1904));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1633 (.I0(bit_ctr[16]), .I1(n1904), .I2(n1909), 
            .I3(GND_net), .O(n20_adj_4919));
    defparam i5_3_lut_adj_1633.LUT_INIT = 16'hecec;
    SB_LUT4 i11_4_lut_adj_1634 (.I0(n1903), .I1(n1907), .I2(n1906), .I3(n1908), 
            .O(n26_adj_4920));
    defparam i11_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1635 (.I0(n1896), .I1(n1895), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4921));
    defparam i1_2_lut_adj_1635.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1636 (.I0(n1897), .I1(n1899), .I2(n1898), .I3(n1900), 
            .O(n24_adj_4922));
    defparam i9_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1637 (.I0(n1901), .I1(n26_adj_4920), .I2(n20_adj_4919), 
            .I3(n1902), .O(n28_adj_4923));
    defparam i13_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1638 (.I0(n1905), .I1(n28_adj_4923), .I2(n24_adj_4922), 
            .I3(n16_adj_4921), .O(n1928));
    defparam i14_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1547_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n38535), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1547_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n38534), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_32 (.CI(n38534), .I0(GND_net), .I1(timer[30]), 
            .CO(n38535));
    SB_LUT4 timer_1547_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n38533), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_31 (.CI(n38533), .I0(GND_net), .I1(timer[29]), 
            .CO(n38534));
    SB_LUT4 timer_1547_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n38532), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_30 (.CI(n38532), .I0(GND_net), .I1(timer[28]), 
            .CO(n38533));
    SB_LUT4 timer_1547_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n38531), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_29 (.CI(n38531), .I0(GND_net), .I1(timer[27]), 
            .CO(n38532));
    SB_LUT4 timer_1547_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n38530), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_28 (.CI(n38530), .I0(GND_net), .I1(timer[26]), 
            .CO(n38531));
    SB_LUT4 timer_1547_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n38529), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_27 (.CI(n38529), .I0(GND_net), .I1(timer[25]), 
            .CO(n38530));
    SB_LUT4 timer_1547_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n38528), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_26 (.CI(n38528), .I0(GND_net), .I1(timer[24]), 
            .CO(n38529));
    SB_LUT4 timer_1547_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n38527), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_25 (.CI(n38527), .I0(GND_net), .I1(timer[23]), 
            .CO(n38528));
    SB_LUT4 timer_1547_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n38526), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_24 (.CI(n38526), .I0(GND_net), .I1(timer[22]), 
            .CO(n38527));
    SB_LUT4 timer_1547_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n38525), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_23 (.CI(n38525), .I0(GND_net), .I1(timer[21]), 
            .CO(n38526));
    SB_LUT4 timer_1547_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n38524), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_22 (.CI(n38524), .I0(GND_net), .I1(timer[20]), 
            .CO(n38525));
    SB_LUT4 timer_1547_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n38523), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_21 (.CI(n38523), .I0(GND_net), .I1(timer[19]), 
            .CO(n38524));
    SB_LUT4 timer_1547_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n38522), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_20 (.CI(n38522), .I0(GND_net), .I1(timer[18]), 
            .CO(n38523));
    SB_LUT4 timer_1547_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n38521), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_19 (.CI(n38521), .I0(GND_net), .I1(timer[17]), 
            .CO(n38522));
    SB_LUT4 timer_1547_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n38520), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_18 (.CI(n38520), .I0(GND_net), .I1(timer[16]), 
            .CO(n38521));
    SB_LUT4 timer_1547_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n38519), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_17 (.CI(n38519), .I0(GND_net), .I1(timer[15]), 
            .CO(n38520));
    SB_LUT4 timer_1547_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n38518), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_16 (.CI(n38518), .I0(GND_net), .I1(timer[14]), 
            .CO(n38519));
    SB_LUT4 timer_1547_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n38517), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_15 (.CI(n38517), .I0(GND_net), .I1(timer[13]), 
            .CO(n38518));
    SB_LUT4 timer_1547_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n38516), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_14 (.CI(n38516), .I0(GND_net), .I1(timer[12]), 
            .CO(n38517));
    SB_LUT4 timer_1547_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n38515), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_13 (.CI(n38515), .I0(GND_net), .I1(timer[11]), 
            .CO(n38516));
    SB_LUT4 timer_1547_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n38514), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_12 (.CI(n38514), .I0(GND_net), .I1(timer[10]), 
            .CO(n38515));
    SB_LUT4 timer_1547_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n38513), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_11 (.CI(n38513), .I0(GND_net), .I1(timer[9]), 
            .CO(n38514));
    SB_LUT4 timer_1547_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n38512), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_10 (.CI(n38512), .I0(GND_net), .I1(timer[8]), 
            .CO(n38513));
    SB_LUT4 timer_1547_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n38511), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_9 (.CI(n38511), .I0(GND_net), .I1(timer[7]), 
            .CO(n38512));
    SB_LUT4 timer_1547_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n38510), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_8 (.CI(n38510), .I0(GND_net), .I1(timer[6]), 
            .CO(n38511));
    SB_LUT4 timer_1547_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n38509), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_7 (.CI(n38509), .I0(GND_net), .I1(timer[5]), 
            .CO(n38510));
    SB_LUT4 timer_1547_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n38508), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_6 (.CI(n38508), .I0(GND_net), .I1(timer[4]), 
            .CO(n38509));
    SB_LUT4 timer_1547_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n38507), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_5 (.CI(n38507), .I0(GND_net), .I1(timer[3]), 
            .CO(n38508));
    SB_LUT4 timer_1547_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n38506), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_4 (.CI(n38506), .I0(GND_net), .I1(timer[2]), 
            .CO(n38507));
    SB_LUT4 timer_1547_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n38505), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_3 (.CI(n38505), .I0(GND_net), .I1(timer[1]), 
            .CO(n38506));
    SB_LUT4 timer_1547_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1547_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1547_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n38505));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n38504), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n38503), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n38503), .I0(n1203), .I1(n1235), .CO(n38504));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n38502), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n38502), .I0(n1204), .I1(n1235), .CO(n38503));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n38501), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n38501), .I0(n1205), .I1(n1235), .CO(n38502));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n38500), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n38500), .I0(n1206), .I1(n1235), .CO(n38501));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n38499), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n38499), .I0(n1207), .I1(n1235), .CO(n38500));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n38498), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n38498), .I0(n1208), .I1(n1235), .CO(n38499));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n49249), 
            .I3(n38497), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n38497), .I0(n1209), .I1(n49249), .CO(n38498));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n49249), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n49249), 
            .CO(n38497));
    SB_LUT4 mod_5_i1219_3_lut (.I0(n1709), .I1(n1763[19]), .I2(n1730), 
            .I3(GND_net), .O(n1808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1216_3_lut (.I0(n1706), .I1(n1763[22]), .I2(n1730), 
            .I3(GND_net), .O(n1805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1215_3_lut (.I0(n1705), .I1(n1763[23]), .I2(n1730), 
            .I3(GND_net), .O(n1804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1212_3_lut (.I0(n1702), .I1(n1763[26]), .I2(n1730), 
            .I3(GND_net), .O(n1801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1213_3_lut (.I0(n1703), .I1(n1763[25]), .I2(n1730), 
            .I3(GND_net), .O(n1802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1217_3_lut (.I0(n1707), .I1(n1763[21]), .I2(n1730), 
            .I3(GND_net), .O(n1806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1211_3_lut (.I0(n1701), .I1(n1763[27]), .I2(n1730), 
            .I3(GND_net), .O(n1800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1218_3_lut (.I0(n1708), .I1(n1763[20]), .I2(n1730), 
            .I3(GND_net), .O(n1807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1214_3_lut (.I0(n1704), .I1(n1763[24]), .I2(n1730), 
            .I3(GND_net), .O(n1803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1209_3_lut (.I0(n1699), .I1(n1763[29]), .I2(n1730), 
            .I3(GND_net), .O(n1798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1208_3_lut (.I0(n1698), .I1(n1763[30]), .I2(n1730), 
            .I3(GND_net), .O(n1797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1220_3_lut (.I0(bit_ctr[18]), .I1(n1763[18]), .I2(n1730), 
            .I3(GND_net), .O(n1809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1210_3_lut (.I0(n1700), .I1(n1763[28]), .I2(n1730), 
            .I3(GND_net), .O(n1799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1639 (.I0(n1807), .I1(n1800), .I2(n1806), .I3(n1802), 
            .O(n24_adj_4924));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n1799), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n17_adj_4925));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i8_4_lut (.I0(n1797), .I1(n1798), .I2(n1796), .I3(n1803), 
            .O(n22_adj_4926));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1640 (.I0(n17_adj_4925), .I1(n24_adj_4924), .I2(n1801), 
            .I3(n1804), .O(n26_adj_4927));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1641 (.I0(n1805), .I1(n26_adj_4927), .I2(n22_adj_4926), 
            .I3(n1808), .O(n1829));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1151_3_lut (.I0(n1609), .I1(n1664[20]), .I2(n1631), 
            .I3(GND_net), .O(n1708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1148_3_lut (.I0(n1606), .I1(n1664[23]), .I2(n1631), 
            .I3(GND_net), .O(n1705));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1147_3_lut (.I0(n1605), .I1(n1664[24]), .I2(n1631), 
            .I3(GND_net), .O(n1704));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1146_3_lut (.I0(n1604), .I1(n1664[25]), .I2(n1631), 
            .I3(GND_net), .O(n1703));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1141_3_lut (.I0(n1599), .I1(n1664[30]), .I2(n1631), 
            .I3(GND_net), .O(n1698));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1150_3_lut (.I0(n1608), .I1(n1664[21]), .I2(n1631), 
            .I3(GND_net), .O(n1707));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1145_3_lut (.I0(n1603), .I1(n1664[26]), .I2(n1631), 
            .I3(GND_net), .O(n1702));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1143_3_lut (.I0(n1601), .I1(n1664[28]), .I2(n1631), 
            .I3(GND_net), .O(n1700));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1144_3_lut (.I0(n1602), .I1(n1664[27]), .I2(n1631), 
            .I3(GND_net), .O(n1701));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1142_3_lut (.I0(n1600), .I1(n1664[29]), .I2(n1631), 
            .I3(GND_net), .O(n1699));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1152_3_lut (.I0(bit_ctr[19]), .I1(n1664[19]), .I2(n1631), 
            .I3(GND_net), .O(n1709));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1149_3_lut (.I0(n1607), .I1(n1664[22]), .I2(n1631), 
            .I3(GND_net), .O(n1706));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1642 (.I0(bit_ctr[18]), .I1(n1706), .I2(n1709), 
            .I3(GND_net), .O(n18_adj_4928));
    defparam i5_3_lut_adj_1642.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1643 (.I0(n1699), .I1(n1701), .I2(n1700), .I3(n1702), 
            .O(n21_adj_4929));
    defparam i8_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1644 (.I0(n1707), .I1(n1698), .I2(n1697), .I3(GND_net), 
            .O(n20_adj_4930));
    defparam i7_3_lut_adj_1644.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1645 (.I0(n21_adj_4929), .I1(n1703), .I2(n18_adj_4928), 
            .I3(n1704), .O(n24_adj_4931));
    defparam i11_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1646 (.I0(n1705), .I1(n24_adj_4931), .I2(n20_adj_4930), 
            .I3(n1708), .O(n1730));
    defparam i12_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1083_3_lut (.I0(n1509), .I1(n1565[21]), .I2(n1532), 
            .I3(GND_net), .O(n1608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1077_3_lut (.I0(n1503), .I1(n1565[27]), .I2(n1532), 
            .I3(GND_net), .O(n1602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1074_3_lut (.I0(n1500), .I1(n1565[30]), .I2(n1532), 
            .I3(GND_net), .O(n1599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1076_3_lut (.I0(n1502), .I1(n1565[28]), .I2(n1532), 
            .I3(GND_net), .O(n1601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1079_3_lut (.I0(n1505), .I1(n1565[25]), .I2(n1532), 
            .I3(GND_net), .O(n1604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1081_3_lut (.I0(n1507), .I1(n1565[23]), .I2(n1532), 
            .I3(GND_net), .O(n1606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1080_3_lut (.I0(n1506), .I1(n1565[24]), .I2(n1532), 
            .I3(GND_net), .O(n1605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1078_3_lut (.I0(n1504), .I1(n1565[26]), .I2(n1532), 
            .I3(GND_net), .O(n1603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1075_3_lut (.I0(n1501), .I1(n1565[29]), .I2(n1532), 
            .I3(GND_net), .O(n1600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1015_3_lut (.I0(n1409), .I1(n1466[22]), .I2(n1433), 
            .I3(GND_net), .O(n1508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1014_3_lut (.I0(n1408), .I1(n1466[23]), .I2(n1433), 
            .I3(GND_net), .O(n1507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1016_3_lut (.I0(bit_ctr[21]), .I1(n1466[21]), .I2(n1433), 
            .I3(GND_net), .O(n1509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1012_3_lut (.I0(n1406), .I1(n1466[25]), .I2(n1433), 
            .I3(GND_net), .O(n1505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1007_3_lut (.I0(n1401), .I1(n1466[30]), .I2(n1433), 
            .I3(GND_net), .O(n1500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1013_3_lut (.I0(n1407), .I1(n1466[24]), .I2(n1433), 
            .I3(GND_net), .O(n1506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1011_3_lut (.I0(n1405), .I1(n1466[26]), .I2(n1433), 
            .I3(GND_net), .O(n1504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1009_3_lut (.I0(n1403), .I1(n1466[28]), .I2(n1433), 
            .I3(GND_net), .O(n1502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1010_3_lut (.I0(n1404), .I1(n1466[27]), .I2(n1433), 
            .I3(GND_net), .O(n1503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1008_3_lut (.I0(n1402), .I1(n1466[29]), .I2(n1433), 
            .I3(GND_net), .O(n1501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1647 (.I0(n1501), .I1(n1503), .I2(n1502), .I3(n1504), 
            .O(n18_adj_4932));
    defparam i7_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1648 (.I0(n1506), .I1(n18_adj_4932), .I2(n1500), 
            .I3(n1499), .O(n20_adj_4933));
    defparam i9_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1649 (.I0(n1505), .I1(bit_ctr[20]), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4934));
    defparam i4_3_lut_adj_1649.LUT_INIT = 16'heaea;
    SB_LUT4 i10_4_lut_adj_1650 (.I0(n15_adj_4934), .I1(n20_adj_4933), .I2(n1507), 
            .I3(n1508), .O(n1532));
    defparam i10_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1084_3_lut (.I0(bit_ctr[20]), .I1(n1565[20]), .I2(n1532), 
            .I3(GND_net), .O(n1609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1082_3_lut (.I0(n1508), .I1(n1565[22]), .I2(n1532), 
            .I3(GND_net), .O(n1607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(bit_ctr[19]), .I1(n1607), .I2(n1609), .I3(GND_net), 
            .O(n14_adj_4935));   // verilog/neopixel.v(22[26:36])
    defparam i2_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1651 (.I0(n1600), .I1(n1603), .I2(n1605), .I3(n1606), 
            .O(n20_adj_4936));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1604), .I1(n1601), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4937));   // verilog/neopixel.v(22[26:36])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1652 (.I0(n1599), .I1(n20_adj_4936), .I2(n14_adj_4935), 
            .I3(n1598), .O(n22_adj_4938));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1653 (.I0(n1602), .I1(n22_adj_4938), .I2(n18_adj_4937), 
            .I3(n1608), .O(n1631));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i34292_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49245));
    defparam i34292_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21341_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n34387));
    defparam i21341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1654 (.I0(n1106), .I1(n1103), .I2(n1108), .I3(n34387), 
            .O(n12_adj_4939));
    defparam i5_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1107), .I1(n12_adj_4939), .I2(n1105), .I3(n1104), 
            .O(n1136));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(one_wire_N_579[3]), .I1(n4_adj_4893), 
            .I2(n147), .I3(GND_net), .O(n45));   // verilog/neopixel.v(6[16:24])
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'hf8f8;
    SB_LUT4 i34291_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49244));
    defparam i34291_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33785_2_lut (.I0(n971[28]), .I1(n2_adj_4905), .I2(GND_net), 
            .I3(GND_net), .O(n48738));   // verilog/neopixel.v(22[26:36])
    defparam i33785_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33784_2_lut (.I0(n971[29]), .I1(n2_adj_4905), .I2(GND_net), 
            .I3(GND_net), .O(n48737));   // verilog/neopixel.v(22[26:36])
    defparam i33784_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33839_2_lut (.I0(n971[30]), .I1(n2_adj_4905), .I2(GND_net), 
            .I3(GND_net), .O(n48792));   // verilog/neopixel.v(22[26:36])
    defparam i33839_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_3_lut_adj_1656 (.I0(n147), .I1(one_wire_N_579[3]), 
            .I2(one_wire_N_579[2]), .I3(GND_net), .O(n30298));
    defparam i2_2_lut_3_lut_adj_1656.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_i673_3_lut (.I0(n27993), .I1(n971[29]), .I2(n2_adj_4905), 
            .I3(GND_net), .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i674_3_lut (.I0(n27950), .I1(n971[28]), .I2(n2_adj_4905), 
            .I3(GND_net), .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2_adj_4905), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n25171), .I1(n971[27]), .I2(n2_adj_4905), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1657 (.I0(n27950), .I1(n27993), .I2(n56), .I3(GND_net), 
            .O(n2_adj_4905));   // verilog/neopixel.v(22[26:36])
    defparam i1_4_lut_adj_1657.LUT_INIT = 16'h1010;
    SB_LUT4 i33912_2_lut (.I0(n971[31]), .I1(n2_adj_4905), .I2(GND_net), 
            .I3(GND_net), .O(n48865));   // verilog/neopixel.v(22[26:36])
    defparam i33912_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[0] ), .I1(n147), .I2(one_wire_N_579[3]), 
            .I3(n4_adj_4893), .O(n14));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i1_3_lut_adj_1658 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n7_adj_4940));
    defparam i1_3_lut_adj_1658.LUT_INIT = 16'heaea;
    SB_LUT4 i5_4_lut_adj_1659 (.I0(n48865), .I1(n7_adj_4940), .I2(n1006), 
            .I3(n8_adj_4906), .O(n1037));
    defparam i5_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i32703_2_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(one_wire_N_579[3]), .I3(one_wire_N_579[2]), .O(n47529));
    defparam i32703_2_lut_4_lut.LUT_INIT = 16'h4440;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32706_2_lut_4_lut (.I0(LED_c), .I1(bit_ctr[3]), .I2(bit_ctr[4]), 
            .I3(n40382), .O(n47530));
    defparam i32706_2_lut_4_lut.LUT_INIT = 16'haa80;
    SB_LUT4 i22_3_lut_4_lut (.I0(n113), .I1(n147), .I2(\state[1] ), .I3(\state[0] ), 
            .O(n11_adj_4883));   // verilog/neopixel.v(16[20:25])
    defparam i22_3_lut_4_lut.LUT_INIT = 16'h0fee;
    SB_LUT4 i1_2_lut_4_lut (.I0(n147), .I1(n4_adj_4823), .I2(start), .I3(\neo_pixel_transmitter.done ), 
            .O(n46404));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0e00;
    SB_LUT4 i32963_3_lut_3_lut (.I0(bit_ctr[27]), .I1(n25173), .I2(n27956), 
            .I3(GND_net), .O(n27950));   // verilog/neopixel.v(22[26:36])
    defparam i32963_3_lut_3_lut.LUT_INIT = 16'h1919;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i606_3_lut_4_lut_3_lut (.I0(bit_ctr[27]), .I1(n25173), 
            .I2(n27956), .I3(GND_net), .O(n27993));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i942_3_lut (.I0(n1304), .I1(n1367[28]), .I2(n1334), 
            .I3(GND_net), .O(n1403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i943_3_lut (.I0(n1305), .I1(n1367[27]), .I2(n1334), 
            .I3(GND_net), .O(n1404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i946_3_lut (.I0(n1308), .I1(n1367[24]), .I2(n1334), 
            .I3(GND_net), .O(n1407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i945_3_lut (.I0(n1307), .I1(n1367[25]), .I2(n1334), 
            .I3(GND_net), .O(n1406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i944_3_lut (.I0(n1306), .I1(n1367[26]), .I2(n1334), 
            .I3(GND_net), .O(n1405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i941_3_lut (.I0(n1303), .I1(n1367[29]), .I2(n1334), 
            .I3(GND_net), .O(n1402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1660 (.I0(n1307), .I1(n1302), .I2(n1301), .I3(GND_net), 
            .O(n14_adj_4941));   // verilog/neopixel.v(22[26:36])
    defparam i5_3_lut_adj_1660.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_2_lut_adj_1661 (.I0(n1305), .I1(n1306), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4942));   // verilog/neopixel.v(22[26:36])
    defparam i3_2_lut_adj_1661.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1662 (.I0(bit_ctr[22]), .I1(n14_adj_4941), .I2(n1308), 
            .I3(n1309), .O(n16_adj_4943));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1662.LUT_INIT = 16'hfefc;
    SB_LUT4 i8_4_lut_adj_1663 (.I0(n1303), .I1(n16_adj_4943), .I2(n12_adj_4942), 
            .I3(n1304), .O(n1334));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i940_3_lut (.I0(n1302), .I1(n1367[30]), .I2(n1334), 
            .I3(GND_net), .O(n1401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i947_3_lut (.I0(n1309), .I1(n1367[23]), .I2(n1334), 
            .I3(GND_net), .O(n1408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i948_3_lut (.I0(bit_ctr[22]), .I1(n1367[22]), .I2(n1334), 
            .I3(GND_net), .O(n1409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_1664 (.I0(n1408), .I1(n1401), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4944));   // verilog/neopixel.v(22[26:36])
    defparam i2_2_lut_adj_1664.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1665 (.I0(bit_ctr[21]), .I1(n12_adj_4944), .I2(n1400), 
            .I3(n1409), .O(n16_adj_4945));   // verilog/neopixel.v(22[26:36])
    defparam i6_4_lut_adj_1665.LUT_INIT = 16'hfefc;
    SB_LUT4 i7_4_lut_adj_1666 (.I0(n1402), .I1(n1405), .I2(n1406), .I3(n1407), 
            .O(n17_adj_4946));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1667 (.I0(n17_adj_4946), .I1(n1404), .I2(n16_adj_4945), 
            .I3(n1403), .O(n1433));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i32732_3_lut_4_lut (.I0(\state[0] ), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n34515), .O(n47534));   // verilog/neopixel.v(16[20:25])
    defparam i32732_3_lut_4_lut.LUT_INIT = 16'hcdcc;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47_3_lut_4_lut (.I0(one_wire_N_579[3]), .I1(n4_adj_4893), .I2(one_wire_N_579[2]), 
            .I3(\neo_pixel_transmitter.done ), .O(n42927));
    defparam i47_3_lut_4_lut.LUT_INIT = 16'hfa88;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1668 (.I0(n147), .I1(\state[1] ), .I2(start), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut_3_lut_adj_1668.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n34515), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n44951));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 bit_ctr_1__bdd_4_lut (.I0(bit_ctr[1]), .I1(n46746), .I2(n46747), 
            .I3(bit_ctr[2]), .O(n49251));
    defparam bit_ctr_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49251_bdd_4_lut (.I0(n49251), .I1(n46744), .I2(n46743), .I3(bit_ctr[2]), 
            .O(n49254));
    defparam n49251_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (\a_new[1] , ENCODER0_B_N_keep, 
            n1188, ENCODER0_A_N_keep, b_prev, n28221, n1152, direction_N_3807, 
            encoder0_position, GND_net, VCC_net) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    input ENCODER0_B_N_keep;
    input n1188;
    input ENCODER0_A_N_keep;
    output b_prev;
    input n28221;
    output n1152;
    output direction_N_3807;
    output [31:0]encoder0_position;
    input GND_net;
    input VCC_net;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire a_prev_N_3813, debounce_cnt, n28223, a_prev, n28222;
    wire [31:0]n133;
    
    wire direction_N_3806, n38643, n38642, n38641, n38640, n38639, 
        n38638, n38637, n38636, n38635, n38634, n38633, n38632, 
        n38631, n38630, n38629, n38628, n38627, n38626, n38625, 
        n38624, n38623, n38622, n38621, n38620, n38619, n38618, 
        n38617, n38616, n38615, n38614, n38613, direction_N_3810;
    
    SB_LUT4 i33586_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(57[8:58])
    defparam i33586_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1188), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1188), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1188), .D(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1188), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1188), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1188), .D(n28223));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1188), .D(n28222));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1152), .C(n1188), .D(n28221));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_1554__i0 (.Q(encoder0_position[0]), .C(n1188), .E(direction_N_3807), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_1554_add_4_33_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[31]), .I3(n38643), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15164_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n28223));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15164_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15163_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(b_new[1]), 
            .I3(b_prev), .O(n28222));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15163_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 position_1554_add_4_32_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[30]), .I3(n38642), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_32 (.CI(n38642), .I0(direction_N_3806), 
            .I1(encoder0_position[30]), .CO(n38643));
    SB_LUT4 position_1554_add_4_31_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[29]), .I3(n38641), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_31 (.CI(n38641), .I0(direction_N_3806), 
            .I1(encoder0_position[29]), .CO(n38642));
    SB_LUT4 position_1554_add_4_30_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[28]), .I3(n38640), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_30 (.CI(n38640), .I0(direction_N_3806), 
            .I1(encoder0_position[28]), .CO(n38641));
    SB_LUT4 position_1554_add_4_29_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[27]), .I3(n38639), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_29 (.CI(n38639), .I0(direction_N_3806), 
            .I1(encoder0_position[27]), .CO(n38640));
    SB_LUT4 position_1554_add_4_28_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[26]), .I3(n38638), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_28 (.CI(n38638), .I0(direction_N_3806), 
            .I1(encoder0_position[26]), .CO(n38639));
    SB_LUT4 position_1554_add_4_27_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[25]), .I3(n38637), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_27 (.CI(n38637), .I0(direction_N_3806), 
            .I1(encoder0_position[25]), .CO(n38638));
    SB_LUT4 position_1554_add_4_26_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[24]), .I3(n38636), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_26 (.CI(n38636), .I0(direction_N_3806), 
            .I1(encoder0_position[24]), .CO(n38637));
    SB_LUT4 position_1554_add_4_25_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[23]), .I3(n38635), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_25 (.CI(n38635), .I0(direction_N_3806), 
            .I1(encoder0_position[23]), .CO(n38636));
    SB_LUT4 position_1554_add_4_24_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[22]), .I3(n38634), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_24 (.CI(n38634), .I0(direction_N_3806), 
            .I1(encoder0_position[22]), .CO(n38635));
    SB_DFFE position_1554__i1 (.Q(encoder0_position[1]), .C(n1188), .E(direction_N_3807), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i2 (.Q(encoder0_position[2]), .C(n1188), .E(direction_N_3807), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i3 (.Q(encoder0_position[3]), .C(n1188), .E(direction_N_3807), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i4 (.Q(encoder0_position[4]), .C(n1188), .E(direction_N_3807), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i5 (.Q(encoder0_position[5]), .C(n1188), .E(direction_N_3807), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i6 (.Q(encoder0_position[6]), .C(n1188), .E(direction_N_3807), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i7 (.Q(encoder0_position[7]), .C(n1188), .E(direction_N_3807), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i8 (.Q(encoder0_position[8]), .C(n1188), .E(direction_N_3807), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i9 (.Q(encoder0_position[9]), .C(n1188), .E(direction_N_3807), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i10 (.Q(encoder0_position[10]), .C(n1188), .E(direction_N_3807), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i11 (.Q(encoder0_position[11]), .C(n1188), .E(direction_N_3807), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i12 (.Q(encoder0_position[12]), .C(n1188), .E(direction_N_3807), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i13 (.Q(encoder0_position[13]), .C(n1188), .E(direction_N_3807), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i14 (.Q(encoder0_position[14]), .C(n1188), .E(direction_N_3807), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i15 (.Q(encoder0_position[15]), .C(n1188), .E(direction_N_3807), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i16 (.Q(encoder0_position[16]), .C(n1188), .E(direction_N_3807), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i17 (.Q(encoder0_position[17]), .C(n1188), .E(direction_N_3807), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i18 (.Q(encoder0_position[18]), .C(n1188), .E(direction_N_3807), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i19 (.Q(encoder0_position[19]), .C(n1188), .E(direction_N_3807), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i20 (.Q(encoder0_position[20]), .C(n1188), .E(direction_N_3807), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i21 (.Q(encoder0_position[21]), .C(n1188), .E(direction_N_3807), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i22 (.Q(encoder0_position[22]), .C(n1188), .E(direction_N_3807), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i23 (.Q(encoder0_position[23]), .C(n1188), .E(direction_N_3807), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i24 (.Q(encoder0_position[24]), .C(n1188), .E(direction_N_3807), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i25 (.Q(encoder0_position[25]), .C(n1188), .E(direction_N_3807), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i26 (.Q(encoder0_position[26]), .C(n1188), .E(direction_N_3807), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i27 (.Q(encoder0_position[27]), .C(n1188), .E(direction_N_3807), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i28 (.Q(encoder0_position[28]), .C(n1188), .E(direction_N_3807), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i29 (.Q(encoder0_position[29]), .C(n1188), .E(direction_N_3807), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i30 (.Q(encoder0_position[30]), .C(n1188), .E(direction_N_3807), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1554__i31 (.Q(encoder0_position[31]), .C(n1188), .E(direction_N_3807), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_1554_add_4_23_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[21]), .I3(n38633), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_23 (.CI(n38633), .I0(direction_N_3806), 
            .I1(encoder0_position[21]), .CO(n38634));
    SB_LUT4 position_1554_add_4_22_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[20]), .I3(n38632), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_22 (.CI(n38632), .I0(direction_N_3806), 
            .I1(encoder0_position[20]), .CO(n38633));
    SB_LUT4 position_1554_add_4_21_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[19]), .I3(n38631), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_21 (.CI(n38631), .I0(direction_N_3806), 
            .I1(encoder0_position[19]), .CO(n38632));
    SB_LUT4 position_1554_add_4_20_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[18]), .I3(n38630), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_20 (.CI(n38630), .I0(direction_N_3806), 
            .I1(encoder0_position[18]), .CO(n38631));
    SB_LUT4 position_1554_add_4_19_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[17]), .I3(n38629), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_19 (.CI(n38629), .I0(direction_N_3806), 
            .I1(encoder0_position[17]), .CO(n38630));
    SB_LUT4 position_1554_add_4_18_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[16]), .I3(n38628), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_18 (.CI(n38628), .I0(direction_N_3806), 
            .I1(encoder0_position[16]), .CO(n38629));
    SB_LUT4 position_1554_add_4_17_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[15]), .I3(n38627), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_17 (.CI(n38627), .I0(direction_N_3806), 
            .I1(encoder0_position[15]), .CO(n38628));
    SB_LUT4 position_1554_add_4_16_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[14]), .I3(n38626), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_16 (.CI(n38626), .I0(direction_N_3806), 
            .I1(encoder0_position[14]), .CO(n38627));
    SB_LUT4 position_1554_add_4_15_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[13]), .I3(n38625), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_15 (.CI(n38625), .I0(direction_N_3806), 
            .I1(encoder0_position[13]), .CO(n38626));
    SB_LUT4 position_1554_add_4_14_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[12]), .I3(n38624), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_14 (.CI(n38624), .I0(direction_N_3806), 
            .I1(encoder0_position[12]), .CO(n38625));
    SB_LUT4 position_1554_add_4_13_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[11]), .I3(n38623), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_13 (.CI(n38623), .I0(direction_N_3806), 
            .I1(encoder0_position[11]), .CO(n38624));
    SB_LUT4 position_1554_add_4_12_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[10]), .I3(n38622), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_12 (.CI(n38622), .I0(direction_N_3806), 
            .I1(encoder0_position[10]), .CO(n38623));
    SB_LUT4 position_1554_add_4_11_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[9]), .I3(n38621), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_11 (.CI(n38621), .I0(direction_N_3806), 
            .I1(encoder0_position[9]), .CO(n38622));
    SB_LUT4 position_1554_add_4_10_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[8]), .I3(n38620), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_10 (.CI(n38620), .I0(direction_N_3806), 
            .I1(encoder0_position[8]), .CO(n38621));
    SB_LUT4 position_1554_add_4_9_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[7]), .I3(n38619), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_9 (.CI(n38619), .I0(direction_N_3806), 
            .I1(encoder0_position[7]), .CO(n38620));
    SB_LUT4 position_1554_add_4_8_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[6]), .I3(n38618), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_8 (.CI(n38618), .I0(direction_N_3806), 
            .I1(encoder0_position[6]), .CO(n38619));
    SB_LUT4 position_1554_add_4_7_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[5]), .I3(n38617), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_7 (.CI(n38617), .I0(direction_N_3806), 
            .I1(encoder0_position[5]), .CO(n38618));
    SB_LUT4 position_1554_add_4_6_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[4]), .I3(n38616), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_6 (.CI(n38616), .I0(direction_N_3806), 
            .I1(encoder0_position[4]), .CO(n38617));
    SB_LUT4 position_1554_add_4_5_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[3]), .I3(n38615), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_5 (.CI(n38615), .I0(direction_N_3806), 
            .I1(encoder0_position[3]), .CO(n38616));
    SB_LUT4 position_1554_add_4_4_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[2]), .I3(n38614), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_4 (.CI(n38614), .I0(direction_N_3806), 
            .I1(encoder0_position[2]), .CO(n38615));
    SB_LUT4 position_1554_add_4_3_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[1]), .I3(n38613), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_3 (.CI(n38613), .I0(direction_N_3806), 
            .I1(encoder0_position[1]), .CO(n38614));
    SB_LUT4 position_1554_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1554_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1554_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n38613));
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3810));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3810), 
            .I3(\a_new[1] ), .O(direction_N_3807));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3806));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (PWMLimit, GND_net, \Ki[8] , \Ki[1] , \Ki[0] , 
            \Ki[2] , \Ki[3] , \Kp[2] , \Ki[4] , \Kp[1] , \Kp[0] , 
            \Ki[5] , \Kp[6] , \Ki[6] , \Ki[7] , \Ki[9] , \Kp[7] , 
            \Kp[3] , \Kp[8] , \Kp[4] , \Kp[5] , \Kp[9] , \Ki[10] , 
            \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , setpoint, 
            motor_state, \Kp[15] , \Ki[11] , \Ki[12] , \Ki[13] , duty, 
            clk32MHz, \Ki[14] , \Ki[15] , IntegralLimit, VCC_net, 
            n49248) /* synthesis syn_module_defined=1 */ ;
    input [23:0]PWMLimit;
    input GND_net;
    input \Ki[8] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Kp[2] ;
    input \Ki[4] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Ki[5] ;
    input \Kp[6] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[9] ;
    input \Kp[7] ;
    input \Kp[3] ;
    input \Kp[8] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[9] ;
    input \Ki[10] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input \Kp[15] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    output [23:0]duty;
    input clk32MHz;
    input \Ki[14] ;
    input \Ki[15] ;
    input [23:0]IntegralLimit;
    input VCC_net;
    output n49248;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]duty_23__N_3647;
    
    wire duty_23__N_3671;
    wire [23:0]duty_23__N_3548;
    wire [23:0]duty_23__N_3672;
    wire [23:0]n257;
    
    wire n256;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3572 ;
    
    wire n630, n116, n47, n189, n262;
    wire [23:0]n1;
    
    wire n168, n335, n74, n5, \PID_CONTROLLER.integral_23__N_3620 ;
    wire [23:0]n3616;
    
    wire n408, n454, n481, n554, n627, n700, n527, n113, n241, 
        n44, n186, n259_adj_4401, n332, n600, n314, n147, n405, 
        n387, n478, n551, n673, n624, n697, n770, n110, n41, 
        n460, n220, n293, n366, n533, n606, n679, n439, n752, 
        n512, n110_adj_4403, n41_adj_4404, n183, n256_adj_4405, n825, 
        n329, n402, n585, n475, n658, n898, n731, n548, n971, 
        n804, n621, n877, n694, n1044;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n37312, n37396, n37397, n767, n950, n1117, n1023, n840, 
        n1096, n92, n23, n37395, n165, n37313, n37311, n238, 
        n311, n37394, n384, n183_adj_4406, n256_adj_4407, n457, 
        n530, n603, n329_adj_4408, n402_adj_4409, n475_adj_4410, n548_adj_4411, 
        n621_adj_4412, n676, n694_adj_4413, n767_adj_4414, n840_adj_4415, 
        n746, n125, n56, n819, n198, n271, n344, n417, n6_adj_4416;
    wire [3:0]n19032;
    wire [4:0]n18983;
    
    wire n892, n749;
    wire [1:0]n19080;
    
    wire n822, n37393, n4_adj_4417;
    wire [2:0]n19063;
    
    wire n490, n12_adj_4418, n8_adj_4419, n11_adj_4420, n6_adj_4421, 
        n37310, n36954, n18, n13_adj_4422, n4_adj_4423, n44192, 
        n895, n965, n107, n38, n1038, n180, n968, n253, n326, 
        n1111, n399, n1041, n472, n545, n618, n691, n764, n837, 
        n910, n104, n35, n177, n250, n86, n17, n323, n159, 
        n396, n469, n232, n542, n615, n305, n1114, n37309, n688, 
        n761, n834, n907, n980, n378, n122, n53, n195, n268, 
        n39, n41_adj_4424, n45, n37, n341, n414, n451, n487, 
        n560, n29, n31, n43, n23_adj_4425, n101, n32, n174, 
        n524, n247, n320, n25_adj_4426, n393, n35_adj_4427, n11_adj_4428, 
        n13_adj_4429, n15, n27, n33, n9_adj_4430, n17_adj_4431, 
        n19_adj_4432, n21_adj_4433, n47880, n47874, n12_adj_4434, 
        n10_adj_4435, n30, n47890, n48128, n48124, n48402, n48242, 
        n48445, n16, n6_adj_4436, n48328, n48329, n8_adj_4437, n24_adj_4438, 
        n47860, n47858, n48308, n48004, n4_adj_4439, n48326, n48327, 
        n47870, n47868, n48412, n48006, n48482, n48483, n48462, 
        n47862, n48430, n48012, n48432, n41_adj_4440, n39_adj_4442, 
        n45_adj_4443, n43_adj_4444, n37_adj_4445, n29_adj_4446, n31_adj_4447, 
        n23_adj_4448, n25_adj_4449, n35_adj_4450, n33_adj_4451, n11_adj_4452, 
        n13_adj_4453, n15_adj_4454, n27_adj_4456, n9_adj_4457, n17_adj_4458, 
        n19_adj_4459, n21_adj_4461, n47845, n47838, n12_adj_4462, 
        n10_adj_4463, n30_adj_4464, n37392, n47855, n48088;
    wire [16:0]n15535;
    wire [15:0]n16112;
    
    wire n38071, n38070, n48082, n48396, n48224, n48443, n16_adj_4465, 
        n597, n466, n6_adj_4466, n48320, n539, n612, n38069, n685, 
        n758, n831, n904, n48321, n37308, n670, n8_adj_4467, n24_adj_4468, 
        n47823, n47821, n48310, n743, n977, n1050, n816, n889, 
        n962, n38068, n98, n37391, n29_adj_4470, n48014, n37390, 
        n4_adj_4472, n38067, n48318, n48319, n38066, n37307, n37389, 
        n47834, n38065, n47832, n48414, n48016, n48484, n48485, 
        n48460, n47825, n48434, n38064, n48022;
    wire [0:0]n9366;
    wire [21:0]n9873;
    
    wire n38208, n48436, n1035;
    wire [47:0]n106;
    
    wire n38207, n171, n244, n317, n37388, n38063, n1108, n390, 
        n463, n38062, n536, n38206, n609, n37387, n682, n755;
    wire [0:0]n8835;
    
    wire n37306, n828, n901, n974, n1047, n1120, n119, n50, 
        n192, n265_adj_4475, n338, n38061, n411, n484, n557, n630_adj_4476, 
        n95, n26_adj_4477, n83, n14_adj_4479, n168_adj_4480, n38060, 
        n38205, n241_adj_4481, n314_adj_4482, n387_adj_4483, n37386, 
        n460_adj_4484, n37385, n533_adj_4485, n156, n606_adj_4486, 
        n679_adj_4487, n752_adj_4488, n825_adj_4489, n37384;
    wire [47:0]n155;
    
    wire n37305, n38204, n38059, n898_adj_4490, n971_adj_4491, n1044_adj_4492, 
        n229, n1117_adj_4493, n92_adj_4494, n23_adj_4495, n165_adj_4496, 
        n238_adj_4497, n311_adj_4498, n384_adj_4499, n302, n38058, 
        n457_adj_4500, n530_adj_4501, n603_adj_4502, n676_adj_4503, 
        n749_adj_4504, n375, n822_adj_4505, n895_adj_4506, n968_adj_4507, 
        n1041_adj_4508, n448, n1114_adj_4509, n116_adj_4510, n47_adj_4511, 
        n189_adj_4512, n262_adj_4513, n335_adj_4514, n408_adj_4515, 
        n481_adj_4516, n521, n554_adj_4517, n627_adj_4518, n700_adj_4519, 
        n38203, n89, n20_adj_4520, n38057, n162, n594, n235, n308, 
        n381, n454_adj_4521, n38202, n38201, n527_adj_4522, n600_adj_4523, 
        n667, n673_adj_4524, n107_adj_4525, n38_adj_4526, n38056, 
        n746_adj_4527, n740, n819_adj_4528, n892_adj_4529, n813, n965_adj_4530, 
        n180_adj_4531, n1038_adj_4532, n1111_adj_4533, n86_adj_4534, 
        n17_adj_4535, n159_adj_4536, n232_adj_4537, n305_adj_4538, n378_adj_4539, 
        n38200, n451_adj_4540, n524_adj_4541, n597_adj_4542;
    wire [10:0]n18087;
    wire [9:0]n18328;
    
    wire n37891;
    wire [14:0]n16623;
    
    wire n38055, n38199, n38054, n253_adj_4543, n38198, n670_adj_4544, 
        n37890, n886, n38053, n37889, n38197, n37888, n38196, 
        n743_adj_4545, n38052, n37304, n37383, n37887, n38195, n38051, 
        n38194, n37886, n38193, n37885, n37884, n38050, n37883, 
        n816_adj_4546, n889_adj_4547, n962_adj_4548, n1035_adj_4549, 
        n1108_adj_4550, n37882, n113_adj_4551, n17_adj_4552, n9_adj_4553, 
        n11_adj_4554, n47666, n47664, n49714, n48178, n47961, n44_adj_4555, 
        n326_adj_4556, n186_adj_4557, n38192, n49696, n259_adj_4559, 
        n332_adj_4560, n47959, n399_adj_4561, n959, n405_adj_4562, 
        n478_adj_4563, n47957, n49689, n27_adj_4564, n15_adj_4565, 
        n13_adj_4566, n11_adj_4567, n47910, n21_adj_4568, n19_adj_4569, 
        n17_adj_4570, n9_adj_4571, n47917, n43_adj_4572, n16_adj_4573, 
        n47892, n8_adj_4574, n45_adj_4575, n24_adj_4576, n7_adj_4577, 
        n5_adj_4578, n47931, n48160, n48156, n25_adj_4579, n23_adj_4580, 
        n48408, n37382, n38049, n31_adj_4581, n29_adj_4582, n48258, 
        n37_adj_4583, n35_adj_4584, n33_adj_4585, n48447, n551_adj_4586, 
        n624_adj_4587, n37303, n47963, n38191, n38048, n38047, n49683, 
        n47951, n37302, n49677, n12_adj_4589, n47636, n38046, n49701, 
        n37381, n38190, n10_adj_4590, n30_adj_4591, n48272, n38189, 
        n47647, n49681, n48172, n49707, n48354, n49672, n48449, 
        n49669, n16_adj_4592, n47934, n24_adj_4593, n38188, n6_adj_4594, 
        n48374, n48375, n47624, n8_adj_4595, n49666, n48304, n48299;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3623 ;
    
    wire n3_adj_4596, n4_adj_4597, n48334, n48335, n12_adj_4598, n38045, 
        n38044, n47903, n38187, n10_adj_4599, n38043, n38042, n30_adj_4600, 
        n38041, n47906, n48410, n472_adj_4601, n47996, n37301, n697_adj_4602, 
        n770_adj_4603, n545_adj_4604, n1032, n83_adj_4605, n26_adj_4606, 
        n95_adj_4607, n48480, n48481, n14_adj_4608, n156_adj_4609;
    wire [20:0]n12116;
    
    wire n38186, n37300, n38185, n39_adj_4611, n48466, n6_adj_4612, 
        n229_adj_4613;
    wire [13:0]n17072;
    
    wire n1120_adj_4614, n38040, n1047_adj_4615, n38039, n38184, n48336, 
        n1105, n302_adj_4616, n618_adj_4617, n48337, n375_adj_4618, 
        n448_adj_4619, n47894, n38183, n48306, n47994, n41_adj_4620, 
        n47896, n974_adj_4621, n38038, n48426, n48002, n48428, n4_adj_4622, 
        n691_adj_4623, n48364, n38182, n48365, n47638, n48441, n48301, 
        n48486, n38181, n48487, n48458, n47627, n521_adj_4624, n48380, 
        n901_adj_4625, n38037, n40, n37299, n38180, n828_adj_4626, 
        n38036, n37298, n594_adj_4627, \PID_CONTROLLER.integral_23__N_3622 , 
        n755_adj_4628, n38035, n764_adj_4629, n682_adj_4630, n38034, 
        n48382, n609_adj_4631, n38033, n1099, n38179, n1026, n38178, 
        n953, n38177, n536_adj_4632, n38032, n463_adj_4633, n38031, 
        n37297, n390_adj_4635, n38030, n880, n38176, n807, n38175, 
        n317_adj_4636, n38029, n244_adj_4637, n38028, n734, n38174, 
        n171_adj_4638, n38027, n661, n38173, n37296, n29_adj_4639, 
        n98_adj_4640, n588, n38172;
    wire [12:0]n17463;
    
    wire n1050_adj_4641, n38026, n977_adj_4642, n38025, n515, n38171, 
        n37295, n667_adj_4643, n740_adj_4644, n837_adj_4645, n813_adj_4646, 
        n886_adj_4647, n910_adj_4648, n104_adj_4649, n35_adj_4650, n80, 
        n11_adj_4651, n959_adj_4652, n153_adj_4653, n177_adj_4654, n442, 
        n38170, n250_adj_4655, n323_adj_4656, n904_adj_4657, n38024;
    wire [23:0]n1_adj_4821;
    
    wire n37294, n369, n38169;
    wire [21:0]n9342;
    
    wire n37801, n37800, n37799, n37798, n37797, n37796, n37795, 
        n37794, n296, n38168, n223, n38167, n831_adj_4664, n38023, 
        n1096_adj_4665, n37793, n758_adj_4666, n38022, n1023_adj_4667, 
        n37792, n950_adj_4669, n37791, n37293, n877_adj_4671, n37790, 
        n804_adj_4672, n37789, n731_adj_4674, n37788, n658_adj_4675, 
        n37787, n685_adj_4677, n38021, n37292, n585_adj_4679, n37786, 
        n512_adj_4681, n37785, n439_adj_4682, n37784, n366_adj_4684, 
        n37783, n1032_adj_4686, n1105_adj_4687, n293_adj_4691, n37782, 
        n220_adj_4694, n37781, n147_adj_4695, n37780, n5_adj_4696, 
        n74_adj_4697;
    wire [20:0]n11631;
    
    wire n37779, n37778, n37777, n37776, n37775;
    wire [23:0]n1_adj_4822;
    
    wire n37774, n612_adj_4707, n38020, n150_adj_4708, n38166, n37773, 
        n1099_adj_4710, n37772, n1026_adj_4711, n37771, n953_adj_4719, 
        n37770, n880_adj_4720, n37769, n37291, n539_adj_4721, n38019, 
        n807_adj_4722, n37768, n734_adj_4723, n37767, n661_adj_4725, 
        n37766, n588_adj_4726, n37765, n515_adj_4727, n37764, n442_adj_4728, 
        n37763, n396_adj_4729, n369_adj_4730, n37762, n8_adj_4731, 
        n77, n37290, n466_adj_4732, n38018, n296_adj_4733, n37761, 
        n393_adj_4735, n38017;
    wire [19:0]n13367;
    
    wire n38165, n38164, n38163, n320_adj_4736, n38016, n38162, 
        n223_adj_4737, n37760, n150_adj_4740, n37759, n8_adj_4741, 
        n77_adj_4742, n247_adj_4743, n38015, n174_adj_4744, n38014, 
        n38161;
    wire [19:0]n12927;
    
    wire n37758, n38160, n1102, n38159, n1029, n38158, n37757, 
        n956, n38157, n32_adj_4749, n101_adj_4750, n37756, n37755, 
        n37754, n37289, n37753, n1102_adj_4752, n37752, n1029_adj_4753, 
        n37751, n956_adj_4754, n37750, n883, n38156, n883_adj_4755, 
        n37749, n810, n38155;
    wire [11:0]n17800;
    
    wire n980_adj_4756, n38013, n810_adj_4757, n37748, n226, n907_adj_4758, 
        n38012, n834_adj_4759, n38011, n737, n38154, n664, n38153, 
        n761_adj_4760, n38010, n591, n38152, n737_adj_4761, n37747, 
        n518, n38151, n664_adj_4762, n37746, n299, n80_adj_4764, 
        n11_adj_4765, n469_adj_4766, n542_adj_4767, n153_adj_4768, n615_adj_4769, 
        n226_adj_4770, n591_adj_4771, n37745, n518_adj_4772, n37744, 
        n445, n37743, n372, n37742, n299_adj_4773, n37741, n688_adj_4774, 
        n445_adj_4775, n38150, n372_adj_4776, n38149, n38009, n37740, 
        n38008, n37739, n38007, n38006;
    wire [18:0]n13768;
    
    wire n37738, n37737, n37736, n37735, n38148, n37734, n38147, 
        n38005, n37733, n37732, n38004, n38003, n38002, n38146, 
        n37731;
    wire [18:0]n14167;
    
    wire n38145, n38001, n37730, n37288, n37729, n38144, n38000, 
        n37728, n37727, n38143, n38142, n37999, n37726, n37725, 
        n38141, n37998, n37724, n37723, n37997, n37722, n38140, 
        n37287, n37721, n37720, n38139, n37996;
    wire [8:0]n18527;
    
    wire n37719, n37718, n37995, n37717, n37716, n37715, n37714, 
        n38138, n37994, n37713, n37712, n37711, n37993;
    wire [17:0]n14528;
    
    wire n37704, n37703, n37702, n37701, n37700, n37699, n37698, 
        n37286, n37697, n37696, n37695, n38137, n37694, n37992, 
        n37693, n37692, n37691, n37690, n37689, n37688, n37687;
    wire [16:0]n15212;
    
    wire n37686, n37685, n37684, n37683, n37682, n37991, n37681, 
        n38136, n37680, n37679, n38135, n37678, n37677, n38134, 
        n37676, n37675, n37674, n37673, n37672, n37671, n38133, 
        n37670;
    wire [7:0]n18688;
    
    wire n37669, n37668, n37667, n38132, n37285, n37666, n37665, 
        n37284, n37664, n37663, n37662;
    wire [15:0]n15824;
    
    wire n37661, n37660, n37659, n38131, n37658, n37657, n37656, 
        n37655, n38130, n37654, n37653, n37652, n37651, n37650, 
        n38129, n37649, n37648, n37647, n37646;
    wire [14:0]n16368;
    
    wire n37645, n37644, n36929;
    wire [1:0]n19072;
    
    wire n4_adj_4778, n38128, n37643, n37642, n37641, n37640, n37639, 
        n37638, n37637, n38127, n37636, n37635, n37634, n37633, 
        n37632, n37631;
    wire [6:0]n18815;
    
    wire n37630, n37629, n37628, n37627;
    wire [2:0]n19048;
    
    wire n37626, n37625, n37624;
    wire [17:0]n14888;
    
    wire n38126;
    wire [13:0]n16848;
    
    wire n37623, n37622, n37621, n37620, n38125, n37619, n37618, 
        n38124, n36970, n4_adj_4779;
    wire [3:0]n19008;
    
    wire n37617, n37616, n38123, n37615, n37614, n37613, n38122, 
        n37612, n37611, n37610, n38121, n38120, n4_adj_4781, n6_adj_4782, 
        n38119;
    wire [4:0]n18948;
    
    wire n38118, n37004;
    wire [12:0]n17268;
    
    wire n37598, n37597, n38117, n38116, n37596, n37595, n37594, 
        n37593, n37592, n37591, n37590, n38115, n37589, n37588, 
        n37587, n38114, n37586;
    wire [5:0]n18912;
    
    wire n37585, n37584, n38113, n37583, n37582, n37581, n37580, 
        n38112;
    wire [11:0]n17632;
    
    wire n37579, n37578, n37577, n37576, n37575, n38111, n37574, 
        n37573, n38110, n37572, n37571, n38109, n37570, n37569, 
        n37568, n38108, n38107;
    wire [10:0]n17944;
    
    wire n37567, n37566, n37565, n38106, n37564, n37563, n37562, 
        n37561, n37560, n38105, n37559, n37558, n37557, n38104, 
        n38103, n37556, n38102, n37555, n37554, n37553, n37552, 
        n38101, n37329, n37328, n38100;
    wire [9:0]n18208;
    
    wire n37539, n37538, n37537, n37536, n37535, n37534, n37533, 
        n37532, n37531, n37530, n37327;
    wire [8:0]n18428;
    
    wire n37529, n37528, n37527, n37326, n38099, n37526, n37525, 
        n37524, n37325, n38098, n37523, n37522, n37521, n38097;
    wire [7:0]n18608;
    
    wire n37520, n37519, n37324, n37518, n37517, n38096, n37516, 
        n37323, n37515, n37514, n37513;
    wire [6:0]n18752;
    
    wire n37512, n557_adj_4785, n37511, n484_adj_4786, n37510, n411_adj_4787, 
        n37509, n338_adj_4788, n37508, n265_adj_4789, n37507, n192_adj_4790, 
        n37506, n50_adj_4791, n119_adj_4792;
    wire [5:0]n18864;
    
    wire n560_adj_4793, n37505, n487_adj_4794, n37504, n414_adj_4795, 
        n37503, n341_adj_4796, n37502, n268_adj_4797, n37501, n195_adj_4798, 
        n37500, n53_adj_4799, n122_adj_4800, n43558, n490_adj_4801, 
        n37499, n417_adj_4802, n37498, n344_adj_4803, n37497, n271_adj_4804, 
        n37496, n198_adj_4805, n37495, n56_adj_4806, n125_adj_4807, 
        n381_adj_4808, n38095, n308_adj_4809, n38094, n235_adj_4810, 
        n38093, n37322, n162_adj_4811, n38092, n20_adj_4812, n89_adj_4813, 
        n37321, n37320, n37319, n37318, n37449, n37317, n37448, 
        n37447, n37446, n37445, n37444, n37443, n37442, n37441, 
        n37440, n37439, n37438, n37437, n37436, n37435, n37434, 
        n37433, n37432, n37431, n37430, n37429, n37428, n37427, 
        n37426, n37316, n37425, n37424, n37423, n37422, n37421, 
        n37420, n37419, n37418, n37417, n37315, n37416, n37415, 
        n37414, n37413, n37412, n37411, n37410, n37409, n37408, 
        n37407, n37406, n37405, n37314, n37404, n37403, n37402, 
        n37401, n37400, n37399, n37398, n4_adj_4814, n37072, n37047, 
        n37106, n12_adj_4815, n8_adj_4816, n11_adj_4817, n6_adj_4818, 
        n36913, n18_adj_4819, n13_adj_4820;
    
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3647[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3672[20]), .I1(n257[20]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3647[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3672[21]), .I1(n257[21]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3647[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3672[22]), .I1(n257[22]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3647[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3672[23]), .I1(n257[23]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3647[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20631_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20631_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20628_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20628_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4401));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20627_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20627_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20626_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20626_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20625_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20625_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4403));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4404));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_711_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n3616[6]), .I3(n37312), .O(\PID_CONTROLLER.integral_23__N_3572 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n37396), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n37397));
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n37395), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_711_8 (.CI(n37312), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n3616[6]), .CO(n37313));
    SB_LUT4 add_711_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n3616[5]), .I3(n37311), .O(\PID_CONTROLLER.integral_23__N_3572 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_7 (.CI(n37311), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n3616[5]), .CO(n37312));
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_17 (.CI(n37395), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n37396));
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n37394), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4406));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4407));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4409));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4410));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4412));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4413));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4414));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4415));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20624_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20624_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20623_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20623_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4416), .I1(\Kp[4] ), .I2(n19032[2]), 
            .I3(n1[18]), .O(n18983[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23943_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n19080[0]));   // verilog/motorControl.v(34[16:22])
    defparam i23943_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i20504_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_16 (.CI(n37394), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n37395));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n37393), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20649_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1514 (.I0(n4_adj_4417), .I1(\Kp[3] ), .I2(n19063[1]), 
            .I3(n1[19]), .O(n19032[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1514.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1515 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_4418));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1515.LUT_INIT = 16'h9c50;
    SB_LUT4 i24111_4_lut (.I0(n19032[2]), .I1(\Kp[4] ), .I2(n6_adj_4416), 
            .I3(n1[18]), .O(n8_adj_4419));   // verilog/motorControl.v(34[16:22])
    defparam i24111_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), .I3(n1[21]), 
            .O(n11_adj_4420));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i24072_4_lut (.I0(n19063[1]), .I1(\Kp[3] ), .I2(n4_adj_4417), 
            .I3(n1[19]), .O(n6_adj_4421));   // verilog/motorControl.v(34[16:22])
    defparam i24072_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_711_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n3616[4]), .I3(n37310), .O(\PID_CONTROLLER.integral_23__N_3572 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23945_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n36954));   // verilog/motorControl.v(34[16:22])
    defparam i23945_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4421), .I1(n11_adj_4420), .I2(n8_adj_4419), 
            .I3(n12_adj_4418), .O(n18));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), .I3(n1[22]), 
            .O(n13_adj_4422));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4422), .I1(n18), .I2(n36954), .I3(n4_adj_4423), 
            .O(n44192));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20648_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20648_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_15 (.CI(n37393), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n37394));
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_711_6 (.CI(n37310), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n3616[4]), .CO(n37311));
    SB_LUT4 add_711_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n3616[3]), .I3(n37309), .O(\PID_CONTROLLER.integral_23__N_3572 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_832_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3672[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3672[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4424));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3672[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3672[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_832_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3672[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3672[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3672[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3672[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4425));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_832_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3672[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4426));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_832_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3672[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4427));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3672[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4428));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3672[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4429));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3672[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3672[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3672[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3672[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4430));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3672[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4431));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3672[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4432));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3672[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4433));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32927_4_lut (.I0(n21_adj_4433), .I1(n19_adj_4432), .I2(n17_adj_4431), 
            .I3(n9_adj_4430), .O(n47880));
    defparam i32927_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32921_4_lut (.I0(n27), .I1(n15), .I2(n13_adj_4429), .I3(n11_adj_4428), 
            .O(n47874));
    defparam i32921_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_832_i12_3_lut (.I0(duty_23__N_3672[7]), .I1(duty_23__N_3672[16]), 
            .I2(n33), .I3(GND_net), .O(n12_adj_4434));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i10_3_lut (.I0(duty_23__N_3672[5]), .I1(duty_23__N_3672[6]), 
            .I2(n13_adj_4429), .I3(GND_net), .O(n10_adj_4435));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i30_3_lut (.I0(n12_adj_4434), .I1(duty_23__N_3672[17]), 
            .I2(n35_adj_4427), .I3(GND_net), .O(n30));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33175_4_lut (.I0(n13_adj_4429), .I1(n11_adj_4428), .I2(n9_adj_4430), 
            .I3(n47890), .O(n48128));
    defparam i33175_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33171_4_lut (.I0(n19_adj_4432), .I1(n17_adj_4431), .I2(n15), 
            .I3(n48128), .O(n48124));
    defparam i33171_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33449_4_lut (.I0(n25_adj_4426), .I1(n23_adj_4425), .I2(n21_adj_4433), 
            .I3(n48124), .O(n48402));
    defparam i33449_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33289_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n48402), 
            .O(n48242));
    defparam i33289_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33492_4_lut (.I0(n37), .I1(n35_adj_4427), .I2(n33), .I3(n48242), 
            .O(n48445));
    defparam i33492_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_832_i16_3_lut (.I0(duty_23__N_3672[9]), .I1(duty_23__N_3672[21]), 
            .I2(n43), .I3(GND_net), .O(n16));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33375_3_lut (.I0(n6_adj_4436), .I1(duty_23__N_3672[10]), .I2(n21_adj_4433), 
            .I3(GND_net), .O(n48328));   // verilog/motorControl.v(36[10:25])
    defparam i33375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33376_3_lut (.I0(n48328), .I1(duty_23__N_3672[11]), .I2(n23_adj_4425), 
            .I3(GND_net), .O(n48329));   // verilog/motorControl.v(36[10:25])
    defparam i33376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i8_3_lut (.I0(duty_23__N_3672[4]), .I1(duty_23__N_3672[8]), 
            .I2(n17_adj_4431), .I3(GND_net), .O(n8_adj_4437));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i24_3_lut (.I0(n16), .I1(duty_23__N_3672[22]), 
            .I2(n45), .I3(GND_net), .O(n24_adj_4438));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32907_4_lut (.I0(n43), .I1(n25_adj_4426), .I2(n23_adj_4425), 
            .I3(n47880), .O(n47860));
    defparam i32907_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33355_4_lut (.I0(n24_adj_4438), .I1(n8_adj_4437), .I2(n45), 
            .I3(n47858), .O(n48308));   // verilog/motorControl.v(36[10:25])
    defparam i33355_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33051_3_lut (.I0(n48329), .I1(duty_23__N_3672[12]), .I2(n25_adj_4426), 
            .I3(GND_net), .O(n48004));   // verilog/motorControl.v(36[10:25])
    defparam i33051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i4_4_lut (.I0(duty_23__N_3672[0]), .I1(duty_23__N_3672[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4439));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i33373_3_lut (.I0(n4_adj_4439), .I1(duty_23__N_3672[13]), .I2(n27), 
            .I3(GND_net), .O(n48326));   // verilog/motorControl.v(36[10:25])
    defparam i33373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33374_3_lut (.I0(n48326), .I1(duty_23__N_3672[14]), .I2(n29), 
            .I3(GND_net), .O(n48327));   // verilog/motorControl.v(36[10:25])
    defparam i33374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32917_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n47874), 
            .O(n47870));
    defparam i32917_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33459_4_lut (.I0(n30), .I1(n10_adj_4435), .I2(n35_adj_4427), 
            .I3(n47868), .O(n48412));   // verilog/motorControl.v(36[10:25])
    defparam i33459_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33053_3_lut (.I0(n48327), .I1(duty_23__N_3672[15]), .I2(n31), 
            .I3(GND_net), .O(n48006));   // verilog/motorControl.v(36[10:25])
    defparam i33053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33529_4_lut (.I0(n48006), .I1(n48412), .I2(n35_adj_4427), 
            .I3(n47870), .O(n48482));   // verilog/motorControl.v(36[10:25])
    defparam i33529_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33530_3_lut (.I0(n48482), .I1(duty_23__N_3672[18]), .I2(n37), 
            .I3(GND_net), .O(n48483));   // verilog/motorControl.v(36[10:25])
    defparam i33530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33509_3_lut (.I0(n48483), .I1(duty_23__N_3672[19]), .I2(n39), 
            .I3(GND_net), .O(n48462));   // verilog/motorControl.v(36[10:25])
    defparam i33509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32909_4_lut (.I0(n43), .I1(n41_adj_4424), .I2(n39), .I3(n48445), 
            .O(n47862));
    defparam i32909_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33477_4_lut (.I0(n48004), .I1(n48308), .I2(n45), .I3(n47860), 
            .O(n48430));   // verilog/motorControl.v(36[10:25])
    defparam i33477_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33059_3_lut (.I0(n48462), .I1(duty_23__N_3672[20]), .I2(n41_adj_4424), 
            .I3(GND_net), .O(n48012));   // verilog/motorControl.v(36[10:25])
    defparam i33059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33479_4_lut (.I0(n48012), .I1(n48430), .I2(n45), .I3(n47862), 
            .O(n48432));   // verilog/motorControl.v(36[10:25])
    defparam i33479_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33480_3_lut (.I0(n48432), .I1(PWMLimit[23]), .I2(duty_23__N_3672[23]), 
            .I3(GND_net), .O(duty_23__N_3671));   // verilog/motorControl.v(36[10:25])
    defparam i33480_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3672[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4440));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3672[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4442));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3672[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4443));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3672[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4444));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3672[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4445));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3672[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4446));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3672[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4447));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3672[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4448));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3672[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4449));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3672[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4450));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3672[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4451));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3672[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4452));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3672[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4453));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3672[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4454));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3672[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4456));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3672[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4457));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3672[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4458));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3672[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4459));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3672[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4461));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32892_4_lut (.I0(n21_adj_4461), .I1(n19_adj_4459), .I2(n17_adj_4458), 
            .I3(n9_adj_4457), .O(n47845));
    defparam i32892_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32885_4_lut (.I0(n27_adj_4456), .I1(n15_adj_4454), .I2(n13_adj_4453), 
            .I3(n11_adj_4452), .O(n47838));
    defparam i32885_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4451), 
            .I3(GND_net), .O(n12_adj_4462));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4453), 
            .I3(GND_net), .O(n10_adj_4463));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4462), .I1(n257[17]), .I2(n35_adj_4450), 
            .I3(GND_net), .O(n30_adj_4464));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n37392), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33135_4_lut (.I0(n13_adj_4453), .I1(n11_adj_4452), .I2(n9_adj_4457), 
            .I3(n47855), .O(n48088));
    defparam i33135_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_5845_18_lut (.I0(GND_net), .I1(n16112[15]), .I2(GND_net), 
            .I3(n38071), .O(n15535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5845_17_lut (.I0(GND_net), .I1(n16112[14]), .I2(GND_net), 
            .I3(n38070), .O(n15535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33129_4_lut (.I0(n19_adj_4459), .I1(n17_adj_4458), .I2(n15_adj_4454), 
            .I3(n48088), .O(n48082));
    defparam i33129_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33443_4_lut (.I0(n25_adj_4449), .I1(n23_adj_4448), .I2(n21_adj_4461), 
            .I3(n48082), .O(n48396));
    defparam i33443_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33271_4_lut (.I0(n31_adj_4447), .I1(n29_adj_4446), .I2(n27_adj_4456), 
            .I3(n48396), .O(n48224));
    defparam i33271_4_lut.LUT_INIT = 16'hfeff;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3548[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_711_5 (.CI(n37309), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n3616[3]), .CO(n37310));
    SB_LUT4 i33490_4_lut (.I0(n37_adj_4445), .I1(n35_adj_4450), .I2(n33_adj_4451), 
            .I3(n48224), .O(n48443));
    defparam i33490_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4444), 
            .I3(GND_net), .O(n16_adj_4465));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5845_17 (.CI(n38070), .I0(n16112[14]), .I1(GND_net), 
            .CO(n38071));
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33367_3_lut (.I0(n6_adj_4466), .I1(n257[10]), .I2(n21_adj_4461), 
            .I3(GND_net), .O(n48320));   // verilog/motorControl.v(38[19:35])
    defparam i33367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5845_16_lut (.I0(GND_net), .I1(n16112[13]), .I2(n1114), 
            .I3(n38069), .O(n15535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33368_3_lut (.I0(n48320), .I1(n257[11]), .I2(n23_adj_4448), 
            .I3(GND_net), .O(n48321));   // verilog/motorControl.v(38[19:35])
    defparam i33368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_711_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n3616[2]), .I3(n37308), .O(\PID_CONTROLLER.integral_23__N_3572 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n37392), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n37393));
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4458), 
            .I3(GND_net), .O(n8_adj_4467));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4465), .I1(n257[22]), .I2(n45_adj_4443), 
            .I3(GND_net), .O(n24_adj_4468));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32870_4_lut (.I0(n43_adj_4444), .I1(n25_adj_4449), .I2(n23_adj_4448), 
            .I3(n47845), .O(n47823));
    defparam i32870_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33357_4_lut (.I0(n24_adj_4468), .I1(n8_adj_4467), .I2(n45_adj_4443), 
            .I3(n47821), .O(n48310));   // verilog/motorControl.v(38[19:35])
    defparam i33357_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5845_16 (.CI(n38069), .I0(n16112[13]), .I1(n1114), .CO(n38070));
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_711_4 (.CI(n37308), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n3616[2]), .CO(n37309));
    SB_LUT4 add_5845_15_lut (.I0(GND_net), .I1(n16112[12]), .I2(n1041), 
            .I3(n38068), .O(n15535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n37391), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4470));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33061_3_lut (.I0(n48321), .I1(n257[12]), .I2(n25_adj_4449), 
            .I3(GND_net), .O(n48014));   // verilog/motorControl.v(38[19:35])
    defparam i33061_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_13 (.CI(n37391), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n37392));
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n37390), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5845_15 (.CI(n38068), .I0(n16112[12]), .I1(n1041), .CO(n38069));
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3672[0]), .I1(n257[1]), 
            .I2(duty_23__N_3672[1]), .I3(n257[0]), .O(n4_adj_4472));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_5845_14_lut (.I0(GND_net), .I1(n16112[11]), .I2(n968), 
            .I3(n38067), .O(n15535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33365_3_lut (.I0(n4_adj_4472), .I1(n257[13]), .I2(n27_adj_4456), 
            .I3(GND_net), .O(n48318));   // verilog/motorControl.v(38[19:35])
    defparam i33365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33366_3_lut (.I0(n48318), .I1(n257[14]), .I2(n29_adj_4446), 
            .I3(GND_net), .O(n48319));   // verilog/motorControl.v(38[19:35])
    defparam i33366_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_12 (.CI(n37390), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n37391));
    SB_CARRY add_5845_14 (.CI(n38067), .I0(n16112[11]), .I1(n968), .CO(n38068));
    SB_LUT4 add_5845_13_lut (.I0(GND_net), .I1(n16112[10]), .I2(n895), 
            .I3(n38066), .O(n15535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5845_13 (.CI(n38066), .I0(n16112[10]), .I1(n895), .CO(n38067));
    SB_LUT4 add_711_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3616[1]), .I3(n37307), .O(\PID_CONTROLLER.integral_23__N_3572 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n37389), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32881_4_lut (.I0(n33_adj_4451), .I1(n31_adj_4447), .I2(n29_adj_4446), 
            .I3(n47838), .O(n47834));
    defparam i32881_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5845_12_lut (.I0(GND_net), .I1(n16112[9]), .I2(n822), 
            .I3(n38065), .O(n15535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_3 (.CI(n37307), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n3616[1]), .CO(n37308));
    SB_CARRY add_5845_12 (.CI(n38065), .I0(n16112[9]), .I1(n822), .CO(n38066));
    SB_LUT4 i33461_4_lut (.I0(n30_adj_4464), .I1(n10_adj_4463), .I2(n35_adj_4450), 
            .I3(n47832), .O(n48414));   // verilog/motorControl.v(38[19:35])
    defparam i33461_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY sub_3_add_2_11 (.CI(n37389), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n37390));
    SB_LUT4 i33063_3_lut (.I0(n48319), .I1(n257[15]), .I2(n31_adj_4447), 
            .I3(GND_net), .O(n48016));   // verilog/motorControl.v(38[19:35])
    defparam i33063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33531_4_lut (.I0(n48016), .I1(n48414), .I2(n35_adj_4450), 
            .I3(n47834), .O(n48484));   // verilog/motorControl.v(38[19:35])
    defparam i33531_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33532_3_lut (.I0(n48484), .I1(n257[18]), .I2(n37_adj_4445), 
            .I3(GND_net), .O(n48485));   // verilog/motorControl.v(38[19:35])
    defparam i33532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33507_3_lut (.I0(n48485), .I1(n257[19]), .I2(n39_adj_4442), 
            .I3(GND_net), .O(n48460));   // verilog/motorControl.v(38[19:35])
    defparam i33507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32872_4_lut (.I0(n43_adj_4444), .I1(n41_adj_4440), .I2(n39_adj_4442), 
            .I3(n48443), .O(n47825));
    defparam i32872_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_711_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n3616[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3572 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33481_4_lut (.I0(n48014), .I1(n48310), .I2(n45_adj_4443), 
            .I3(n47823), .O(n48434));   // verilog/motorControl.v(38[19:35])
    defparam i33481_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5845_11_lut (.I0(GND_net), .I1(n16112[8]), .I2(n749), 
            .I3(n38064), .O(n15535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33069_3_lut (.I0(n48460), .I1(n257[20]), .I2(n41_adj_4440), 
            .I3(GND_net), .O(n48022));   // verilog/motorControl.v(38[19:35])
    defparam i33069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n9873[21]), .I2(GND_net), 
            .I3(n38208), .O(n9366[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33483_4_lut (.I0(n48022), .I1(n48434), .I2(n45_adj_4443), 
            .I3(n47825), .O(n48436));   // verilog/motorControl.v(38[19:35])
    defparam i33483_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33484_3_lut (.I0(n48436), .I1(duty_23__N_3672[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(38[19:35])
    defparam i33484_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3672[0]), .I1(n257[0]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3647[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n9873[20]), .I2(GND_net), 
            .I3(n38207), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5845_11 (.CI(n38064), .I0(n16112[8]), .I1(n749), .CO(n38065));
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n37388), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5845_10_lut (.I0(GND_net), .I1(n16112[7]), .I2(n676), 
            .I3(n38063), .O(n15535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_23 (.CI(n38207), .I0(n9873[20]), .I1(GND_net), 
            .CO(n38208));
    SB_CARRY add_5845_10 (.CI(n38063), .I0(n16112[7]), .I1(n676), .CO(n38064));
    SB_CARRY add_711_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n3616[0]), .CO(n37307));
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5845_9_lut (.I0(GND_net), .I1(n16112[6]), .I2(n603), .I3(n38062), 
            .O(n15535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5845_9 (.CI(n38062), .I0(n16112[6]), .I1(n603), .CO(n38063));
    SB_CARRY sub_3_add_2_10 (.CI(n37388), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n37389));
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n9873[19]), .I2(GND_net), 
            .I3(n38206), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n37387), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n9366[0]), .I2(n8835[0]), 
            .I3(n37306), .O(duty_23__N_3672[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5845_8_lut (.I0(GND_net), .I1(n16112[5]), .I2(n530), .I3(n38061), 
            .O(n15535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_22 (.CI(n38206), .I0(n9873[19]), .I1(GND_net), 
            .CO(n38207));
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5845_8 (.CI(n38061), .I0(n16112[5]), .I1(n530), .CO(n38062));
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4476));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4477));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4479));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4480));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_9 (.CI(n37387), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n37388));
    SB_LUT4 add_5845_7_lut (.I0(GND_net), .I1(n16112[4]), .I2(n457), .I3(n38060), 
            .O(n15535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n9873[18]), .I2(GND_net), 
            .I3(n38205), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4482));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4483));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n37386), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_8 (.CI(n37386), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n37387));
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n37385), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5845_7 (.CI(n38060), .I0(n16112[4]), .I1(n457), .CO(n38061));
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4485));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4486));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_7 (.CI(n37385), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n37386));
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4488));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4489));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n37384), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n37305), .O(duty_23__N_3672[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n38205), .I0(n9873[18]), .I1(GND_net), 
            .CO(n38206));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n9873[17]), .I2(GND_net), 
            .I3(n38204), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5845_6_lut (.I0(GND_net), .I1(n16112[3]), .I2(n384), .I3(n38059), 
            .O(n15535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4491));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_20 (.CI(n38204), .I0(n9873[17]), .I1(GND_net), 
            .CO(n38205));
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4492));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4493));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4494));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4495));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4496));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5845_6 (.CI(n38059), .I0(n16112[3]), .I1(n384), .CO(n38060));
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4497));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4498));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4499));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_24 (.CI(n37305), .I0(n106[22]), .I1(n155[22]), .CO(n37306));
    SB_LUT4 add_5845_5_lut (.I0(GND_net), .I1(n16112[2]), .I2(n311), .I3(n38058), 
            .O(n15535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4500));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4501));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4502));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4503));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4504));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4505));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4506));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4507));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4508));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4509));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4510));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4511));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4513));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4514));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4516));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4517));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4519));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n9873[16]), .I2(GND_net), 
            .I3(n38203), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_19 (.CI(n38203), .I0(n9873[16]), .I1(GND_net), 
            .CO(n38204));
    SB_CARRY add_5845_5 (.CI(n38058), .I0(n16112[2]), .I1(n311), .CO(n38059));
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4520));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5845_4_lut (.I0(GND_net), .I1(n16112[1]), .I2(n238), .I3(n38057), 
            .O(n15535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20647_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n9873[15]), .I2(GND_net), 
            .I3(n38202), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n38202), .I0(n9873[15]), .I1(GND_net), 
            .CO(n38203));
    SB_CARRY add_5845_4 (.CI(n38057), .I0(n16112[1]), .I1(n238), .CO(n38058));
    SB_LUT4 i20646_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20646_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n9873[14]), .I2(GND_net), 
            .I3(n38201), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4522));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4523));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4525));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4526));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5845_3_lut (.I0(GND_net), .I1(n16112[0]), .I2(n165), .I3(n38056), 
            .O(n15535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5845_3 (.CI(n38056), .I0(n16112[0]), .I1(n165), .CO(n38057));
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4528));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4529));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4531));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4532));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4534));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4535));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5845_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n15535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5845_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4537));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_17 (.CI(n38201), .I0(n9873[14]), .I1(GND_net), 
            .CO(n38202));
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4538));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n9873[13]), .I2(n1096), 
            .I3(n38200), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4540));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20645_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4541));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5845_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n38056));
    SB_CARRY mult_10_add_1225_16 (.CI(n38200), .I0(n9873[13]), .I1(n1096), 
            .CO(n38201));
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6007_12_lut (.I0(GND_net), .I1(n18328[9]), .I2(n840), 
            .I3(n37891), .O(n18087[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5877_17_lut (.I0(GND_net), .I1(n16623[14]), .I2(GND_net), 
            .I3(n38055), .O(n16112[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n9873[12]), .I2(n1023), 
            .I3(n38199), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n38199), .I0(n9873[12]), .I1(n1023), 
            .CO(n38200));
    SB_LUT4 add_5877_16_lut (.I0(GND_net), .I1(n16623[13]), .I2(n1117), 
            .I3(n38054), .O(n16112[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_16 (.CI(n38054), .I0(n16623[13]), .I1(n1117), .CO(n38055));
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4543));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n9873[11]), .I2(n950), 
            .I3(n38198), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n38198), .I0(n9873[11]), .I1(n950), 
            .CO(n38199));
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4544));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6007_11_lut (.I0(GND_net), .I1(n18328[8]), .I2(n767), 
            .I3(n37890), .O(n18087[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_11 (.CI(n37890), .I0(n18328[8]), .I1(n767), .CO(n37891));
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5877_15_lut (.I0(GND_net), .I1(n16623[12]), .I2(n1044), 
            .I3(n38053), .O(n16112[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6007_10_lut (.I0(GND_net), .I1(n18328[7]), .I2(n694), 
            .I3(n37889), .O(n18087[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_10 (.CI(n37889), .I0(n18328[7]), .I1(n694), .CO(n37890));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n9873[10]), .I2(n877), 
            .I3(n38197), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6007_9_lut (.I0(GND_net), .I1(n18328[6]), .I2(n621), .I3(n37888), 
            .O(n18087[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n37384), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n37385));
    SB_CARRY mult_10_add_1225_13 (.CI(n38197), .I0(n9873[10]), .I1(n877), 
            .CO(n38198));
    SB_CARRY add_6007_9 (.CI(n37888), .I0(n18328[6]), .I1(n621), .CO(n37889));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n9873[9]), .I2(n804), 
            .I3(n38196), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_12 (.CI(n38196), .I0(n9873[9]), .I1(n804), 
            .CO(n38197));
    SB_CARRY add_5877_15 (.CI(n38053), .I0(n16623[12]), .I1(n1044), .CO(n38054));
    SB_LUT4 add_5877_14_lut (.I0(GND_net), .I1(n16623[11]), .I2(n971), 
            .I3(n38052), .O(n16112[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n37304), .O(duty_23__N_3672[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n37383), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6007_8_lut (.I0(GND_net), .I1(n18328[5]), .I2(n548), .I3(n37887), 
            .O(n18087[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n9873[8]), .I2(n731), 
            .I3(n38195), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_5 (.CI(n37383), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n37384));
    SB_CARRY add_5877_14 (.CI(n38052), .I0(n16623[11]), .I1(n971), .CO(n38053));
    SB_LUT4 add_5877_13_lut (.I0(GND_net), .I1(n16623[10]), .I2(n898), 
            .I3(n38051), .O(n16112[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n38195), .I0(n9873[8]), .I1(n731), 
            .CO(n38196));
    SB_CARRY add_6007_8 (.CI(n37887), .I0(n18328[5]), .I1(n548), .CO(n37888));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n9873[7]), .I2(n658), 
            .I3(n38194), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n38194), .I0(n9873[7]), .I1(n658), 
            .CO(n38195));
    SB_LUT4 add_6007_7_lut (.I0(GND_net), .I1(n18328[4]), .I2(n475), .I3(n37886), 
            .O(n18087[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_13 (.CI(n38051), .I0(n16623[10]), .I1(n898), .CO(n38052));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n9873[6]), .I2(n585), 
            .I3(n38193), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_7 (.CI(n37886), .I0(n18328[4]), .I1(n475), .CO(n37887));
    SB_LUT4 add_6007_6_lut (.I0(GND_net), .I1(n18328[3]), .I2(n402), .I3(n37885), 
            .O(n18087[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_6 (.CI(n37885), .I0(n18328[3]), .I1(n402), .CO(n37886));
    SB_LUT4 add_6007_5_lut (.I0(GND_net), .I1(n18328[2]), .I2(n329), .I3(n37884), 
            .O(n18087[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_5 (.CI(n37884), .I0(n18328[2]), .I1(n329), .CO(n37885));
    SB_LUT4 i20641_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5877_12_lut (.I0(GND_net), .I1(n16623[9]), .I2(n825), 
            .I3(n38050), .O(n16112[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6007_4_lut (.I0(GND_net), .I1(n18328[1]), .I2(n256_adj_4405), 
            .I3(n37883), .O(n18087[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_4 (.CI(n37883), .I0(n18328[1]), .I1(n256_adj_4405), 
            .CO(n37884));
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4546));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4547));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4549));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4550));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6007_3_lut (.I0(GND_net), .I1(n18328[0]), .I2(n183), .I3(n37882), 
            .O(n18087[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_3 (.CI(n37882), .I0(n18328[0]), .I1(n183), .CO(n37883));
    SB_LUT4 add_6007_2_lut (.I0(GND_net), .I1(n41_adj_4404), .I2(n110_adj_4403), 
            .I3(GND_net), .O(n18087[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6007_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6007_2 (.CI(GND_net), .I0(n41_adj_4404), .I1(n110_adj_4403), 
            .CO(n37882));
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4552));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_9 (.CI(n38193), .I0(n9873[6]), .I1(n585), 
            .CO(n38194));
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4553));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4554));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5877_12 (.CI(n38050), .I0(n16623[9]), .I1(n825), .CO(n38051));
    SB_LUT4 i32713_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n47666));
    defparam i32713_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i32711_3_lut (.I0(n11_adj_4554), .I1(n9_adj_4553), .I2(n47666), 
            .I3(GND_net), .O(n47664));
    defparam i32711_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_172_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n49714));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_172_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33225_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n49714), 
            .I2(IntegralLimit[7]), .I3(n47664), .O(n48178));
    defparam i33225_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i33008_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4552), 
            .I2(IntegralLimit[9]), .I3(n48178), .O(n47961));
    defparam i33008_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4555));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4556));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n9873[5]), .I2(n512), 
            .I3(n38192), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_154_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n49696));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_154_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4559));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33006_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4552), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4553), .O(n47959));
    defparam i33006_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4561));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4562));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4563));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33004_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n49696), 
            .I2(IntegralLimit[11]), .I3(n47959), .O(n47957));
    defparam i33004_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_147_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n49689));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_147_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32957_4_lut (.I0(n27_adj_4564), .I1(n15_adj_4565), .I2(n13_adj_4566), 
            .I3(n11_adj_4567), .O(n47910));
    defparam i32957_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32964_4_lut (.I0(n21_adj_4568), .I1(n19_adj_4569), .I2(n17_adj_4570), 
            .I3(n9_adj_4571), .O(n47917));
    defparam i32964_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_4572), .I3(GND_net), 
            .O(n16_adj_4573));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i32939_2_lut (.I0(n43_adj_4572), .I1(n19_adj_4569), .I2(GND_net), 
            .I3(GND_net), .O(n47892));
    defparam i32939_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4570), .I3(GND_net), 
            .O(n8_adj_4574));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4573), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_4575), .I3(GND_net), 
            .O(n24_adj_4576));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i32978_2_lut (.I0(n7_adj_4577), .I1(n5_adj_4578), .I2(GND_net), 
            .I3(GND_net), .O(n47931));
    defparam i32978_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33207_4_lut (.I0(n13_adj_4566), .I1(n11_adj_4567), .I2(n9_adj_4571), 
            .I3(n47931), .O(n48160));
    defparam i33207_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY mult_10_add_1225_8 (.CI(n38192), .I0(n9873[5]), .I1(n512), 
            .CO(n38193));
    SB_LUT4 i33203_4_lut (.I0(n19_adj_4569), .I1(n17_adj_4570), .I2(n15_adj_4565), 
            .I3(n48160), .O(n48156));
    defparam i33203_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33455_4_lut (.I0(n25_adj_4579), .I1(n23_adj_4580), .I2(n21_adj_4568), 
            .I3(n48156), .O(n48408));
    defparam i33455_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_12_23 (.CI(n37304), .I0(n106[21]), .I1(n155[21]), .CO(n37305));
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n37382), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5877_11_lut (.I0(GND_net), .I1(n16623[8]), .I2(n752), 
            .I3(n38049), .O(n16112[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33305_4_lut (.I0(n31_adj_4581), .I1(n29_adj_4582), .I2(n27_adj_4564), 
            .I3(n48408), .O(n48258));
    defparam i33305_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33494_4_lut (.I0(n37_adj_4583), .I1(n35_adj_4584), .I2(n33_adj_4585), 
            .I3(n48258), .O(n48447));
    defparam i33494_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4586));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4587));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5877_11 (.CI(n38049), .I0(n16623[8]), .I1(n752), .CO(n38050));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n37303), .O(duty_23__N_3672[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33010_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n49714), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4554), .O(n47963));
    defparam i33010_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n9873[4]), .I2(n439), 
            .I3(n38191), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n38191), .I0(n9873[4]), .I1(n439), 
            .CO(n38192));
    SB_LUT4 add_5877_10_lut (.I0(GND_net), .I1(n16623[7]), .I2(n679), 
            .I3(n38048), .O(n16112[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_10 (.CI(n38048), .I0(n16623[7]), .I1(n679), .CO(n38049));
    SB_LUT4 add_5877_9_lut (.I0(GND_net), .I1(n16623[6]), .I2(n606), .I3(n38047), 
            .O(n16112[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_141_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n49683));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_141_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_22 (.CI(n37303), .I0(n106[20]), .I1(n155[20]), .CO(n37304));
    SB_LUT4 i32998_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n49683), 
            .I2(IntegralLimit[14]), .I3(n47963), .O(n47951));
    defparam i32998_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n37302), .O(duty_23__N_3672[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_135_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n49677));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_135_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4589));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32683_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n47636));
    defparam i32683_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_5877_9 (.CI(n38047), .I0(n16623[6]), .I1(n606), .CO(n38048));
    SB_LUT4 add_5877_8_lut (.I0(GND_net), .I1(n16623[5]), .I2(n533), .I3(n38046), 
            .O(n16112[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_159_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n49701));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_159_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_3_add_2_4 (.CI(n37382), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n37383));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n37381), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n9873[3]), .I2(n366), 
            .I3(n38190), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n38190), .I0(n9873[3]), .I1(n366), 
            .CO(n38191));
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4590));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4589), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_4591));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33319_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n49696), 
            .I2(IntegralLimit[11]), .I3(n47961), .O(n48272));
    defparam i33319_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n9873[2]), .I2(n293), 
            .I3(n38189), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32694_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n49689), 
            .I2(IntegralLimit[13]), .I3(n48272), .O(n47647));
    defparam i32694_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_139_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n49681));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_139_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33219_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n49681), 
            .I2(IntegralLimit[15]), .I3(n47647), .O(n48172));
    defparam i33219_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_165_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n49707));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_165_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33401_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n49707), 
            .I2(IntegralLimit[17]), .I3(n48172), .O(n48354));
    defparam i33401_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_130_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n49672));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_130_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33496_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n49672), 
            .I2(IntegralLimit[19]), .I3(n48354), .O(n48449));
    defparam i33496_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_127_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n49669));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_127_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4592));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32981_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n47934));
    defparam i32981_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY mult_10_add_1225_5 (.CI(n38189), .I0(n9873[2]), .I1(n293), 
            .CO(n38190));
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4592), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4593));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n9873[1]), .I2(n220), 
            .I3(n38188), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4594));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5877_8 (.CI(n38046), .I0(n16623[5]), .I1(n533), .CO(n38047));
    SB_LUT4 i33421_3_lut (.I0(n6_adj_4594), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n48374));   // verilog/motorControl.v(31[10:34])
    defparam i33421_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33422_3_lut (.I0(n48374), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n48375));   // verilog/motorControl.v(31[10:34])
    defparam i33422_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_3_add_2_3 (.CI(n37381), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n37382));
    SB_LUT4 i32671_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n49689), 
            .I2(IntegralLimit[21]), .I3(n47957), .O(n47624));
    defparam i32671_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i33351_4_lut (.I0(n24_adj_4593), .I1(n8_adj_4595), .I2(n49666), 
            .I3(n47934), .O(n48304));   // verilog/motorControl.v(31[10:34])
    defparam i33351_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33346_3_lut (.I0(n48375), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n48299));   // verilog/motorControl.v(31[10:34])
    defparam i33346_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3623 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4596), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4597));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i33381_3_lut (.I0(n4_adj_4597), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27_adj_4564), .I3(GND_net), .O(n48334));   // verilog/motorControl.v(31[38:63])
    defparam i33381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33382_3_lut (.I0(n48334), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4582), .I3(GND_net), .O(n48335));   // verilog/motorControl.v(31[38:63])
    defparam i33382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33_adj_4585), .I3(GND_net), 
            .O(n12_adj_4598));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_5877_7_lut (.I0(GND_net), .I1(n16623[4]), .I2(n460), .I3(n38045), 
            .O(n16112[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_7 (.CI(n38045), .I0(n16623[4]), .I1(n460), .CO(n38046));
    SB_CARRY mult_10_add_1225_4 (.CI(n38188), .I0(n9873[1]), .I1(n220), 
            .CO(n38189));
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5877_6_lut (.I0(GND_net), .I1(n16623[3]), .I2(n387), .I3(n38044), 
            .O(n16112[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32950_2_lut (.I0(n33_adj_4585), .I1(n15_adj_4565), .I2(GND_net), 
            .I3(GND_net), .O(n47903));
    defparam i32950_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n9873[0]), .I2(n147), 
            .I3(n38187), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_6 (.CI(n38044), .I0(n16623[3]), .I1(n387), .CO(n38045));
    SB_CARRY mult_10_add_1225_3 (.CI(n38187), .I0(n9873[0]), .I1(n147), 
            .CO(n38188));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4566), .I3(GND_net), 
            .O(n10_adj_4599));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_5877_5_lut (.I0(GND_net), .I1(n16623[2]), .I2(n314), .I3(n38043), 
            .O(n16112[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_5 (.CI(n38043), .I0(n16623[2]), .I1(n314), .CO(n38044));
    SB_LUT4 add_5877_4_lut (.I0(GND_net), .I1(n16623[1]), .I2(n241), .I3(n38042), 
            .O(n16112[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_4 (.CI(n38042), .I0(n16623[1]), .I1(n241), .CO(n38043));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4598), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4584), .I3(GND_net), 
            .O(n30_adj_4600));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_5877_3_lut (.I0(GND_net), .I1(n16623[0]), .I2(n168), .I3(n38041), 
            .O(n16112[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32953_4_lut (.I0(n33_adj_4585), .I1(n31_adj_4581), .I2(n29_adj_4582), 
            .I3(n47910), .O(n47906));
    defparam i32953_4_lut.LUT_INIT = 16'haaab;
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_12_21 (.CI(n37302), .I0(n106[19]), .I1(n155[19]), .CO(n37303));
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5877_3 (.CI(n38041), .I0(n16623[0]), .I1(n168), .CO(n38042));
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n38187));
    SB_LUT4 i33457_4_lut (.I0(n30_adj_4600), .I1(n10_adj_4599), .I2(n35_adj_4584), 
            .I3(n47903), .O(n48410));   // verilog/motorControl.v(31[38:63])
    defparam i33457_4_lut.LUT_INIT = 16'haaac;
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n37381));
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3548[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3548[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3548[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3548[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3548[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3548[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3548[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3548[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3548[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4601));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33043_3_lut (.I0(n48335), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_4581), .I3(GND_net), .O(n47996));   // verilog/motorControl.v(31[38:63])
    defparam i33043_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3548[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3548[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3548[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3548[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n37301), .O(duty_23__N_3672[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3548[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3548[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3548[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3548[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4602));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3548[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3548[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3548[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3548[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3548[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3548[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4604));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4605));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_20 (.CI(n37301), .I0(n106[18]), .I1(n155[18]), .CO(n37302));
    SB_LUT4 add_5877_2_lut (.I0(GND_net), .I1(n26_adj_4606), .I2(n95_adj_4607), 
            .I3(GND_net), .O(n16112[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5877_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33527_4_lut (.I0(n47996), .I1(n48410), .I2(n35_adj_4584), 
            .I3(n47906), .O(n48480));   // verilog/motorControl.v(31[38:63])
    defparam i33527_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33528_3_lut (.I0(n48480), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37_adj_4583), .I3(GND_net), .O(n48481));   // verilog/motorControl.v(31[38:63])
    defparam i33528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4608));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4081_23_lut (.I0(GND_net), .I1(n12116[20]), .I2(GND_net), 
            .I3(n38186), .O(n9873[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n37300), .O(duty_23__N_3672[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4081_22_lut (.I0(GND_net), .I1(n12116[19]), .I2(GND_net), 
            .I3(n38185), .O(n9873[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5877_2 (.CI(GND_net), .I0(n26_adj_4606), .I1(n95_adj_4607), 
            .CO(n38041));
    SB_LUT4 i33513_3_lut (.I0(n48481), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_4611), .I3(GND_net), .O(n48466));   // verilog/motorControl.v(31[38:63])
    defparam i33513_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_12_19 (.CI(n37300), .I0(n106[17]), .I1(n155[17]), .CO(n37301));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4577), .I3(GND_net), 
            .O(n6_adj_4612));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4613));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5907_16_lut (.I0(GND_net), .I1(n17072[13]), .I2(n1120_adj_4614), 
            .I3(n38040), .O(n16623[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5907_15_lut (.I0(GND_net), .I1(n17072[12]), .I2(n1047_adj_4615), 
            .I3(n38039), .O(n16623[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_22 (.CI(n38185), .I0(n12116[19]), .I1(GND_net), 
            .CO(n38186));
    SB_LUT4 add_4081_21_lut (.I0(GND_net), .I1(n12116[18]), .I2(GND_net), 
            .I3(n38184), .O(n9873[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33383_3_lut (.I0(n6_adj_4612), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4568), .I3(GND_net), .O(n48336));   // verilog/motorControl.v(31[38:63])
    defparam i33383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4616));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4617));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33384_3_lut (.I0(n48336), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4580), .I3(GND_net), .O(n48337));   // verilog/motorControl.v(31[38:63])
    defparam i33384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4619));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32941_4_lut (.I0(n43_adj_4572), .I1(n25_adj_4579), .I2(n23_adj_4580), 
            .I3(n47917), .O(n47894));
    defparam i32941_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4081_21 (.CI(n38184), .I0(n12116[18]), .I1(GND_net), 
            .CO(n38185));
    SB_CARRY add_5907_15 (.CI(n38039), .I0(n17072[12]), .I1(n1047_adj_4615), 
            .CO(n38040));
    SB_LUT4 add_4081_20_lut (.I0(GND_net), .I1(n12116[17]), .I2(GND_net), 
            .I3(n38183), .O(n9873[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33353_4_lut (.I0(n24_adj_4576), .I1(n8_adj_4574), .I2(n45_adj_4575), 
            .I3(n47892), .O(n48306));   // verilog/motorControl.v(31[38:63])
    defparam i33353_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4081_20 (.CI(n38183), .I0(n12116[17]), .I1(GND_net), 
            .CO(n38184));
    SB_LUT4 i33041_3_lut (.I0(n48337), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4579), .I3(GND_net), .O(n47994));   // verilog/motorControl.v(31[38:63])
    defparam i33041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32943_4_lut (.I0(n43_adj_4572), .I1(n41_adj_4620), .I2(n39_adj_4611), 
            .I3(n48447), .O(n47896));
    defparam i32943_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5907_14_lut (.I0(GND_net), .I1(n17072[11]), .I2(n974_adj_4621), 
            .I3(n38038), .O(n16623[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33473_4_lut (.I0(n47994), .I1(n48306), .I2(n45_adj_4575), 
            .I3(n47894), .O(n48426));   // verilog/motorControl.v(31[38:63])
    defparam i33473_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33049_3_lut (.I0(n48466), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4620), .I3(GND_net), .O(n48002));   // verilog/motorControl.v(31[38:63])
    defparam i33049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33475_4_lut (.I0(n48002), .I1(n48426), .I2(n45_adj_4575), 
            .I3(n47896), .O(n48428));   // verilog/motorControl.v(31[38:63])
    defparam i33475_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4622));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4623));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5907_14 (.CI(n38038), .I0(n17072[11]), .I1(n974_adj_4621), 
            .CO(n38039));
    SB_LUT4 i33411_3_lut (.I0(n4_adj_4622), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n48364));   // verilog/motorControl.v(31[10:34])
    defparam i33411_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4081_19_lut (.I0(GND_net), .I1(n12116[16]), .I2(GND_net), 
            .I3(n38182), .O(n9873[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33412_3_lut (.I0(n48364), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n48365));   // verilog/motorControl.v(31[10:34])
    defparam i33412_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32685_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n49677), 
            .I2(IntegralLimit[16]), .I3(n47951), .O(n47638));
    defparam i32685_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_4081_19 (.CI(n38182), .I0(n12116[16]), .I1(GND_net), 
            .CO(n38183));
    SB_LUT4 i33488_4_lut (.I0(n30_adj_4591), .I1(n10_adj_4590), .I2(n49701), 
            .I3(n47636), .O(n48441));   // verilog/motorControl.v(31[10:34])
    defparam i33488_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33348_3_lut (.I0(n48365), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n48301));   // verilog/motorControl.v(31[10:34])
    defparam i33348_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33533_4_lut (.I0(n48301), .I1(n48441), .I2(n49701), .I3(n47638), 
            .O(n48486));   // verilog/motorControl.v(31[10:34])
    defparam i33533_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4081_18_lut (.I0(GND_net), .I1(n12116[15]), .I2(GND_net), 
            .I3(n38181), .O(n9873[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33534_3_lut (.I0(n48486), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n48487));   // verilog/motorControl.v(31[10:34])
    defparam i33534_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33505_3_lut (.I0(n48487), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n48458));   // verilog/motorControl.v(31[10:34])
    defparam i33505_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32674_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n49669), 
            .I2(IntegralLimit[21]), .I3(n48449), .O(n47627));
    defparam i32674_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_124_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n49666));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_124_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33427_4_lut (.I0(n48299), .I1(n48304), .I2(n49666), .I3(n47624), 
            .O(n48380));   // verilog/motorControl.v(31[10:34])
    defparam i33427_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5907_13_lut (.I0(GND_net), .I1(n17072[10]), .I2(n901_adj_4625), 
            .I3(n38037), .O(n16623[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33503_3_lut (.I0(n48458), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[10:34])
    defparam i33503_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n37299), .O(duty_23__N_3672[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_18 (.CI(n37299), .I0(n106[16]), .I1(n155[16]), .CO(n37300));
    SB_CARRY add_4081_18 (.CI(n38181), .I0(n12116[15]), .I1(GND_net), 
            .CO(n38182));
    SB_CARRY add_5907_13 (.CI(n38037), .I0(n17072[10]), .I1(n901_adj_4625), 
            .CO(n38038));
    SB_LUT4 add_4081_17_lut (.I0(GND_net), .I1(n12116[14]), .I2(GND_net), 
            .I3(n38180), .O(n9873[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5907_12_lut (.I0(GND_net), .I1(n17072[9]), .I2(n828_adj_4626), 
            .I3(n38036), .O(n16623[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n37298), .O(duty_23__N_3672[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5907_12 (.CI(n38036), .I0(n17072[9]), .I1(n828_adj_4626), 
            .CO(n38037));
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33476_3_lut (.I0(n48428), .I1(\PID_CONTROLLER.integral_23__N_3623 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3622 ));   // verilog/motorControl.v(31[38:63])
    defparam i33476_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5907_11_lut (.I0(GND_net), .I1(n17072[8]), .I2(n755_adj_4628), 
            .I3(n38035), .O(n16623[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5907_11 (.CI(n38035), .I0(n17072[8]), .I1(n755_adj_4628), 
            .CO(n38036));
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4629));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5907_10_lut (.I0(GND_net), .I1(n17072[7]), .I2(n682_adj_4630), 
            .I3(n38034), .O(n16623[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33429_4_lut (.I0(n40), .I1(n48380), .I2(n49666), .I3(n47627), 
            .O(n48382));   // verilog/motorControl.v(31[10:34])
    defparam i33429_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5907_10 (.CI(n38034), .I0(n17072[7]), .I1(n682_adj_4630), 
            .CO(n38035));
    SB_LUT4 add_5907_9_lut (.I0(GND_net), .I1(n17072[6]), .I2(n609_adj_4631), 
            .I3(n38033), .O(n16623[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_831_4_lut  (.I0(n48382), .I1(\PID_CONTROLLER.integral_23__N_3622 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3620 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_831_4_lut .LUT_INIT = 16'h80c8;
    SB_CARRY add_4081_17 (.CI(n38180), .I0(n12116[14]), .I1(GND_net), 
            .CO(n38181));
    SB_CARRY add_12_17 (.CI(n37298), .I0(n106[15]), .I1(n155[15]), .CO(n37299));
    SB_LUT4 add_4081_16_lut (.I0(GND_net), .I1(n12116[13]), .I2(n1099), 
            .I3(n38179), .O(n9873[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_16 (.CI(n38179), .I0(n12116[13]), .I1(n1099), .CO(n38180));
    SB_CARRY add_5907_9 (.CI(n38033), .I0(n17072[6]), .I1(n609_adj_4631), 
            .CO(n38034));
    SB_LUT4 add_4081_15_lut (.I0(GND_net), .I1(n12116[12]), .I2(n1026), 
            .I3(n38178), .O(n9873[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_15 (.CI(n38178), .I0(n12116[12]), .I1(n1026), .CO(n38179));
    SB_LUT4 add_4081_14_lut (.I0(GND_net), .I1(n12116[11]), .I2(n953), 
            .I3(n38177), .O(n9873[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5907_8_lut (.I0(GND_net), .I1(n17072[5]), .I2(n536_adj_4632), 
            .I3(n38032), .O(n16623[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_14 (.CI(n38177), .I0(n12116[11]), .I1(n953), .CO(n38178));
    SB_CARRY add_5907_8 (.CI(n38032), .I0(n17072[5]), .I1(n536_adj_4632), 
            .CO(n38033));
    SB_LUT4 add_5907_7_lut (.I0(GND_net), .I1(n17072[4]), .I2(n463_adj_4633), 
            .I3(n38031), .O(n16623[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n37297), .O(duty_23__N_3672[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5907_7 (.CI(n38031), .I0(n17072[4]), .I1(n463_adj_4633), 
            .CO(n38032));
    SB_LUT4 add_5907_6_lut (.I0(GND_net), .I1(n17072[3]), .I2(n390_adj_4635), 
            .I3(n38030), .O(n16623[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5907_6 (.CI(n38030), .I0(n17072[3]), .I1(n390_adj_4635), 
            .CO(n38031));
    SB_LUT4 add_4081_13_lut (.I0(GND_net), .I1(n12116[10]), .I2(n880), 
            .I3(n38176), .O(n9873[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_13 (.CI(n38176), .I0(n12116[10]), .I1(n880), .CO(n38177));
    SB_LUT4 add_4081_12_lut (.I0(GND_net), .I1(n12116[9]), .I2(n807), 
            .I3(n38175), .O(n9873[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5907_5_lut (.I0(GND_net), .I1(n17072[2]), .I2(n317_adj_4636), 
            .I3(n38029), .O(n16623[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5907_5 (.CI(n38029), .I0(n17072[2]), .I1(n317_adj_4636), 
            .CO(n38030));
    SB_LUT4 add_5907_4_lut (.I0(GND_net), .I1(n17072[1]), .I2(n244_adj_4637), 
            .I3(n38028), .O(n16623[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_16 (.CI(n37297), .I0(n106[14]), .I1(n155[14]), .CO(n37298));
    SB_CARRY add_5907_4 (.CI(n38028), .I0(n17072[1]), .I1(n244_adj_4637), 
            .CO(n38029));
    SB_CARRY add_4081_12 (.CI(n38175), .I0(n12116[9]), .I1(n807), .CO(n38176));
    SB_LUT4 add_4081_11_lut (.I0(GND_net), .I1(n12116[8]), .I2(n734), 
            .I3(n38174), .O(n9873[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_11 (.CI(n38174), .I0(n12116[8]), .I1(n734), .CO(n38175));
    SB_LUT4 add_5907_3_lut (.I0(GND_net), .I1(n17072[0]), .I2(n171_adj_4638), 
            .I3(n38027), .O(n16623[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4081_10_lut (.I0(GND_net), .I1(n12116[7]), .I2(n661), 
            .I3(n38173), .O(n9873[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_10 (.CI(n38173), .I0(n12116[7]), .I1(n661), .CO(n38174));
    SB_CARRY add_5907_3 (.CI(n38027), .I0(n17072[0]), .I1(n171_adj_4638), 
            .CO(n38028));
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n37296), .O(duty_23__N_3672[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5907_2_lut (.I0(GND_net), .I1(n29_adj_4639), .I2(n98_adj_4640), 
            .I3(GND_net), .O(n16623[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5907_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_15 (.CI(n37296), .I0(n106[13]), .I1(n155[13]), .CO(n37297));
    SB_LUT4 add_4081_9_lut (.I0(GND_net), .I1(n12116[6]), .I2(n588), .I3(n38172), 
            .O(n9873[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_9 (.CI(n38172), .I0(n12116[6]), .I1(n588), .CO(n38173));
    SB_CARRY add_5907_2 (.CI(GND_net), .I0(n29_adj_4639), .I1(n98_adj_4640), 
            .CO(n38027));
    SB_LUT4 add_5935_15_lut (.I0(GND_net), .I1(n17463[12]), .I2(n1050_adj_4641), 
            .I3(n38026), .O(n17072[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5935_14_lut (.I0(GND_net), .I1(n17463[11]), .I2(n977_adj_4642), 
            .I3(n38025), .O(n17072[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4081_8_lut (.I0(GND_net), .I1(n12116[5]), .I2(n515), .I3(n38171), 
            .O(n9873[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n37295), .O(duty_23__N_3672[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5935_14 (.CI(n38025), .I0(n17463[11]), .I1(n977_adj_4642), 
            .CO(n38026));
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4643));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4644));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4645));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4646));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4647));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4648));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4649));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4650));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4651));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4652));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4653));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4654));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4081_8 (.CI(n38171), .I0(n12116[5]), .I1(n515), .CO(n38172));
    SB_LUT4 add_4081_7_lut (.I0(GND_net), .I1(n12116[4]), .I2(n442), .I3(n38170), 
            .O(n9873[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4655));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4656));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_14 (.CI(n37295), .I0(n106[12]), .I1(n155[12]), .CO(n37296));
    SB_LUT4 add_5935_13_lut (.I0(GND_net), .I1(n17463[10]), .I2(n904_adj_4657), 
            .I3(n38024), .O(n17072[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n37294), .O(duty_23__N_3672[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_7 (.CI(n38170), .I0(n12116[4]), .I1(n442), .CO(n38171));
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4081_6_lut (.I0(GND_net), .I1(n12116[3]), .I2(n369), .I3(n38169), 
            .O(n9873[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_13 (.CI(n37294), .I0(n106[11]), .I1(n155[11]), .CO(n37295));
    SB_LUT4 i20640_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20640_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20642_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20642_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4081_6 (.CI(n38169), .I0(n12116[3]), .I1(n369), .CO(n38170));
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3572 [23]), 
            .I1(n9342[21]), .I2(GND_net), .I3(n37801), .O(n8835[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n9342[20]), .I2(GND_net), 
            .I3(n37800), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n37800), .I0(n9342[20]), .I1(GND_net), 
            .CO(n37801));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n9342[19]), .I2(GND_net), 
            .I3(n37799), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n37799), .I0(n9342[19]), .I1(GND_net), 
            .CO(n37800));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n9342[18]), .I2(GND_net), 
            .I3(n37798), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_21 (.CI(n37798), .I0(n9342[18]), .I1(GND_net), 
            .CO(n37799));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n9342[17]), .I2(GND_net), 
            .I3(n37797), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n37797), .I0(n9342[17]), .I1(GND_net), 
            .CO(n37798));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n9342[16]), .I2(GND_net), 
            .I3(n37796), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n37796), .I0(n9342[16]), .I1(GND_net), 
            .CO(n37797));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n9342[15]), .I2(GND_net), 
            .I3(n37795), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_18 (.CI(n37795), .I0(n9342[15]), .I1(GND_net), 
            .CO(n37796));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n9342[14]), .I2(GND_net), 
            .I3(n37794), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5935_13 (.CI(n38024), .I0(n17463[10]), .I1(n904_adj_4657), 
            .CO(n38025));
    SB_LUT4 add_4081_5_lut (.I0(GND_net), .I1(n12116[2]), .I2(n296), .I3(n38168), 
            .O(n9873[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_5 (.CI(n38168), .I0(n12116[2]), .I1(n296), .CO(n38169));
    SB_LUT4 add_4081_4_lut (.I0(GND_net), .I1(n12116[1]), .I2(n223), .I3(n38167), 
            .O(n9873[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5935_12_lut (.I0(GND_net), .I1(n17463[9]), .I2(n831_adj_4664), 
            .I3(n38023), .O(n17072[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n37794), .I0(n9342[14]), .I1(GND_net), 
            .CO(n37795));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n9342[13]), .I2(n1096_adj_4665), 
            .I3(n37793), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n37793), .I0(n9342[13]), .I1(n1096_adj_4665), 
            .CO(n37794));
    SB_CARRY add_5935_12 (.CI(n38023), .I0(n17463[9]), .I1(n831_adj_4664), 
            .CO(n38024));
    SB_LUT4 add_5935_11_lut (.I0(GND_net), .I1(n17463[8]), .I2(n758_adj_4666), 
            .I3(n38022), .O(n17072[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n9342[12]), .I2(n1023_adj_4667), 
            .I3(n37792), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_15 (.CI(n37792), .I0(n9342[12]), .I1(n1023_adj_4667), 
            .CO(n37793));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n9342[11]), .I2(n950_adj_4669), 
            .I3(n37791), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n37791), .I0(n9342[11]), .I1(n950_adj_4669), 
            .CO(n37792));
    SB_CARRY add_5935_11 (.CI(n38022), .I0(n17463[8]), .I1(n758_adj_4666), 
            .CO(n38023));
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n37293), .O(duty_23__N_3672[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n9342[10]), .I2(n877_adj_4671), 
            .I3(n37790), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n37293), .I0(n106[10]), .I1(n155[10]), .CO(n37294));
    SB_CARRY mult_11_add_1225_13 (.CI(n37790), .I0(n9342[10]), .I1(n877_adj_4671), 
            .CO(n37791));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n9342[9]), .I2(n804_adj_4672), 
            .I3(n37789), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n37789), .I0(n9342[9]), .I1(n804_adj_4672), 
            .CO(n37790));
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n9342[8]), .I2(n731_adj_4674), 
            .I3(n37788), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n37788), .I0(n9342[8]), .I1(n731_adj_4674), 
            .CO(n37789));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n9342[7]), .I2(n658_adj_4675), 
            .I3(n37787), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_4 (.CI(n38167), .I0(n12116[1]), .I1(n223), .CO(n38168));
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5935_10_lut (.I0(GND_net), .I1(n17463[7]), .I2(n685_adj_4677), 
            .I3(n38021), .O(n17072[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n37292), 
            .O(duty_23__N_3672[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n37787), .I0(n9342[7]), .I1(n658_adj_4675), 
            .CO(n37788));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n9342[6]), .I2(n585_adj_4679), 
            .I3(n37786), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_9 (.CI(n37786), .I0(n9342[6]), .I1(n585_adj_4679), 
            .CO(n37787));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n9342[5]), .I2(n512_adj_4681), 
            .I3(n37785), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n37785), .I0(n9342[5]), .I1(n512_adj_4681), 
            .CO(n37786));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n9342[4]), .I2(n439_adj_4682), 
            .I3(n37784), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n37784), .I0(n9342[4]), .I1(n439_adj_4682), 
            .CO(n37785));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n9342[3]), .I2(n366_adj_4684), 
            .I3(n37783), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4686));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4687));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_6 (.CI(n37783), .I0(n9342[3]), .I1(n366_adj_4684), 
            .CO(n37784));
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20639_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n9342[2]), .I2(n293_adj_4691), 
            .I3(n37782), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_5 (.CI(n37782), .I0(n9342[2]), .I1(n293_adj_4691), 
            .CO(n37783));
    SB_CARRY add_5935_10 (.CI(n38021), .I0(n17463[7]), .I1(n685_adj_4677), 
            .CO(n38022));
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n9342[1]), .I2(n220_adj_4694), 
            .I3(n37781), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n37781), .I0(n9342[1]), .I1(n220_adj_4694), 
            .CO(n37782));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n9342[0]), .I2(n147_adj_4695), 
            .I3(n37780), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n37780), .I0(n9342[0]), .I1(n147_adj_4695), 
            .CO(n37781));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4696), .I2(n74_adj_4697), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4696), .I1(n74_adj_4697), 
            .CO(n37780));
    SB_LUT4 add_4058_23_lut (.I0(GND_net), .I1(n11631[20]), .I2(GND_net), 
            .I3(n37779), .O(n9342[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4058_22_lut (.I0(GND_net), .I1(n11631[19]), .I2(GND_net), 
            .I3(n37778), .O(n9342[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_22 (.CI(n37778), .I0(n11631[19]), .I1(GND_net), 
            .CO(n37779));
    SB_LUT4 add_4058_21_lut (.I0(GND_net), .I1(n11631[18]), .I2(GND_net), 
            .I3(n37777), .O(n9342[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n37292), .I0(n106[9]), .I1(n155[9]), .CO(n37293));
    SB_CARRY add_4058_21 (.CI(n37777), .I0(n11631[18]), .I1(GND_net), 
            .CO(n37778));
    SB_LUT4 add_4058_20_lut (.I0(GND_net), .I1(n11631[17]), .I2(GND_net), 
            .I3(n37776), .O(n9342[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4058_20 (.CI(n37776), .I0(n11631[17]), .I1(GND_net), 
            .CO(n37777));
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4058_19_lut (.I0(GND_net), .I1(n11631[16]), .I2(GND_net), 
            .I3(n37775), .O(n9342[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4058_19 (.CI(n37775), .I0(n11631[16]), .I1(GND_net), 
            .CO(n37776));
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20638_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20638_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4821[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4058_18_lut (.I0(GND_net), .I1(n11631[15]), .I2(GND_net), 
            .I3(n37774), .O(n9342[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5935_9_lut (.I0(GND_net), .I1(n17463[6]), .I2(n612_adj_4707), 
            .I3(n38020), .O(n17072[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_18 (.CI(n37774), .I0(n11631[15]), .I1(GND_net), 
            .CO(n37775));
    SB_LUT4 add_4081_3_lut (.I0(GND_net), .I1(n12116[0]), .I2(n150_adj_4708), 
            .I3(n38166), .O(n9873[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4058_17_lut (.I0(GND_net), .I1(n11631[14]), .I2(GND_net), 
            .I3(n37773), .O(n9342[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_17 (.CI(n37773), .I0(n11631[14]), .I1(GND_net), 
            .CO(n37774));
    SB_LUT4 add_4058_16_lut (.I0(GND_net), .I1(n11631[13]), .I2(n1099_adj_4710), 
            .I3(n37772), .O(n9342[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5935_9 (.CI(n38020), .I0(n17463[6]), .I1(n612_adj_4707), 
            .CO(n38021));
    SB_CARRY add_4058_16 (.CI(n37772), .I0(n11631[13]), .I1(n1099_adj_4710), 
            .CO(n37773));
    SB_LUT4 add_4058_15_lut (.I0(GND_net), .I1(n11631[12]), .I2(n1026_adj_4711), 
            .I3(n37771), .O(n9342[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4058_15 (.CI(n37771), .I0(n11631[12]), .I1(n1026_adj_4711), 
            .CO(n37772));
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4058_14_lut (.I0(GND_net), .I1(n11631[11]), .I2(n953_adj_4719), 
            .I3(n37770), .O(n9342[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_14 (.CI(n37770), .I0(n11631[11]), .I1(n953_adj_4719), 
            .CO(n37771));
    SB_LUT4 add_4058_13_lut (.I0(GND_net), .I1(n11631[10]), .I2(n880_adj_4720), 
            .I3(n37769), .O(n9342[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n37291), 
            .O(duty_23__N_3672[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5935_8_lut (.I0(GND_net), .I1(n17463[5]), .I2(n539_adj_4721), 
            .I3(n38019), .O(n17072[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_13 (.CI(n37769), .I0(n11631[10]), .I1(n880_adj_4720), 
            .CO(n37770));
    SB_LUT4 add_4058_12_lut (.I0(GND_net), .I1(n11631[9]), .I2(n807_adj_4722), 
            .I3(n37768), .O(n9342[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_12 (.CI(n37768), .I0(n11631[9]), .I1(n807_adj_4722), 
            .CO(n37769));
    SB_CARRY add_12_10 (.CI(n37291), .I0(n106[8]), .I1(n155[8]), .CO(n37292));
    SB_CARRY add_5935_8 (.CI(n38019), .I0(n17463[5]), .I1(n539_adj_4721), 
            .CO(n38020));
    SB_CARRY add_4081_3 (.CI(n38166), .I0(n12116[0]), .I1(n150_adj_4708), 
            .CO(n38167));
    SB_LUT4 add_4058_11_lut (.I0(GND_net), .I1(n11631[8]), .I2(n734_adj_4723), 
            .I3(n37767), .O(n9342[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_11 (.CI(n37767), .I0(n11631[8]), .I1(n734_adj_4723), 
            .CO(n37768));
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4058_10_lut (.I0(GND_net), .I1(n11631[7]), .I2(n661_adj_4725), 
            .I3(n37766), .O(n9342[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_10 (.CI(n37766), .I0(n11631[7]), .I1(n661_adj_4725), 
            .CO(n37767));
    SB_LUT4 add_4058_9_lut (.I0(GND_net), .I1(n11631[6]), .I2(n588_adj_4726), 
            .I3(n37765), .O(n9342[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_9 (.CI(n37765), .I0(n11631[6]), .I1(n588_adj_4726), 
            .CO(n37766));
    SB_LUT4 add_4058_8_lut (.I0(GND_net), .I1(n11631[5]), .I2(n515_adj_4727), 
            .I3(n37764), .O(n9342[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_8 (.CI(n37764), .I0(n11631[5]), .I1(n515_adj_4727), 
            .CO(n37765));
    SB_LUT4 add_4058_7_lut (.I0(GND_net), .I1(n11631[4]), .I2(n442_adj_4728), 
            .I3(n37763), .O(n9342[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4729));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4058_7 (.CI(n37763), .I0(n11631[4]), .I1(n442_adj_4728), 
            .CO(n37764));
    SB_LUT4 add_4058_6_lut (.I0(GND_net), .I1(n11631[3]), .I2(n369_adj_4730), 
            .I3(n37762), .O(n9342[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_6 (.CI(n37762), .I0(n11631[3]), .I1(n369_adj_4730), 
            .CO(n37763));
    SB_LUT4 add_4081_2_lut (.I0(GND_net), .I1(n8_adj_4731), .I2(n77), 
            .I3(GND_net), .O(n9873[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4081_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n37290), 
            .O(duty_23__N_3672[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5935_7_lut (.I0(GND_net), .I1(n17463[4]), .I2(n466_adj_4732), 
            .I3(n38018), .O(n17072[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5935_7 (.CI(n38018), .I0(n17463[4]), .I1(n466_adj_4732), 
            .CO(n38019));
    SB_LUT4 add_4058_5_lut (.I0(GND_net), .I1(n11631[2]), .I2(n296_adj_4733), 
            .I3(n37761), .O(n9342[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_5 (.CI(n37761), .I0(n11631[2]), .I1(n296_adj_4733), 
            .CO(n37762));
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5935_6_lut (.I0(GND_net), .I1(n17463[3]), .I2(n393_adj_4735), 
            .I3(n38017), .O(n17072[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4081_2 (.CI(GND_net), .I0(n8_adj_4731), .I1(n77), .CO(n38166));
    SB_LUT4 add_5326_22_lut (.I0(GND_net), .I1(n13367[19]), .I2(GND_net), 
            .I3(n38165), .O(n12116[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5935_6 (.CI(n38017), .I0(n17463[3]), .I1(n393_adj_4735), 
            .CO(n38018));
    SB_LUT4 add_5326_21_lut (.I0(GND_net), .I1(n13367[18]), .I2(GND_net), 
            .I3(n38164), .O(n12116[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_21 (.CI(n38164), .I0(n13367[18]), .I1(GND_net), 
            .CO(n38165));
    SB_LUT4 add_5326_20_lut (.I0(GND_net), .I1(n13367[17]), .I2(GND_net), 
            .I3(n38163), .O(n12116[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_20 (.CI(n38163), .I0(n13367[17]), .I1(GND_net), 
            .CO(n38164));
    SB_LUT4 add_5935_5_lut (.I0(GND_net), .I1(n17463[2]), .I2(n320_adj_4736), 
            .I3(n38016), .O(n17072[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5326_19_lut (.I0(GND_net), .I1(n13367[16]), .I2(GND_net), 
            .I3(n38162), .O(n12116[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4058_4_lut (.I0(GND_net), .I1(n11631[1]), .I2(n223_adj_4737), 
            .I3(n37760), .O(n9342[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4058_4 (.CI(n37760), .I0(n11631[1]), .I1(n223_adj_4737), 
            .CO(n37761));
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4058_3_lut (.I0(GND_net), .I1(n11631[0]), .I2(n150_adj_4740), 
            .I3(n37759), .O(n9342[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_3 (.CI(n37759), .I0(n11631[0]), .I1(n150_adj_4740), 
            .CO(n37760));
    SB_LUT4 add_4058_2_lut (.I0(GND_net), .I1(n8_adj_4741), .I2(n77_adj_4742), 
            .I3(GND_net), .O(n9342[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4058_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4058_2 (.CI(GND_net), .I0(n8_adj_4741), .I1(n77_adj_4742), 
            .CO(n37759));
    SB_CARRY add_5935_5 (.CI(n38016), .I0(n17463[2]), .I1(n320_adj_4736), 
            .CO(n38017));
    SB_LUT4 add_5935_4_lut (.I0(GND_net), .I1(n17463[1]), .I2(n247_adj_4743), 
            .I3(n38015), .O(n17072[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5935_4 (.CI(n38015), .I0(n17463[1]), .I1(n247_adj_4743), 
            .CO(n38016));
    SB_CARRY add_5326_19 (.CI(n38162), .I0(n13367[16]), .I1(GND_net), 
            .CO(n38163));
    SB_LUT4 add_5935_3_lut (.I0(GND_net), .I1(n17463[0]), .I2(n174_adj_4744), 
            .I3(n38014), .O(n17072[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5326_18_lut (.I0(GND_net), .I1(n13367[15]), .I2(GND_net), 
            .I3(n38161), .O(n12116[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5303_22_lut (.I0(GND_net), .I1(n12927[19]), .I2(GND_net), 
            .I3(n37758), .O(n11631[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_18 (.CI(n38161), .I0(n13367[15]), .I1(GND_net), 
            .CO(n38162));
    SB_LUT4 add_5326_17_lut (.I0(GND_net), .I1(n13367[14]), .I2(GND_net), 
            .I3(n38160), .O(n12116[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_17 (.CI(n38160), .I0(n13367[14]), .I1(GND_net), 
            .CO(n38161));
    SB_LUT4 add_5326_16_lut (.I0(GND_net), .I1(n13367[13]), .I2(n1102), 
            .I3(n38159), .O(n12116[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_16 (.CI(n38159), .I0(n13367[13]), .I1(n1102), .CO(n38160));
    SB_LUT4 add_5326_15_lut (.I0(GND_net), .I1(n13367[12]), .I2(n1029), 
            .I3(n38158), .O(n12116[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_15 (.CI(n38158), .I0(n13367[12]), .I1(n1029), .CO(n38159));
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5303_21_lut (.I0(GND_net), .I1(n12927[18]), .I2(GND_net), 
            .I3(n37757), .O(n11631[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5303_21 (.CI(n37757), .I0(n12927[18]), .I1(GND_net), 
            .CO(n37758));
    SB_CARRY add_5935_3 (.CI(n38014), .I0(n17463[0]), .I1(n174_adj_4744), 
            .CO(n38015));
    SB_LUT4 add_5326_14_lut (.I0(GND_net), .I1(n13367[11]), .I2(n956), 
            .I3(n38157), .O(n12116[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5935_2_lut (.I0(GND_net), .I1(n32_adj_4749), .I2(n101_adj_4750), 
            .I3(GND_net), .O(n17072[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5935_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5303_20_lut (.I0(GND_net), .I1(n12927[17]), .I2(GND_net), 
            .I3(n37756), .O(n11631[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_20 (.CI(n37756), .I0(n12927[17]), .I1(GND_net), 
            .CO(n37757));
    SB_LUT4 add_5303_19_lut (.I0(GND_net), .I1(n12927[16]), .I2(GND_net), 
            .I3(n37755), .O(n11631[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_9 (.CI(n37290), .I0(n106[7]), .I1(n155[7]), .CO(n37291));
    SB_CARRY add_5303_19 (.CI(n37755), .I0(n12927[16]), .I1(GND_net), 
            .CO(n37756));
    SB_LUT4 add_5303_18_lut (.I0(GND_net), .I1(n12927[15]), .I2(GND_net), 
            .I3(n37754), .O(n11631[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n37289), 
            .O(duty_23__N_3672[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_18 (.CI(n37754), .I0(n12927[15]), .I1(GND_net), 
            .CO(n37755));
    SB_LUT4 add_5303_17_lut (.I0(GND_net), .I1(n12927[14]), .I2(GND_net), 
            .I3(n37753), .O(n11631[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_17 (.CI(n37753), .I0(n12927[14]), .I1(GND_net), 
            .CO(n37754));
    SB_LUT4 add_5303_16_lut (.I0(GND_net), .I1(n12927[13]), .I2(n1102_adj_4752), 
            .I3(n37752), .O(n11631[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_16 (.CI(n37752), .I0(n12927[13]), .I1(n1102_adj_4752), 
            .CO(n37753));
    SB_LUT4 add_5303_15_lut (.I0(GND_net), .I1(n12927[12]), .I2(n1029_adj_4753), 
            .I3(n37751), .O(n11631[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_15 (.CI(n37751), .I0(n12927[12]), .I1(n1029_adj_4753), 
            .CO(n37752));
    SB_CARRY add_5326_14 (.CI(n38157), .I0(n13367[11]), .I1(n956), .CO(n38158));
    SB_LUT4 add_5303_14_lut (.I0(GND_net), .I1(n12927[11]), .I2(n956_adj_4754), 
            .I3(n37750), .O(n11631[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_14 (.CI(n37750), .I0(n12927[11]), .I1(n956_adj_4754), 
            .CO(n37751));
    SB_LUT4 add_5326_13_lut (.I0(GND_net), .I1(n13367[10]), .I2(n883), 
            .I3(n38156), .O(n12116[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_13_lut (.I0(GND_net), .I1(n12927[10]), .I2(n883_adj_4755), 
            .I3(n37749), .O(n11631[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_8 (.CI(n37289), .I0(n106[6]), .I1(n155[6]), .CO(n37290));
    SB_CARRY add_5935_2 (.CI(GND_net), .I0(n32_adj_4749), .I1(n101_adj_4750), 
            .CO(n38014));
    SB_CARRY add_5326_13 (.CI(n38156), .I0(n13367[10]), .I1(n883), .CO(n38157));
    SB_LUT4 add_5326_12_lut (.I0(GND_net), .I1(n13367[9]), .I2(n810), 
            .I3(n38155), .O(n12116[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5961_14_lut (.I0(GND_net), .I1(n17800[11]), .I2(n980_adj_4756), 
            .I3(n38013), .O(n17463[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_13 (.CI(n37749), .I0(n12927[10]), .I1(n883_adj_4755), 
            .CO(n37750));
    SB_LUT4 add_5303_12_lut (.I0(GND_net), .I1(n12927[9]), .I2(n810_adj_4757), 
            .I3(n37748), .O(n11631[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_12 (.CI(n37748), .I0(n12927[9]), .I1(n810_adj_4757), 
            .CO(n37749));
    SB_CARRY add_5326_12 (.CI(n38155), .I0(n13367[9]), .I1(n810), .CO(n38156));
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5961_13_lut (.I0(GND_net), .I1(n17800[10]), .I2(n907_adj_4758), 
            .I3(n38012), .O(n17463[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_13 (.CI(n38012), .I0(n17800[10]), .I1(n907_adj_4758), 
            .CO(n38013));
    SB_LUT4 add_5961_12_lut (.I0(GND_net), .I1(n17800[9]), .I2(n834_adj_4759), 
            .I3(n38011), .O(n17463[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5326_11_lut (.I0(GND_net), .I1(n13367[8]), .I2(n737), 
            .I3(n38154), .O(n12116[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_12 (.CI(n38011), .I0(n17800[9]), .I1(n834_adj_4759), 
            .CO(n38012));
    SB_CARRY add_5326_11 (.CI(n38154), .I0(n13367[8]), .I1(n737), .CO(n38155));
    SB_LUT4 add_5326_10_lut (.I0(GND_net), .I1(n13367[7]), .I2(n664), 
            .I3(n38153), .O(n12116[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_10 (.CI(n38153), .I0(n13367[7]), .I1(n664), .CO(n38154));
    SB_LUT4 add_5961_11_lut (.I0(GND_net), .I1(n17800[8]), .I2(n761_adj_4760), 
            .I3(n38010), .O(n17463[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5326_9_lut (.I0(GND_net), .I1(n13367[6]), .I2(n591), .I3(n38152), 
            .O(n12116[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_11_lut (.I0(GND_net), .I1(n12927[8]), .I2(n737_adj_4761), 
            .I3(n37747), .O(n11631[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_11 (.CI(n38010), .I0(n17800[8]), .I1(n761_adj_4760), 
            .CO(n38011));
    SB_CARRY add_5326_9 (.CI(n38152), .I0(n13367[6]), .I1(n591), .CO(n38153));
    SB_LUT4 add_5326_8_lut (.I0(GND_net), .I1(n13367[5]), .I2(n518), .I3(n38151), 
            .O(n12116[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_11 (.CI(n37747), .I0(n12927[8]), .I1(n737_adj_4761), 
            .CO(n37748));
    SB_LUT4 add_5303_10_lut (.I0(GND_net), .I1(n12927[7]), .I2(n664_adj_4762), 
            .I3(n37746), .O(n11631[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4765));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4766));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4768));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4769));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5303_10 (.CI(n37746), .I0(n12927[7]), .I1(n664_adj_4762), 
            .CO(n37747));
    SB_LUT4 add_5303_9_lut (.I0(GND_net), .I1(n12927[6]), .I2(n591_adj_4771), 
            .I3(n37745), .O(n11631[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_9 (.CI(n37745), .I0(n12927[6]), .I1(n591_adj_4771), 
            .CO(n37746));
    SB_LUT4 add_5303_8_lut (.I0(GND_net), .I1(n12927[5]), .I2(n518_adj_4772), 
            .I3(n37744), .O(n11631[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_8 (.CI(n37744), .I0(n12927[5]), .I1(n518_adj_4772), 
            .CO(n37745));
    SB_LUT4 add_5303_7_lut (.I0(GND_net), .I1(n12927[4]), .I2(n445), .I3(n37743), 
            .O(n11631[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_7 (.CI(n37743), .I0(n12927[4]), .I1(n445), .CO(n37744));
    SB_LUT4 add_5303_6_lut (.I0(GND_net), .I1(n12927[3]), .I2(n372), .I3(n37742), 
            .O(n11631[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_6 (.CI(n37742), .I0(n12927[3]), .I1(n372), .CO(n37743));
    SB_CARRY add_5326_8 (.CI(n38151), .I0(n13367[5]), .I1(n518), .CO(n38152));
    SB_LUT4 add_5303_5_lut (.I0(GND_net), .I1(n12927[2]), .I2(n299_adj_4773), 
            .I3(n37741), .O(n11631[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4774));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5326_7_lut (.I0(GND_net), .I1(n13367[4]), .I2(n445_adj_4775), 
            .I3(n38150), .O(n12116[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_7 (.CI(n38150), .I0(n13367[4]), .I1(n445_adj_4775), 
            .CO(n38151));
    SB_CARRY add_5303_5 (.CI(n37741), .I0(n12927[2]), .I1(n299_adj_4773), 
            .CO(n37742));
    SB_LUT4 add_5326_6_lut (.I0(GND_net), .I1(n13367[3]), .I2(n372_adj_4776), 
            .I3(n38149), .O(n12116[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5961_10_lut (.I0(GND_net), .I1(n17800[7]), .I2(n688_adj_4774), 
            .I3(n38009), .O(n17463[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_4_lut (.I0(GND_net), .I1(n12927[1]), .I2(n226_adj_4770), 
            .I3(n37740), .O(n11631[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_10 (.CI(n38009), .I0(n17800[7]), .I1(n688_adj_4774), 
            .CO(n38010));
    SB_LUT4 add_5961_9_lut (.I0(GND_net), .I1(n17800[6]), .I2(n615_adj_4769), 
            .I3(n38008), .O(n17463[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_4 (.CI(n37740), .I0(n12927[1]), .I1(n226_adj_4770), 
            .CO(n37741));
    SB_LUT4 add_5303_3_lut (.I0(GND_net), .I1(n12927[0]), .I2(n153_adj_4768), 
            .I3(n37739), .O(n11631[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_6 (.CI(n38149), .I0(n13367[3]), .I1(n372_adj_4776), 
            .CO(n38150));
    SB_CARRY add_5961_9 (.CI(n38008), .I0(n17800[6]), .I1(n615_adj_4769), 
            .CO(n38009));
    SB_LUT4 add_5961_8_lut (.I0(GND_net), .I1(n17800[5]), .I2(n542_adj_4767), 
            .I3(n38007), .O(n17463[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_8 (.CI(n38007), .I0(n17800[5]), .I1(n542_adj_4767), 
            .CO(n38008));
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4776));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5303_3 (.CI(n37739), .I0(n12927[0]), .I1(n153_adj_4768), 
            .CO(n37740));
    SB_LUT4 add_5961_7_lut (.I0(GND_net), .I1(n17800[4]), .I2(n469_adj_4766), 
            .I3(n38006), .O(n17463[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_2_lut (.I0(GND_net), .I1(n11_adj_4765), .I2(n80_adj_4764), 
            .I3(GND_net), .O(n11631[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_2 (.CI(GND_net), .I0(n11_adj_4765), .I1(n80_adj_4764), 
            .CO(n37739));
    SB_LUT4 add_5716_21_lut (.I0(GND_net), .I1(n13768[18]), .I2(GND_net), 
            .I3(n37738), .O(n12927[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5716_20_lut (.I0(GND_net), .I1(n13768[17]), .I2(GND_net), 
            .I3(n37737), .O(n12927[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_20 (.CI(n37737), .I0(n13768[17]), .I1(GND_net), 
            .CO(n37738));
    SB_LUT4 add_5716_19_lut (.I0(GND_net), .I1(n13768[16]), .I2(GND_net), 
            .I3(n37736), .O(n12927[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_7 (.CI(n38006), .I0(n17800[4]), .I1(n469_adj_4766), 
            .CO(n38007));
    SB_CARRY add_5716_19 (.CI(n37736), .I0(n13768[16]), .I1(GND_net), 
            .CO(n37737));
    SB_LUT4 add_5716_18_lut (.I0(GND_net), .I1(n13768[15]), .I2(GND_net), 
            .I3(n37735), .O(n12927[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_18 (.CI(n37735), .I0(n13768[15]), .I1(GND_net), 
            .CO(n37736));
    SB_LUT4 add_5326_5_lut (.I0(GND_net), .I1(n13367[2]), .I2(n299), .I3(n38148), 
            .O(n12116[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_5 (.CI(n38148), .I0(n13367[2]), .I1(n299), .CO(n38149));
    SB_LUT4 add_5716_17_lut (.I0(GND_net), .I1(n13768[14]), .I2(GND_net), 
            .I3(n37734), .O(n12927[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5326_4_lut (.I0(GND_net), .I1(n13367[1]), .I2(n226), .I3(n38147), 
            .O(n12116[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_4 (.CI(n38147), .I0(n13367[1]), .I1(n226), .CO(n38148));
    SB_LUT4 add_5961_6_lut (.I0(GND_net), .I1(n17800[3]), .I2(n396_adj_4729), 
            .I3(n38005), .O(n17463[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_17 (.CI(n37734), .I0(n13768[14]), .I1(GND_net), 
            .CO(n37735));
    SB_CARRY add_5961_6 (.CI(n38005), .I0(n17800[3]), .I1(n396_adj_4729), 
            .CO(n38006));
    SB_LUT4 add_5716_16_lut (.I0(GND_net), .I1(n13768[13]), .I2(n1105_adj_4687), 
            .I3(n37733), .O(n12927[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_16 (.CI(n37733), .I0(n13768[13]), .I1(n1105_adj_4687), 
            .CO(n37734));
    SB_LUT4 add_5716_15_lut (.I0(GND_net), .I1(n13768[12]), .I2(n1032_adj_4686), 
            .I3(n37732), .O(n12927[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5961_5_lut (.I0(GND_net), .I1(n17800[2]), .I2(n323_adj_4656), 
            .I3(n38004), .O(n17463[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_5 (.CI(n38004), .I0(n17800[2]), .I1(n323_adj_4656), 
            .CO(n38005));
    SB_LUT4 add_5961_4_lut (.I0(GND_net), .I1(n17800[1]), .I2(n250_adj_4655), 
            .I3(n38003), .O(n17463[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_4 (.CI(n38003), .I0(n17800[1]), .I1(n250_adj_4655), 
            .CO(n38004));
    SB_LUT4 add_5961_3_lut (.I0(GND_net), .I1(n17800[0]), .I2(n177_adj_4654), 
            .I3(n38002), .O(n17463[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_3 (.CI(n38002), .I0(n17800[0]), .I1(n177_adj_4654), 
            .CO(n38003));
    SB_LUT4 add_5326_3_lut (.I0(GND_net), .I1(n13367[0]), .I2(n153_adj_4653), 
            .I3(n38146), .O(n12116[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_3 (.CI(n38146), .I0(n13367[0]), .I1(n153_adj_4653), 
            .CO(n38147));
    SB_CARRY add_5716_15 (.CI(n37732), .I0(n13768[12]), .I1(n1032_adj_4686), 
            .CO(n37733));
    SB_LUT4 add_5716_14_lut (.I0(GND_net), .I1(n13768[11]), .I2(n959_adj_4652), 
            .I3(n37731), .O(n12927[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5326_2_lut (.I0(GND_net), .I1(n11_adj_4651), .I2(n80), 
            .I3(GND_net), .O(n12116[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_2 (.CI(GND_net), .I0(n11_adj_4651), .I1(n80), .CO(n38146));
    SB_LUT4 add_5961_2_lut (.I0(GND_net), .I1(n35_adj_4650), .I2(n104_adj_4649), 
            .I3(GND_net), .O(n17463[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_2 (.CI(GND_net), .I0(n35_adj_4650), .I1(n104_adj_4649), 
            .CO(n38002));
    SB_LUT4 add_5736_21_lut (.I0(GND_net), .I1(n14167[18]), .I2(GND_net), 
            .I3(n38145), .O(n13367[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_14 (.CI(n37731), .I0(n13768[11]), .I1(n959_adj_4652), 
            .CO(n37732));
    SB_LUT4 add_5985_13_lut (.I0(GND_net), .I1(n18087[10]), .I2(n910_adj_4648), 
            .I3(n38001), .O(n17800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5716_13_lut (.I0(GND_net), .I1(n13768[10]), .I2(n886_adj_4647), 
            .I3(n37730), .O(n12927[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n37288), 
            .O(duty_23__N_3672[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_13 (.CI(n37730), .I0(n13768[10]), .I1(n886_adj_4647), 
            .CO(n37731));
    SB_LUT4 add_5716_12_lut (.I0(GND_net), .I1(n13768[9]), .I2(n813_adj_4646), 
            .I3(n37729), .O(n12927[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5736_20_lut (.I0(GND_net), .I1(n14167[17]), .I2(GND_net), 
            .I3(n38144), .O(n13367[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5985_12_lut (.I0(GND_net), .I1(n18087[9]), .I2(n837_adj_4645), 
            .I3(n38000), .O(n17800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_12 (.CI(n37729), .I0(n13768[9]), .I1(n813_adj_4646), 
            .CO(n37730));
    SB_LUT4 add_5716_11_lut (.I0(GND_net), .I1(n13768[8]), .I2(n740_adj_4644), 
            .I3(n37728), .O(n12927[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_11 (.CI(n37728), .I0(n13768[8]), .I1(n740_adj_4644), 
            .CO(n37729));
    SB_LUT4 add_5716_10_lut (.I0(GND_net), .I1(n13768[7]), .I2(n667_adj_4643), 
            .I3(n37727), .O(n12927[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_20 (.CI(n38144), .I0(n14167[17]), .I1(GND_net), 
            .CO(n38145));
    SB_CARRY add_5985_12 (.CI(n38000), .I0(n18087[9]), .I1(n837_adj_4645), 
            .CO(n38001));
    SB_LUT4 add_5736_19_lut (.I0(GND_net), .I1(n14167[16]), .I2(GND_net), 
            .I3(n38143), .O(n13367[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_19 (.CI(n38143), .I0(n14167[16]), .I1(GND_net), 
            .CO(n38144));
    SB_LUT4 add_5736_18_lut (.I0(GND_net), .I1(n14167[15]), .I2(GND_net), 
            .I3(n38142), .O(n13367[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5985_11_lut (.I0(GND_net), .I1(n18087[8]), .I2(n764_adj_4629), 
            .I3(n37999), .O(n17800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_10 (.CI(n37727), .I0(n13768[7]), .I1(n667_adj_4643), 
            .CO(n37728));
    SB_LUT4 add_5716_9_lut (.I0(GND_net), .I1(n13768[6]), .I2(n594_adj_4627), 
            .I3(n37726), .O(n12927[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_9 (.CI(n37726), .I0(n13768[6]), .I1(n594_adj_4627), 
            .CO(n37727));
    SB_CARRY add_5736_18 (.CI(n38142), .I0(n14167[15]), .I1(GND_net), 
            .CO(n38143));
    SB_CARRY add_5985_11 (.CI(n37999), .I0(n18087[8]), .I1(n764_adj_4629), 
            .CO(n38000));
    SB_LUT4 add_5716_8_lut (.I0(GND_net), .I1(n13768[5]), .I2(n521_adj_4624), 
            .I3(n37725), .O(n12927[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5736_17_lut (.I0(GND_net), .I1(n14167[14]), .I2(GND_net), 
            .I3(n38141), .O(n13367[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5985_10_lut (.I0(GND_net), .I1(n18087[7]), .I2(n691_adj_4623), 
            .I3(n37998), .O(n17800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_8 (.CI(n37725), .I0(n13768[5]), .I1(n521_adj_4624), 
            .CO(n37726));
    SB_LUT4 add_5716_7_lut (.I0(GND_net), .I1(n13768[4]), .I2(n448_adj_4619), 
            .I3(n37724), .O(n12927[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_7 (.CI(n37724), .I0(n13768[4]), .I1(n448_adj_4619), 
            .CO(n37725));
    SB_LUT4 add_5716_6_lut (.I0(GND_net), .I1(n13768[3]), .I2(n375_adj_4618), 
            .I3(n37723), .O(n12927[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_17 (.CI(n38141), .I0(n14167[14]), .I1(GND_net), 
            .CO(n38142));
    SB_CARRY add_5985_10 (.CI(n37998), .I0(n18087[7]), .I1(n691_adj_4623), 
            .CO(n37999));
    SB_CARRY add_5716_6 (.CI(n37723), .I0(n13768[3]), .I1(n375_adj_4618), 
            .CO(n37724));
    SB_LUT4 add_5985_9_lut (.I0(GND_net), .I1(n18087[6]), .I2(n618_adj_4617), 
            .I3(n37997), .O(n17800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n37288), .I0(n106[5]), .I1(n155[5]), .CO(n37289));
    SB_LUT4 add_5716_5_lut (.I0(GND_net), .I1(n13768[2]), .I2(n302_adj_4616), 
            .I3(n37722), .O(n12927[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_5 (.CI(n37722), .I0(n13768[2]), .I1(n302_adj_4616), 
            .CO(n37723));
    SB_LUT4 add_5736_16_lut (.I0(GND_net), .I1(n14167[13]), .I2(n1105), 
            .I3(n38140), .O(n13367[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5985_9 (.CI(n37997), .I0(n18087[6]), .I1(n618_adj_4617), 
            .CO(n37998));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n37287), 
            .O(duty_23__N_3672[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5716_4_lut (.I0(GND_net), .I1(n13768[1]), .I2(n229_adj_4613), 
            .I3(n37721), .O(n12927[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_4 (.CI(n37721), .I0(n13768[1]), .I1(n229_adj_4613), 
            .CO(n37722));
    SB_LUT4 add_5716_3_lut (.I0(GND_net), .I1(n13768[0]), .I2(n156_adj_4609), 
            .I3(n37720), .O(n12927[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5716_3 (.CI(n37720), .I0(n13768[0]), .I1(n156_adj_4609), 
            .CO(n37721));
    SB_LUT4 add_5716_2_lut (.I0(GND_net), .I1(n14_adj_4608), .I2(n83_adj_4605), 
            .I3(GND_net), .O(n12927[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5716_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_16 (.CI(n38140), .I0(n14167[13]), .I1(n1105), .CO(n38141));
    SB_LUT4 add_5736_15_lut (.I0(GND_net), .I1(n14167[12]), .I2(n1032), 
            .I3(n38139), .O(n13367[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5985_8_lut (.I0(GND_net), .I1(n18087[5]), .I2(n545_adj_4604), 
            .I3(n37996), .O(n17800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5985_8 (.CI(n37996), .I0(n18087[5]), .I1(n545_adj_4604), 
            .CO(n37997));
    SB_CARRY add_5716_2 (.CI(GND_net), .I0(n14_adj_4608), .I1(n83_adj_4605), 
            .CO(n37720));
    SB_LUT4 add_6027_11_lut (.I0(GND_net), .I1(n18527[8]), .I2(n770_adj_4603), 
            .I3(n37719), .O(n18328[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_15 (.CI(n38139), .I0(n14167[12]), .I1(n1032), .CO(n38140));
    SB_LUT4 add_6027_10_lut (.I0(GND_net), .I1(n18527[7]), .I2(n697_adj_4602), 
            .I3(n37718), .O(n18328[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5985_7_lut (.I0(GND_net), .I1(n18087[4]), .I2(n472_adj_4601), 
            .I3(n37995), .O(n17800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_10 (.CI(n37718), .I0(n18527[7]), .I1(n697_adj_4602), 
            .CO(n37719));
    SB_LUT4 add_6027_9_lut (.I0(GND_net), .I1(n18527[6]), .I2(n624_adj_4587), 
            .I3(n37717), .O(n18328[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_9 (.CI(n37717), .I0(n18527[6]), .I1(n624_adj_4587), 
            .CO(n37718));
    SB_LUT4 add_6027_8_lut (.I0(GND_net), .I1(n18527[5]), .I2(n551_adj_4586), 
            .I3(n37716), .O(n18328[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_8 (.CI(n37716), .I0(n18527[5]), .I1(n551_adj_4586), 
            .CO(n37717));
    SB_CARRY add_5985_7 (.CI(n37995), .I0(n18087[4]), .I1(n472_adj_4601), 
            .CO(n37996));
    SB_CARRY add_12_6 (.CI(n37287), .I0(n106[4]), .I1(n155[4]), .CO(n37288));
    SB_LUT4 add_6027_7_lut (.I0(GND_net), .I1(n18527[4]), .I2(n478_adj_4563), 
            .I3(n37715), .O(n18328[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_7 (.CI(n37715), .I0(n18527[4]), .I1(n478_adj_4563), 
            .CO(n37716));
    SB_LUT4 add_6027_6_lut (.I0(GND_net), .I1(n18527[3]), .I2(n405_adj_4562), 
            .I3(n37714), .O(n18328[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5736_14_lut (.I0(GND_net), .I1(n14167[11]), .I2(n959), 
            .I3(n38138), .O(n13367[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5985_6_lut (.I0(GND_net), .I1(n18087[3]), .I2(n399_adj_4561), 
            .I3(n37994), .O(n17800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_6 (.CI(n37714), .I0(n18527[3]), .I1(n405_adj_4562), 
            .CO(n37715));
    SB_LUT4 add_6027_5_lut (.I0(GND_net), .I1(n18527[2]), .I2(n332_adj_4560), 
            .I3(n37713), .O(n18328[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_14 (.CI(n38138), .I0(n14167[11]), .I1(n959), .CO(n38139));
    SB_CARRY add_5985_6 (.CI(n37994), .I0(n18087[3]), .I1(n399_adj_4561), 
            .CO(n37995));
    SB_CARRY add_6027_5 (.CI(n37713), .I0(n18527[2]), .I1(n332_adj_4560), 
            .CO(n37714));
    SB_LUT4 add_6027_4_lut (.I0(GND_net), .I1(n18527[1]), .I2(n259_adj_4559), 
            .I3(n37712), .O(n18328[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_4 (.CI(n37712), .I0(n18527[1]), .I1(n259_adj_4559), 
            .CO(n37713));
    SB_LUT4 add_6027_3_lut (.I0(GND_net), .I1(n18527[0]), .I2(n186_adj_4557), 
            .I3(n37711), .O(n18328[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_3 (.CI(n37711), .I0(n18527[0]), .I1(n186_adj_4557), 
            .CO(n37712));
    SB_LUT4 add_5985_5_lut (.I0(GND_net), .I1(n18087[2]), .I2(n326_adj_4556), 
            .I3(n37993), .O(n17800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6027_2_lut (.I0(GND_net), .I1(n44_adj_4555), .I2(n113_adj_4551), 
            .I3(GND_net), .O(n18328[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6027_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6027_2 (.CI(GND_net), .I0(n44_adj_4555), .I1(n113_adj_4551), 
            .CO(n37711));
    SB_LUT4 add_5756_20_lut (.I0(GND_net), .I1(n14528[17]), .I2(GND_net), 
            .I3(n37704), .O(n13768[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5756_19_lut (.I0(GND_net), .I1(n14528[16]), .I2(GND_net), 
            .I3(n37703), .O(n13768[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_19 (.CI(n37703), .I0(n14528[16]), .I1(GND_net), 
            .CO(n37704));
    SB_LUT4 add_5756_18_lut (.I0(GND_net), .I1(n14528[15]), .I2(GND_net), 
            .I3(n37702), .O(n13768[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_18 (.CI(n37702), .I0(n14528[15]), .I1(GND_net), 
            .CO(n37703));
    SB_LUT4 add_5756_17_lut (.I0(GND_net), .I1(n14528[14]), .I2(GND_net), 
            .I3(n37701), .O(n13768[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_17 (.CI(n37701), .I0(n14528[14]), .I1(GND_net), 
            .CO(n37702));
    SB_LUT4 add_5756_16_lut (.I0(GND_net), .I1(n14528[13]), .I2(n1108_adj_4550), 
            .I3(n37700), .O(n13768[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_16 (.CI(n37700), .I0(n14528[13]), .I1(n1108_adj_4550), 
            .CO(n37701));
    SB_LUT4 add_5756_15_lut (.I0(GND_net), .I1(n14528[12]), .I2(n1035_adj_4549), 
            .I3(n37699), .O(n13768[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_15 (.CI(n37699), .I0(n14528[12]), .I1(n1035_adj_4549), 
            .CO(n37700));
    SB_LUT4 add_5756_14_lut (.I0(GND_net), .I1(n14528[11]), .I2(n962_adj_4548), 
            .I3(n37698), .O(n13768[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n37286), 
            .O(duty_23__N_3672[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_14 (.CI(n37698), .I0(n14528[11]), .I1(n962_adj_4548), 
            .CO(n37699));
    SB_LUT4 add_5756_13_lut (.I0(GND_net), .I1(n14528[10]), .I2(n889_adj_4547), 
            .I3(n37697), .O(n13768[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_13 (.CI(n37697), .I0(n14528[10]), .I1(n889_adj_4547), 
            .CO(n37698));
    SB_LUT4 add_5756_12_lut (.I0(GND_net), .I1(n14528[9]), .I2(n816_adj_4546), 
            .I3(n37696), .O(n13768[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_12 (.CI(n37696), .I0(n14528[9]), .I1(n816_adj_4546), 
            .CO(n37697));
    SB_LUT4 add_5756_11_lut (.I0(GND_net), .I1(n14528[8]), .I2(n743_adj_4545), 
            .I3(n37695), .O(n13768[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_11 (.CI(n37695), .I0(n14528[8]), .I1(n743_adj_4545), 
            .CO(n37696));
    SB_CARRY add_5985_5 (.CI(n37993), .I0(n18087[2]), .I1(n326_adj_4556), 
            .CO(n37994));
    SB_LUT4 add_5736_13_lut (.I0(GND_net), .I1(n14167[10]), .I2(n886), 
            .I3(n38137), .O(n13367[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5756_10_lut (.I0(GND_net), .I1(n14528[7]), .I2(n670_adj_4544), 
            .I3(n37694), .O(n13768[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5985_4_lut (.I0(GND_net), .I1(n18087[1]), .I2(n253_adj_4543), 
            .I3(n37992), .O(n17800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_10 (.CI(n37694), .I0(n14528[7]), .I1(n670_adj_4544), 
            .CO(n37695));
    SB_LUT4 add_5756_9_lut (.I0(GND_net), .I1(n14528[6]), .I2(n597_adj_4542), 
            .I3(n37693), .O(n13768[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_9 (.CI(n37693), .I0(n14528[6]), .I1(n597_adj_4542), 
            .CO(n37694));
    SB_LUT4 add_5756_8_lut (.I0(GND_net), .I1(n14528[5]), .I2(n524_adj_4541), 
            .I3(n37692), .O(n13768[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_8 (.CI(n37692), .I0(n14528[5]), .I1(n524_adj_4541), 
            .CO(n37693));
    SB_LUT4 add_5756_7_lut (.I0(GND_net), .I1(n14528[4]), .I2(n451_adj_4540), 
            .I3(n37691), .O(n13768[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_7 (.CI(n37691), .I0(n14528[4]), .I1(n451_adj_4540), 
            .CO(n37692));
    SB_LUT4 add_5756_6_lut (.I0(GND_net), .I1(n14528[3]), .I2(n378_adj_4539), 
            .I3(n37690), .O(n13768[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_6 (.CI(n37690), .I0(n14528[3]), .I1(n378_adj_4539), 
            .CO(n37691));
    SB_LUT4 add_5756_5_lut (.I0(GND_net), .I1(n14528[2]), .I2(n305_adj_4538), 
            .I3(n37689), .O(n13768[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_5 (.CI(n37689), .I0(n14528[2]), .I1(n305_adj_4538), 
            .CO(n37690));
    SB_LUT4 add_5756_4_lut (.I0(GND_net), .I1(n14528[1]), .I2(n232_adj_4537), 
            .I3(n37688), .O(n13768[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_4 (.CI(n37688), .I0(n14528[1]), .I1(n232_adj_4537), 
            .CO(n37689));
    SB_LUT4 add_5756_3_lut (.I0(GND_net), .I1(n14528[0]), .I2(n159_adj_4536), 
            .I3(n37687), .O(n13768[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_3 (.CI(n37687), .I0(n14528[0]), .I1(n159_adj_4536), 
            .CO(n37688));
    SB_LUT4 add_5756_2_lut (.I0(GND_net), .I1(n17_adj_4535), .I2(n86_adj_4534), 
            .I3(GND_net), .O(n13768[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5756_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5756_2 (.CI(GND_net), .I0(n17_adj_4535), .I1(n86_adj_4534), 
            .CO(n37687));
    SB_LUT4 add_5793_19_lut (.I0(GND_net), .I1(n15212[16]), .I2(GND_net), 
            .I3(n37686), .O(n14528[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5793_18_lut (.I0(GND_net), .I1(n15212[15]), .I2(GND_net), 
            .I3(n37685), .O(n14528[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_18 (.CI(n37685), .I0(n15212[15]), .I1(GND_net), 
            .CO(n37686));
    SB_LUT4 add_5793_17_lut (.I0(GND_net), .I1(n15212[14]), .I2(GND_net), 
            .I3(n37684), .O(n14528[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_17 (.CI(n37684), .I0(n15212[14]), .I1(GND_net), 
            .CO(n37685));
    SB_LUT4 add_5793_16_lut (.I0(GND_net), .I1(n15212[13]), .I2(n1111_adj_4533), 
            .I3(n37683), .O(n14528[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5736_13 (.CI(n38137), .I0(n14167[10]), .I1(n886), .CO(n38138));
    SB_CARRY add_5985_4 (.CI(n37992), .I0(n18087[1]), .I1(n253_adj_4543), 
            .CO(n37993));
    SB_CARRY add_5793_16 (.CI(n37683), .I0(n15212[13]), .I1(n1111_adj_4533), 
            .CO(n37684));
    SB_LUT4 add_5793_15_lut (.I0(GND_net), .I1(n15212[12]), .I2(n1038_adj_4532), 
            .I3(n37682), .O(n14528[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_15 (.CI(n37682), .I0(n15212[12]), .I1(n1038_adj_4532), 
            .CO(n37683));
    SB_LUT4 add_5985_3_lut (.I0(GND_net), .I1(n18087[0]), .I2(n180_adj_4531), 
            .I3(n37991), .O(n17800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5793_14_lut (.I0(GND_net), .I1(n15212[11]), .I2(n965_adj_4530), 
            .I3(n37681), .O(n14528[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_14 (.CI(n37681), .I0(n15212[11]), .I1(n965_adj_4530), 
            .CO(n37682));
    SB_LUT4 add_5736_12_lut (.I0(GND_net), .I1(n14167[9]), .I2(n813), 
            .I3(n38136), .O(n13367[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5985_3 (.CI(n37991), .I0(n18087[0]), .I1(n180_adj_4531), 
            .CO(n37992));
    SB_LUT4 add_5793_13_lut (.I0(GND_net), .I1(n15212[10]), .I2(n892_adj_4529), 
            .I3(n37680), .O(n14528[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_12 (.CI(n38136), .I0(n14167[9]), .I1(n813), .CO(n38137));
    SB_CARRY add_5793_13 (.CI(n37680), .I0(n15212[10]), .I1(n892_adj_4529), 
            .CO(n37681));
    SB_LUT4 add_5793_12_lut (.I0(GND_net), .I1(n15212[9]), .I2(n819_adj_4528), 
            .I3(n37679), .O(n14528[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5736_11_lut (.I0(GND_net), .I1(n14167[8]), .I2(n740), 
            .I3(n38135), .O(n13367[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_12 (.CI(n37679), .I0(n15212[9]), .I1(n819_adj_4528), 
            .CO(n37680));
    SB_LUT4 add_5793_11_lut (.I0(GND_net), .I1(n15212[8]), .I2(n746_adj_4527), 
            .I3(n37678), .O(n14528[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_11 (.CI(n37678), .I0(n15212[8]), .I1(n746_adj_4527), 
            .CO(n37679));
    SB_LUT4 add_5985_2_lut (.I0(GND_net), .I1(n38_adj_4526), .I2(n107_adj_4525), 
            .I3(GND_net), .O(n17800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5985_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_11 (.CI(n38135), .I0(n14167[8]), .I1(n740), .CO(n38136));
    SB_LUT4 add_5793_10_lut (.I0(GND_net), .I1(n15212[7]), .I2(n673_adj_4524), 
            .I3(n37677), .O(n14528[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4775));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5793_10 (.CI(n37677), .I0(n15212[7]), .I1(n673_adj_4524), 
            .CO(n37678));
    SB_LUT4 add_5736_10_lut (.I0(GND_net), .I1(n14167[7]), .I2(n667), 
            .I3(n38134), .O(n13367[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5793_9_lut (.I0(GND_net), .I1(n15212[6]), .I2(n600_adj_4523), 
            .I3(n37676), .O(n14528[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_9 (.CI(n37676), .I0(n15212[6]), .I1(n600_adj_4523), 
            .CO(n37677));
    SB_LUT4 add_5793_8_lut (.I0(GND_net), .I1(n15212[5]), .I2(n527_adj_4522), 
            .I3(n37675), .O(n14528[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_10 (.CI(n38134), .I0(n14167[7]), .I1(n667), .CO(n38135));
    SB_CARRY add_5793_8 (.CI(n37675), .I0(n15212[5]), .I1(n527_adj_4522), 
            .CO(n37676));
    SB_LUT4 add_5793_7_lut (.I0(GND_net), .I1(n15212[4]), .I2(n454_adj_4521), 
            .I3(n37674), .O(n14528[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_7 (.CI(n37674), .I0(n15212[4]), .I1(n454_adj_4521), 
            .CO(n37675));
    SB_CARRY add_5985_2 (.CI(GND_net), .I0(n38_adj_4526), .I1(n107_adj_4525), 
            .CO(n37991));
    SB_LUT4 add_5793_6_lut (.I0(GND_net), .I1(n15212[3]), .I2(n381), .I3(n37673), 
            .O(n14528[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_6 (.CI(n37673), .I0(n15212[3]), .I1(n381), .CO(n37674));
    SB_LUT4 add_5793_5_lut (.I0(GND_net), .I1(n15212[2]), .I2(n308), .I3(n37672), 
            .O(n14528[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_5 (.CI(n37672), .I0(n15212[2]), .I1(n308), .CO(n37673));
    SB_LUT4 add_5793_4_lut (.I0(GND_net), .I1(n15212[1]), .I2(n235), .I3(n37671), 
            .O(n14528[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5736_9_lut (.I0(GND_net), .I1(n14167[6]), .I2(n594), .I3(n38133), 
            .O(n13367[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_4 (.CI(n37671), .I0(n15212[1]), .I1(n235), .CO(n37672));
    SB_LUT4 add_5793_3_lut (.I0(GND_net), .I1(n15212[0]), .I2(n162), .I3(n37670), 
            .O(n14528[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_3 (.CI(n37670), .I0(n15212[0]), .I1(n162), .CO(n37671));
    SB_CARRY add_12_5 (.CI(n37286), .I0(n106[3]), .I1(n155[3]), .CO(n37287));
    SB_LUT4 add_5793_2_lut (.I0(GND_net), .I1(n20_adj_4520), .I2(n89), 
            .I3(GND_net), .O(n14528[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5793_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5793_2 (.CI(GND_net), .I0(n20_adj_4520), .I1(n89), .CO(n37670));
    SB_LUT4 add_6045_10_lut (.I0(GND_net), .I1(n18688[7]), .I2(n700_adj_4519), 
            .I3(n37669), .O(n18527[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6045_9_lut (.I0(GND_net), .I1(n18688[6]), .I2(n627_adj_4518), 
            .I3(n37668), .O(n18527[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_9 (.CI(n38133), .I0(n14167[6]), .I1(n594), .CO(n38134));
    SB_CARRY add_6045_9 (.CI(n37668), .I0(n18688[6]), .I1(n627_adj_4518), 
            .CO(n37669));
    SB_LUT4 add_6045_8_lut (.I0(GND_net), .I1(n18688[5]), .I2(n554_adj_4517), 
            .I3(n37667), .O(n18527[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6045_8 (.CI(n37667), .I0(n18688[5]), .I1(n554_adj_4517), 
            .CO(n37668));
    SB_LUT4 add_5736_8_lut (.I0(GND_net), .I1(n14167[5]), .I2(n521), .I3(n38132), 
            .O(n13367[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n37285), 
            .O(duty_23__N_3672[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6045_7_lut (.I0(GND_net), .I1(n18688[4]), .I2(n481_adj_4516), 
            .I3(n37666), .O(n18527[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6045_7 (.CI(n37666), .I0(n18688[4]), .I1(n481_adj_4516), 
            .CO(n37667));
    SB_CARRY add_12_4 (.CI(n37285), .I0(n106[2]), .I1(n155[2]), .CO(n37286));
    SB_LUT4 add_6045_6_lut (.I0(GND_net), .I1(n18688[3]), .I2(n408_adj_4515), 
            .I3(n37665), .O(n18527[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n37284), 
            .O(duty_23__N_3672[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6045_6 (.CI(n37665), .I0(n18688[3]), .I1(n408_adj_4515), 
            .CO(n37666));
    SB_LUT4 add_6045_5_lut (.I0(GND_net), .I1(n18688[2]), .I2(n335_adj_4514), 
            .I3(n37664), .O(n18527[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6045_5 (.CI(n37664), .I0(n18688[2]), .I1(n335_adj_4514), 
            .CO(n37665));
    SB_LUT4 add_6045_4_lut (.I0(GND_net), .I1(n18688[1]), .I2(n262_adj_4513), 
            .I3(n37663), .O(n18527[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6045_4 (.CI(n37663), .I0(n18688[1]), .I1(n262_adj_4513), 
            .CO(n37664));
    SB_CARRY add_5736_8 (.CI(n38132), .I0(n14167[5]), .I1(n521), .CO(n38133));
    SB_LUT4 add_6045_3_lut (.I0(GND_net), .I1(n18688[0]), .I2(n189_adj_4512), 
            .I3(n37662), .O(n18527[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6045_3 (.CI(n37662), .I0(n18688[0]), .I1(n189_adj_4512), 
            .CO(n37663));
    SB_LUT4 add_6045_2_lut (.I0(GND_net), .I1(n47_adj_4511), .I2(n116_adj_4510), 
            .I3(GND_net), .O(n18527[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6045_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6045_2 (.CI(GND_net), .I0(n47_adj_4511), .I1(n116_adj_4510), 
            .CO(n37662));
    SB_CARRY add_12_3 (.CI(n37284), .I0(n106[1]), .I1(n155[1]), .CO(n37285));
    SB_LUT4 add_5828_18_lut (.I0(GND_net), .I1(n15824[15]), .I2(GND_net), 
            .I3(n37661), .O(n15212[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5828_17_lut (.I0(GND_net), .I1(n15824[14]), .I2(GND_net), 
            .I3(n37660), .O(n15212[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_17 (.CI(n37660), .I0(n15824[14]), .I1(GND_net), 
            .CO(n37661));
    SB_LUT4 add_5828_16_lut (.I0(GND_net), .I1(n15824[13]), .I2(n1114_adj_4509), 
            .I3(n37659), .O(n15212[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5736_7_lut (.I0(GND_net), .I1(n14167[4]), .I2(n448), .I3(n38131), 
            .O(n13367[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_16 (.CI(n37659), .I0(n15824[13]), .I1(n1114_adj_4509), 
            .CO(n37660));
    SB_LUT4 add_5828_15_lut (.I0(GND_net), .I1(n15824[12]), .I2(n1041_adj_4508), 
            .I3(n37658), .O(n15212[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_15 (.CI(n37658), .I0(n15824[12]), .I1(n1041_adj_4508), 
            .CO(n37659));
    SB_LUT4 add_5828_14_lut (.I0(GND_net), .I1(n15824[11]), .I2(n968_adj_4507), 
            .I3(n37657), .O(n15212[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_14 (.CI(n37657), .I0(n15824[11]), .I1(n968_adj_4507), 
            .CO(n37658));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3672[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5828_13_lut (.I0(GND_net), .I1(n15824[10]), .I2(n895_adj_4506), 
            .I3(n37656), .O(n15212[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_13 (.CI(n37656), .I0(n15824[10]), .I1(n895_adj_4506), 
            .CO(n37657));
    SB_LUT4 add_5828_12_lut (.I0(GND_net), .I1(n15824[9]), .I2(n822_adj_4505), 
            .I3(n37655), .O(n15212[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_7 (.CI(n38131), .I0(n14167[4]), .I1(n448), .CO(n38132));
    SB_LUT4 add_5736_6_lut (.I0(GND_net), .I1(n14167[3]), .I2(n375), .I3(n38130), 
            .O(n13367[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_6 (.CI(n38130), .I0(n14167[3]), .I1(n375), .CO(n38131));
    SB_CARRY add_5828_12 (.CI(n37655), .I0(n15824[9]), .I1(n822_adj_4505), 
            .CO(n37656));
    SB_LUT4 add_5828_11_lut (.I0(GND_net), .I1(n15824[8]), .I2(n749_adj_4504), 
            .I3(n37654), .O(n15212[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_11 (.CI(n37654), .I0(n15824[8]), .I1(n749_adj_4504), 
            .CO(n37655));
    SB_LUT4 add_5828_10_lut (.I0(GND_net), .I1(n15824[7]), .I2(n676_adj_4503), 
            .I3(n37653), .O(n15212[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_10 (.CI(n37653), .I0(n15824[7]), .I1(n676_adj_4503), 
            .CO(n37654));
    SB_LUT4 add_5828_9_lut (.I0(GND_net), .I1(n15824[6]), .I2(n603_adj_4502), 
            .I3(n37652), .O(n15212[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_9 (.CI(n37652), .I0(n15824[6]), .I1(n603_adj_4502), 
            .CO(n37653));
    SB_LUT4 add_5828_8_lut (.I0(GND_net), .I1(n15824[5]), .I2(n530_adj_4501), 
            .I3(n37651), .O(n15212[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_8 (.CI(n37651), .I0(n15824[5]), .I1(n530_adj_4501), 
            .CO(n37652));
    SB_LUT4 add_5828_7_lut (.I0(GND_net), .I1(n15824[4]), .I2(n457_adj_4500), 
            .I3(n37650), .O(n15212[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_7 (.CI(n37650), .I0(n15824[4]), .I1(n457_adj_4500), 
            .CO(n37651));
    SB_LUT4 add_5736_5_lut (.I0(GND_net), .I1(n14167[2]), .I2(n302), .I3(n38129), 
            .O(n13367[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5828_6_lut (.I0(GND_net), .I1(n15824[3]), .I2(n384_adj_4499), 
            .I3(n37649), .O(n15212[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_6 (.CI(n37649), .I0(n15824[3]), .I1(n384_adj_4499), 
            .CO(n37650));
    SB_LUT4 add_5828_5_lut (.I0(GND_net), .I1(n15824[2]), .I2(n311_adj_4498), 
            .I3(n37648), .O(n15212[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_5 (.CI(n37648), .I0(n15824[2]), .I1(n311_adj_4498), 
            .CO(n37649));
    SB_LUT4 add_5828_4_lut (.I0(GND_net), .I1(n15824[1]), .I2(n238_adj_4497), 
            .I3(n37647), .O(n15212[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_4 (.CI(n37647), .I0(n15824[1]), .I1(n238_adj_4497), 
            .CO(n37648));
    SB_LUT4 add_5828_3_lut (.I0(GND_net), .I1(n15824[0]), .I2(n165_adj_4496), 
            .I3(n37646), .O(n15212[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_3 (.CI(n37646), .I0(n15824[0]), .I1(n165_adj_4496), 
            .CO(n37647));
    SB_LUT4 add_5828_2_lut (.I0(GND_net), .I1(n23_adj_4495), .I2(n92_adj_4494), 
            .I3(GND_net), .O(n15212[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5828_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5828_2 (.CI(GND_net), .I0(n23_adj_4495), .I1(n92_adj_4494), 
            .CO(n37646));
    SB_LUT4 add_5861_17_lut (.I0(GND_net), .I1(n16368[14]), .I2(GND_net), 
            .I3(n37645), .O(n15824[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5861_16_lut (.I0(GND_net), .I1(n16368[13]), .I2(n1117_adj_4493), 
            .I3(n37644), .O(n15824[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23933_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(n36929), .I3(n19072[0]), .O(n4_adj_4778));   // verilog/motorControl.v(34[25:36])
    defparam i23933_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n37284));
    SB_CARRY add_5861_16 (.CI(n37644), .I0(n16368[13]), .I1(n1117_adj_4493), 
            .CO(n37645));
    SB_CARRY add_5736_5 (.CI(n38129), .I0(n14167[2]), .I1(n302), .CO(n38130));
    SB_LUT4 add_5736_4_lut (.I0(GND_net), .I1(n14167[1]), .I2(n229), .I3(n38128), 
            .O(n13367[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5861_15_lut (.I0(GND_net), .I1(n16368[12]), .I2(n1044_adj_4492), 
            .I3(n37643), .O(n15824[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_15 (.CI(n37643), .I0(n16368[12]), .I1(n1044_adj_4492), 
            .CO(n37644));
    SB_LUT4 add_5861_14_lut (.I0(GND_net), .I1(n16368[11]), .I2(n971_adj_4491), 
            .I3(n37642), .O(n15824[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_14 (.CI(n37642), .I0(n16368[11]), .I1(n971_adj_4491), 
            .CO(n37643));
    SB_LUT4 add_5861_13_lut (.I0(GND_net), .I1(n16368[10]), .I2(n898_adj_4490), 
            .I3(n37641), .O(n15824[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_13 (.CI(n37641), .I0(n16368[10]), .I1(n898_adj_4490), 
            .CO(n37642));
    SB_LUT4 add_5861_12_lut (.I0(GND_net), .I1(n16368[9]), .I2(n825_adj_4489), 
            .I3(n37640), .O(n15824[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_12 (.CI(n37640), .I0(n16368[9]), .I1(n825_adj_4489), 
            .CO(n37641));
    SB_LUT4 add_5861_11_lut (.I0(GND_net), .I1(n16368[8]), .I2(n752_adj_4488), 
            .I3(n37639), .O(n15824[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_11 (.CI(n37639), .I0(n16368[8]), .I1(n752_adj_4488), 
            .CO(n37640));
    SB_LUT4 add_5861_10_lut (.I0(GND_net), .I1(n16368[7]), .I2(n679_adj_4487), 
            .I3(n37638), .O(n15824[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_4 (.CI(n38128), .I0(n14167[1]), .I1(n229), .CO(n38129));
    SB_CARRY add_5861_10 (.CI(n37638), .I0(n16368[7]), .I1(n679_adj_4487), 
            .CO(n37639));
    SB_LUT4 add_5861_9_lut (.I0(GND_net), .I1(n16368[6]), .I2(n606_adj_4486), 
            .I3(n37637), .O(n15824[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_9 (.CI(n37637), .I0(n16368[6]), .I1(n606_adj_4486), 
            .CO(n37638));
    SB_LUT4 add_5736_3_lut (.I0(GND_net), .I1(n14167[0]), .I2(n156), .I3(n38127), 
            .O(n13367[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5861_8_lut (.I0(GND_net), .I1(n16368[5]), .I2(n533_adj_4485), 
            .I3(n37636), .O(n15824[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_8 (.CI(n37636), .I0(n16368[5]), .I1(n533_adj_4485), 
            .CO(n37637));
    SB_LUT4 add_5861_7_lut (.I0(GND_net), .I1(n16368[4]), .I2(n460_adj_4484), 
            .I3(n37635), .O(n15824[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5736_3 (.CI(n38127), .I0(n14167[0]), .I1(n156), .CO(n38128));
    SB_CARRY add_5861_7 (.CI(n37635), .I0(n16368[4]), .I1(n460_adj_4484), 
            .CO(n37636));
    SB_LUT4 add_5861_6_lut (.I0(GND_net), .I1(n16368[3]), .I2(n387_adj_4483), 
            .I3(n37634), .O(n15824[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_6 (.CI(n37634), .I0(n16368[3]), .I1(n387_adj_4483), 
            .CO(n37635));
    SB_LUT4 add_5861_5_lut (.I0(GND_net), .I1(n16368[2]), .I2(n314_adj_4482), 
            .I3(n37633), .O(n15824[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_5 (.CI(n37633), .I0(n16368[2]), .I1(n314_adj_4482), 
            .CO(n37634));
    SB_LUT4 add_5861_4_lut (.I0(GND_net), .I1(n16368[1]), .I2(n241_adj_4481), 
            .I3(n37632), .O(n15824[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_4 (.CI(n37632), .I0(n16368[1]), .I1(n241_adj_4481), 
            .CO(n37633));
    SB_LUT4 add_5861_3_lut (.I0(GND_net), .I1(n16368[0]), .I2(n168_adj_4480), 
            .I3(n37631), .O(n15824[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5736_2_lut (.I0(GND_net), .I1(n14_adj_4479), .I2(n83), 
            .I3(GND_net), .O(n13367[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5736_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_3 (.CI(n37631), .I0(n16368[0]), .I1(n168_adj_4480), 
            .CO(n37632));
    SB_CARRY add_5736_2 (.CI(GND_net), .I0(n14_adj_4479), .I1(n83), .CO(n38127));
    SB_LUT4 add_5861_2_lut (.I0(GND_net), .I1(n26_adj_4477), .I2(n95), 
            .I3(GND_net), .O(n15824[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5861_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5861_2 (.CI(GND_net), .I0(n26_adj_4477), .I1(n95), .CO(n37631));
    SB_LUT4 add_6061_9_lut (.I0(GND_net), .I1(n18815[6]), .I2(n630_adj_4476), 
            .I3(n37630), .O(n18688[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6061_8_lut (.I0(GND_net), .I1(n18815[5]), .I2(n557), .I3(n37629), 
            .O(n18688[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_8 (.CI(n37629), .I0(n18815[5]), .I1(n557), .CO(n37630));
    SB_LUT4 add_6061_7_lut (.I0(GND_net), .I1(n18815[4]), .I2(n484), .I3(n37628), 
            .O(n18688[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_7 (.CI(n37628), .I0(n18815[4]), .I1(n484), .CO(n37629));
    SB_LUT4 add_6061_6_lut (.I0(GND_net), .I1(n18815[3]), .I2(n411), .I3(n37627), 
            .O(n18688[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(n19072[0]), .I3(n36929), .O(n19048[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_CARRY add_6061_6 (.CI(n37627), .I0(n18815[3]), .I1(n411), .CO(n37628));
    SB_LUT4 i23920_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [20]), .I3(\Ki[1] ), 
            .O(n19048[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23920_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_6061_5_lut (.I0(GND_net), .I1(n18815[2]), .I2(n338), .I3(n37626), 
            .O(n18688[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23922_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [20]), .I3(\Ki[1] ), 
            .O(n36929));   // verilog/motorControl.v(34[25:36])
    defparam i23922_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_6061_5 (.CI(n37626), .I0(n18815[2]), .I1(n338), .CO(n37627));
    SB_LUT4 add_6061_4_lut (.I0(GND_net), .I1(n18815[1]), .I2(n265_adj_4475), 
            .I3(n37625), .O(n18688[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_4 (.CI(n37625), .I0(n18815[1]), .I1(n265_adj_4475), 
            .CO(n37626));
    SB_LUT4 add_6061_3_lut (.I0(GND_net), .I1(n18815[0]), .I2(n192), .I3(n37624), 
            .O(n18688[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_3 (.CI(n37624), .I0(n18815[0]), .I1(n192), .CO(n37625));
    SB_LUT4 add_6061_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n18688[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5775_20_lut (.I0(GND_net), .I1(n14888[17]), .I2(GND_net), 
            .I3(n38126), .O(n14167[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n37624));
    SB_LUT4 add_5892_16_lut (.I0(GND_net), .I1(n16848[13]), .I2(n1120), 
            .I3(n37623), .O(n16368[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5892_15_lut (.I0(GND_net), .I1(n16848[12]), .I2(n1047), 
            .I3(n37622), .O(n16368[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_15 (.CI(n37622), .I0(n16848[12]), .I1(n1047), .CO(n37623));
    SB_LUT4 add_5892_14_lut (.I0(GND_net), .I1(n16848[11]), .I2(n974), 
            .I3(n37621), .O(n16368[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_14 (.CI(n37621), .I0(n16848[11]), .I1(n974), .CO(n37622));
    SB_LUT4 add_5892_13_lut (.I0(GND_net), .I1(n16848[10]), .I2(n901), 
            .I3(n37620), .O(n16368[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_13 (.CI(n37620), .I0(n16848[10]), .I1(n901), .CO(n37621));
    SB_LUT4 add_5775_19_lut (.I0(GND_net), .I1(n14888[16]), .I2(GND_net), 
            .I3(n38125), .O(n14167[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5892_12_lut (.I0(GND_net), .I1(n16848[9]), .I2(n828), 
            .I3(n37619), .O(n16368[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_12 (.CI(n37619), .I0(n16848[9]), .I1(n828), .CO(n37620));
    SB_CARRY add_5775_19 (.CI(n38125), .I0(n14888[16]), .I1(GND_net), 
            .CO(n38126));
    SB_LUT4 add_5892_11_lut (.I0(GND_net), .I1(n16848[8]), .I2(n755), 
            .I3(n37618), .O(n16368[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_11 (.CI(n37618), .I0(n16848[8]), .I1(n755), .CO(n37619));
    SB_LUT4 add_5775_18_lut (.I0(GND_net), .I1(n14888[15]), .I2(GND_net), 
            .I3(n38124), .O(n14167[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23971_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(n36970), .I3(n19048[0]), .O(n4_adj_4779));   // verilog/motorControl.v(34[25:36])
    defparam i23971_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_5775_18 (.CI(n38124), .I0(n14888[15]), .I1(GND_net), 
            .CO(n38125));
    SB_LUT4 i2_3_lut_4_lut_adj_1516 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(n19048[0]), .I3(n36970), .O(n19008[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1516.LUT_INIT = 16'h8778;
    SB_LUT4 add_5892_10_lut (.I0(GND_net), .I1(n16848[7]), .I2(n682), 
            .I3(n37617), .O(n16368[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_10 (.CI(n37617), .I0(n16848[7]), .I1(n682), .CO(n37618));
    SB_LUT4 add_5892_9_lut (.I0(GND_net), .I1(n16848[6]), .I2(n609), .I3(n37616), 
            .O(n16368[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5775_17_lut (.I0(GND_net), .I1(n14888[14]), .I2(GND_net), 
            .I3(n38123), .O(n14167[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_9 (.CI(n37616), .I0(n16848[6]), .I1(n609), .CO(n37617));
    SB_LUT4 add_5892_8_lut (.I0(GND_net), .I1(n16848[5]), .I2(n536), .I3(n37615), 
            .O(n16368[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_8 (.CI(n37615), .I0(n16848[5]), .I1(n536), .CO(n37616));
    SB_LUT4 add_5892_7_lut (.I0(GND_net), .I1(n16848[4]), .I2(n463), .I3(n37614), 
            .O(n16368[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_7 (.CI(n37614), .I0(n16848[4]), .I1(n463), .CO(n37615));
    SB_LUT4 add_5892_6_lut (.I0(GND_net), .I1(n16848[3]), .I2(n390), .I3(n37613), 
            .O(n16368[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_17 (.CI(n38123), .I0(n14888[14]), .I1(GND_net), 
            .CO(n38124));
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5892_6 (.CI(n37613), .I0(n16848[3]), .I1(n390), .CO(n37614));
    SB_LUT4 add_5775_16_lut (.I0(GND_net), .I1(n14888[13]), .I2(n1108), 
            .I3(n38122), .O(n14167[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5892_5_lut (.I0(GND_net), .I1(n16848[2]), .I2(n317), .I3(n37612), 
            .O(n16368[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_5 (.CI(n37612), .I0(n16848[2]), .I1(n317), .CO(n37613));
    SB_LUT4 add_5892_4_lut (.I0(GND_net), .I1(n16848[1]), .I2(n244), .I3(n37611), 
            .O(n16368[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_4 (.CI(n37611), .I0(n16848[1]), .I1(n244), .CO(n37612));
    SB_LUT4 add_5892_3_lut (.I0(GND_net), .I1(n16848[0]), .I2(n171), .I3(n37610), 
            .O(n16368[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5892_3 (.CI(n37610), .I0(n16848[0]), .I1(n171), .CO(n37611));
    SB_CARRY add_5775_16 (.CI(n38122), .I0(n14888[13]), .I1(n1108), .CO(n38123));
    SB_LUT4 i23958_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [19]), .I3(\Ki[1] ), 
            .O(n19008[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23958_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_5775_15_lut (.I0(GND_net), .I1(n14888[12]), .I2(n1035), 
            .I3(n38121), .O(n14167[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5892_2_lut (.I0(GND_net), .I1(n29_adj_4470), .I2(n98), 
            .I3(GND_net), .O(n16368[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5892_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_15 (.CI(n38121), .I0(n14888[12]), .I1(n1035), .CO(n38122));
    SB_CARRY add_5892_2 (.CI(GND_net), .I0(n29_adj_4470), .I1(n98), .CO(n37610));
    SB_LUT4 i23960_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [19]), .I3(\Ki[1] ), 
            .O(n36970));   // verilog/motorControl.v(34[25:36])
    defparam i23960_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_5775_14_lut (.I0(GND_net), .I1(n14888[11]), .I2(n962), 
            .I3(n38120), .O(n14167[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24010_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n4_adj_4781), .I3(n19008[1]), .O(n6_adj_4782));   // verilog/motorControl.v(34[25:36])
    defparam i24010_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_5775_14 (.CI(n38120), .I0(n14888[11]), .I1(n962), .CO(n38121));
    SB_LUT4 add_5775_13_lut (.I0(GND_net), .I1(n14888[10]), .I2(n889), 
            .I3(n38119), .O(n14167[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1517 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n19008[1]), .I3(n4_adj_4781), .O(n18948[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1517.LUT_INIT = 16'h8778;
    SB_CARRY add_5775_13 (.CI(n38119), .I0(n14888[10]), .I1(n889), .CO(n38120));
    SB_LUT4 add_5775_12_lut (.I0(GND_net), .I1(n14888[9]), .I2(n816), 
            .I3(n38118), .O(n14167[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4773));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5775_12 (.CI(n38118), .I0(n14888[9]), .I1(n816), .CO(n38119));
    SB_LUT4 i2_3_lut_4_lut_adj_1518 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n19008[0]), .I3(n37004), .O(n18948[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1518.LUT_INIT = 16'h8778;
    SB_LUT4 add_5921_15_lut (.I0(GND_net), .I1(n17268[12]), .I2(n1050), 
            .I3(n37598), .O(n16848[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5921_14_lut (.I0(GND_net), .I1(n17268[11]), .I2(n977), 
            .I3(n37597), .O(n16848[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24002_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n37004), .I3(n19008[0]), .O(n4_adj_4781));   // verilog/motorControl.v(34[25:36])
    defparam i24002_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_5775_11_lut (.I0(GND_net), .I1(n14888[8]), .I2(n743), 
            .I3(n38117), .O(n14167[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_11 (.CI(n38117), .I0(n14888[8]), .I1(n743), .CO(n38118));
    SB_CARRY add_5921_14 (.CI(n37597), .I0(n17268[11]), .I1(n977), .CO(n37598));
    SB_LUT4 add_5775_10_lut (.I0(GND_net), .I1(n14888[7]), .I2(n670), 
            .I3(n38116), .O(n14167[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5921_13_lut (.I0(GND_net), .I1(n17268[10]), .I2(n904), 
            .I3(n37596), .O(n16848[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_13 (.CI(n37596), .I0(n17268[10]), .I1(n904), .CO(n37597));
    SB_LUT4 add_5921_12_lut (.I0(GND_net), .I1(n17268[9]), .I2(n831), 
            .I3(n37595), .O(n16848[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_12 (.CI(n37595), .I0(n17268[9]), .I1(n831), .CO(n37596));
    SB_LUT4 add_5921_11_lut (.I0(GND_net), .I1(n17268[8]), .I2(n758), 
            .I3(n37594), .O(n16848[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_11 (.CI(n37594), .I0(n17268[8]), .I1(n758), .CO(n37595));
    SB_LUT4 add_5921_10_lut (.I0(GND_net), .I1(n17268[7]), .I2(n685), 
            .I3(n37593), .O(n16848[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_10 (.CI(n37593), .I0(n17268[7]), .I1(n685), .CO(n37594));
    SB_CARRY add_5775_10 (.CI(n38116), .I0(n14888[7]), .I1(n670), .CO(n38117));
    SB_LUT4 add_5921_9_lut (.I0(GND_net), .I1(n17268[6]), .I2(n612), .I3(n37592), 
            .O(n16848[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_9 (.CI(n37592), .I0(n17268[6]), .I1(n612), .CO(n37593));
    SB_LUT4 add_5921_8_lut (.I0(GND_net), .I1(n17268[5]), .I2(n539), .I3(n37591), 
            .O(n16848[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_8 (.CI(n37591), .I0(n17268[5]), .I1(n539), .CO(n37592));
    SB_LUT4 add_5921_7_lut (.I0(GND_net), .I1(n17268[4]), .I2(n466), .I3(n37590), 
            .O(n16848[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5775_9_lut (.I0(GND_net), .I1(n14888[6]), .I2(n597), .I3(n38115), 
            .O(n14167[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_9 (.CI(n38115), .I0(n14888[6]), .I1(n597), .CO(n38116));
    SB_CARRY add_5921_7 (.CI(n37590), .I0(n17268[4]), .I1(n466), .CO(n37591));
    SB_LUT4 add_5921_6_lut (.I0(GND_net), .I1(n17268[3]), .I2(n393), .I3(n37589), 
            .O(n16848[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_6 (.CI(n37589), .I0(n17268[3]), .I1(n393), .CO(n37590));
    SB_LUT4 add_5921_5_lut (.I0(GND_net), .I1(n17268[2]), .I2(n320), .I3(n37588), 
            .O(n16848[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5921_5 (.CI(n37588), .I0(n17268[2]), .I1(n320), .CO(n37589));
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5921_4_lut (.I0(GND_net), .I1(n17268[1]), .I2(n247), .I3(n37587), 
            .O(n16848[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5775_8_lut (.I0(GND_net), .I1(n14888[5]), .I2(n524), .I3(n38114), 
            .O(n14167[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4772));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5921_4 (.CI(n37587), .I0(n17268[1]), .I1(n247), .CO(n37588));
    SB_LUT4 add_5921_3_lut (.I0(GND_net), .I1(n17268[0]), .I2(n174), .I3(n37586), 
            .O(n16848[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20637_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20637_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5921_3 (.CI(n37586), .I0(n17268[0]), .I1(n174), .CO(n37587));
    SB_LUT4 add_5921_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n16848[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5921_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_8 (.CI(n38114), .I0(n14888[5]), .I1(n524), .CO(n38115));
    SB_CARRY add_5921_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n37586));
    SB_LUT4 add_6075_8_lut (.I0(GND_net), .I1(n18912[5]), .I2(n560), .I3(n37585), 
            .O(n18815[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6075_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6075_7_lut (.I0(GND_net), .I1(n18912[4]), .I2(n487), .I3(n37584), 
            .O(n18815[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6075_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5775_7_lut (.I0(GND_net), .I1(n14888[4]), .I2(n451), .I3(n38113), 
            .O(n14167[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6075_7 (.CI(n37584), .I0(n18912[4]), .I1(n487), .CO(n37585));
    SB_LUT4 add_6075_6_lut (.I0(GND_net), .I1(n18912[3]), .I2(n414), .I3(n37583), 
            .O(n18815[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6075_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6075_6 (.CI(n37583), .I0(n18912[3]), .I1(n414), .CO(n37584));
    SB_LUT4 add_6075_5_lut (.I0(GND_net), .I1(n18912[2]), .I2(n341), .I3(n37582), 
            .O(n18815[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6075_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6075_5 (.CI(n37582), .I0(n18912[2]), .I1(n341), .CO(n37583));
    SB_LUT4 add_6075_4_lut (.I0(GND_net), .I1(n18912[1]), .I2(n268), .I3(n37581), 
            .O(n18815[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6075_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_7 (.CI(n38113), .I0(n14888[4]), .I1(n451), .CO(n38114));
    SB_CARRY add_6075_4 (.CI(n37581), .I0(n18912[1]), .I1(n268), .CO(n37582));
    SB_LUT4 add_6075_3_lut (.I0(GND_net), .I1(n18912[0]), .I2(n195), .I3(n37580), 
            .O(n18815[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6075_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6075_3 (.CI(n37580), .I0(n18912[0]), .I1(n195), .CO(n37581));
    SB_LUT4 add_6075_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n18815[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6075_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6075_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n37580));
    SB_LUT4 add_5775_6_lut (.I0(GND_net), .I1(n14888[3]), .I2(n378), .I3(n38112), 
            .O(n14167[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5948_14_lut (.I0(GND_net), .I1(n17632[11]), .I2(n980), 
            .I3(n37579), .O(n17268[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5948_13_lut (.I0(GND_net), .I1(n17632[10]), .I2(n907), 
            .I3(n37578), .O(n17268[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_13 (.CI(n37578), .I0(n17632[10]), .I1(n907), .CO(n37579));
    SB_LUT4 add_5948_12_lut (.I0(GND_net), .I1(n17632[9]), .I2(n834), 
            .I3(n37577), .O(n17268[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_12 (.CI(n37577), .I0(n17632[9]), .I1(n834), .CO(n37578));
    SB_LUT4 add_5948_11_lut (.I0(GND_net), .I1(n17632[8]), .I2(n761), 
            .I3(n37576), .O(n17268[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_11 (.CI(n37576), .I0(n17632[8]), .I1(n761), .CO(n37577));
    SB_CARRY add_5775_6 (.CI(n38112), .I0(n14888[3]), .I1(n378), .CO(n38113));
    SB_LUT4 add_5948_10_lut (.I0(GND_net), .I1(n17632[7]), .I2(n688), 
            .I3(n37575), .O(n17268[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4822[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5775_5_lut (.I0(GND_net), .I1(n14888[2]), .I2(n305), .I3(n38111), 
            .O(n14167[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_10 (.CI(n37575), .I0(n17632[7]), .I1(n688), .CO(n37576));
    SB_CARRY add_5775_5 (.CI(n38111), .I0(n14888[2]), .I1(n305), .CO(n38112));
    SB_LUT4 add_5948_9_lut (.I0(GND_net), .I1(n17632[6]), .I2(n615), .I3(n37574), 
            .O(n17268[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_9 (.CI(n37574), .I0(n17632[6]), .I1(n615), .CO(n37575));
    SB_LUT4 add_5948_8_lut (.I0(GND_net), .I1(n17632[5]), .I2(n542), .I3(n37573), 
            .O(n17268[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_8 (.CI(n37573), .I0(n17632[5]), .I1(n542), .CO(n37574));
    SB_LUT4 add_5775_4_lut (.I0(GND_net), .I1(n14888[1]), .I2(n232), .I3(n38110), 
            .O(n14167[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5948_7_lut (.I0(GND_net), .I1(n17632[4]), .I2(n469), .I3(n37572), 
            .O(n17268[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_7 (.CI(n37572), .I0(n17632[4]), .I1(n469), .CO(n37573));
    SB_LUT4 add_5948_6_lut (.I0(GND_net), .I1(n17632[3]), .I2(n396), .I3(n37571), 
            .O(n17268[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_6 (.CI(n37571), .I0(n17632[3]), .I1(n396), .CO(n37572));
    SB_CARRY add_5775_4 (.CI(n38110), .I0(n14888[1]), .I1(n232), .CO(n38111));
    SB_LUT4 add_5775_3_lut (.I0(GND_net), .I1(n14888[0]), .I2(n159), .I3(n38109), 
            .O(n14167[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_3 (.CI(n38109), .I0(n14888[0]), .I1(n159), .CO(n38110));
    SB_LUT4 add_5948_5_lut (.I0(GND_net), .I1(n17632[2]), .I2(n323), .I3(n37570), 
            .O(n17268[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_5 (.CI(n37570), .I0(n17632[2]), .I1(n323), .CO(n37571));
    SB_LUT4 add_5775_2_lut (.I0(GND_net), .I1(n17), .I2(n86), .I3(GND_net), 
            .O(n14167[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5775_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5948_4_lut (.I0(GND_net), .I1(n17632[1]), .I2(n250), .I3(n37569), 
            .O(n17268[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_4 (.CI(n37569), .I0(n17632[1]), .I1(n250), .CO(n37570));
    SB_LUT4 add_5948_3_lut (.I0(GND_net), .I1(n17632[0]), .I2(n177), .I3(n37568), 
            .O(n17268[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5775_2 (.CI(GND_net), .I0(n17), .I1(n86), .CO(n38109));
    SB_CARRY add_5948_3 (.CI(n37568), .I0(n17632[0]), .I1(n177), .CO(n37569));
    SB_LUT4 add_5811_19_lut (.I0(GND_net), .I1(n15535[16]), .I2(GND_net), 
            .I3(n38108), .O(n14888[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5948_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n17268[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5948_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5948_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n37568));
    SB_LUT4 add_5811_18_lut (.I0(GND_net), .I1(n15535[15]), .I2(GND_net), 
            .I3(n38107), .O(n14888[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23989_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [18]), .I3(\Ki[1] ), 
            .O(n18948[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23989_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_5811_18 (.CI(n38107), .I0(n15535[15]), .I1(GND_net), 
            .CO(n38108));
    SB_LUT4 add_5973_13_lut (.I0(GND_net), .I1(n17944[10]), .I2(n910), 
            .I3(n37567), .O(n17632[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5973_12_lut (.I0(GND_net), .I1(n17944[9]), .I2(n837), 
            .I3(n37566), .O(n17632[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_12 (.CI(n37566), .I0(n17944[9]), .I1(n837), .CO(n37567));
    SB_LUT4 add_5973_11_lut (.I0(GND_net), .I1(n17944[8]), .I2(n764), 
            .I3(n37565), .O(n17632[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5811_17_lut (.I0(GND_net), .I1(n15535[14]), .I2(GND_net), 
            .I3(n38106), .O(n14888[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_17 (.CI(n38106), .I0(n15535[14]), .I1(GND_net), 
            .CO(n38107));
    SB_CARRY add_5973_11 (.CI(n37565), .I0(n17944[8]), .I1(n764), .CO(n37566));
    SB_LUT4 i23991_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [18]), .I3(\Ki[1] ), 
            .O(n37004));   // verilog/motorControl.v(34[25:36])
    defparam i23991_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_5973_10_lut (.I0(GND_net), .I1(n17944[7]), .I2(n691), 
            .I3(n37564), .O(n17632[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_10 (.CI(n37564), .I0(n17944[7]), .I1(n691), .CO(n37565));
    SB_LUT4 add_5973_9_lut (.I0(GND_net), .I1(n17944[6]), .I2(n618), .I3(n37563), 
            .O(n17632[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_9 (.CI(n37563), .I0(n17944[6]), .I1(n618), .CO(n37564));
    SB_LUT4 add_5973_8_lut (.I0(GND_net), .I1(n17944[5]), .I2(n545), .I3(n37562), 
            .O(n17632[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_8 (.CI(n37562), .I0(n17944[5]), .I1(n545), .CO(n37563));
    SB_LUT4 add_5973_7_lut (.I0(GND_net), .I1(n17944[4]), .I2(n472), .I3(n37561), 
            .O(n17632[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_7 (.CI(n37561), .I0(n17944[4]), .I1(n472), .CO(n37562));
    SB_LUT4 add_5973_6_lut (.I0(GND_net), .I1(n17944[3]), .I2(n399), .I3(n37560), 
            .O(n17632[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_6 (.CI(n37560), .I0(n17944[3]), .I1(n399), .CO(n37561));
    SB_LUT4 add_5811_16_lut (.I0(GND_net), .I1(n15535[13]), .I2(n1111), 
            .I3(n38105), .O(n14888[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5973_5_lut (.I0(GND_net), .I1(n17944[2]), .I2(n326), .I3(n37559), 
            .O(n17632[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_5 (.CI(n37559), .I0(n17944[2]), .I1(n326), .CO(n37560));
    SB_LUT4 add_5973_4_lut (.I0(GND_net), .I1(n17944[1]), .I2(n253), .I3(n37558), 
            .O(n17632[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_4 (.CI(n37558), .I0(n17944[1]), .I1(n253), .CO(n37559));
    SB_CARRY add_5811_16 (.CI(n38105), .I0(n15535[13]), .I1(n1111), .CO(n38106));
    SB_LUT4 add_5973_3_lut (.I0(GND_net), .I1(n17944[0]), .I2(n180), .I3(n37557), 
            .O(n17632[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5973_3 (.CI(n37557), .I0(n17944[0]), .I1(n180), .CO(n37558));
    SB_LUT4 add_5811_15_lut (.I0(GND_net), .I1(n15535[12]), .I2(n1038), 
            .I3(n38104), .O(n14888[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5973_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n17632[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5973_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_15 (.CI(n38104), .I0(n15535[12]), .I1(n1038), .CO(n38105));
    SB_CARRY add_5973_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n37557));
    SB_LUT4 add_5811_14_lut (.I0(GND_net), .I1(n15535[11]), .I2(n965), 
            .I3(n38103), .O(n14888[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_14 (.CI(n38103), .I0(n15535[11]), .I1(n965), .CO(n38104));
    SB_LUT4 add_6087_7_lut (.I0(GND_net), .I1(n44192), .I2(n490), .I3(n37556), 
            .O(n18912[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5811_13_lut (.I0(GND_net), .I1(n15535[10]), .I2(n892), 
            .I3(n38102), .O(n14888[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_6_lut (.I0(GND_net), .I1(n18983[3]), .I2(n417), .I3(n37555), 
            .O(n18912[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_6 (.CI(n37555), .I0(n18983[3]), .I1(n417), .CO(n37556));
    SB_LUT4 add_6087_5_lut (.I0(GND_net), .I1(n18983[2]), .I2(n344), .I3(n37554), 
            .O(n18912[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_13 (.CI(n38102), .I0(n15535[10]), .I1(n892), .CO(n38103));
    SB_CARRY add_6087_5 (.CI(n37554), .I0(n18983[2]), .I1(n344), .CO(n37555));
    SB_LUT4 add_6087_4_lut (.I0(GND_net), .I1(n18983[1]), .I2(n271), .I3(n37553), 
            .O(n18912[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_4 (.CI(n37553), .I0(n18983[1]), .I1(n271), .CO(n37554));
    SB_LUT4 add_6087_3_lut (.I0(GND_net), .I1(n18983[0]), .I2(n198), .I3(n37552), 
            .O(n18912[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_3 (.CI(n37552), .I0(n18983[0]), .I1(n198), .CO(n37553));
    SB_LUT4 add_5811_12_lut (.I0(GND_net), .I1(n15535[9]), .I2(n819), 
            .I3(n38101), .O(n14888[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_12 (.CI(n38101), .I0(n15535[9]), .I1(n819), .CO(n38102));
    SB_LUT4 add_711_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n3616[23]), .I3(n37329), .O(\PID_CONTROLLER.integral_23__N_3572 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6087_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n18912[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6087_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_711_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n3616[22]), .I3(n37328), .O(\PID_CONTROLLER.integral_23__N_3572 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6087_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n37552));
    SB_LUT4 add_5811_11_lut (.I0(GND_net), .I1(n15535[8]), .I2(n746), 
            .I3(n38100), .O(n14888[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5996_12_lut (.I0(GND_net), .I1(n18208[9]), .I2(n840_adj_4415), 
            .I3(n37539), .O(n17944[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5996_11_lut (.I0(GND_net), .I1(n18208[8]), .I2(n767_adj_4414), 
            .I3(n37538), .O(n17944[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_11 (.CI(n37538), .I0(n18208[8]), .I1(n767_adj_4414), 
            .CO(n37539));
    SB_LUT4 add_5996_10_lut (.I0(GND_net), .I1(n18208[7]), .I2(n694_adj_4413), 
            .I3(n37537), .O(n17944[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_10 (.CI(n37537), .I0(n18208[7]), .I1(n694_adj_4413), 
            .CO(n37538));
    SB_LUT4 add_5996_9_lut (.I0(GND_net), .I1(n18208[6]), .I2(n621_adj_4412), 
            .I3(n37536), .O(n17944[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_9 (.CI(n37536), .I0(n18208[6]), .I1(n621_adj_4412), 
            .CO(n37537));
    SB_LUT4 add_5996_8_lut (.I0(GND_net), .I1(n18208[5]), .I2(n548_adj_4411), 
            .I3(n37535), .O(n17944[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_8 (.CI(n37535), .I0(n18208[5]), .I1(n548_adj_4411), 
            .CO(n37536));
    SB_LUT4 add_5996_7_lut (.I0(GND_net), .I1(n18208[4]), .I2(n475_adj_4410), 
            .I3(n37534), .O(n17944[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_7 (.CI(n37534), .I0(n18208[4]), .I1(n475_adj_4410), 
            .CO(n37535));
    SB_LUT4 add_5996_6_lut (.I0(GND_net), .I1(n18208[3]), .I2(n402_adj_4409), 
            .I3(n37533), .O(n17944[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_6 (.CI(n37533), .I0(n18208[3]), .I1(n402_adj_4409), 
            .CO(n37534));
    SB_LUT4 add_5996_5_lut (.I0(GND_net), .I1(n18208[2]), .I2(n329_adj_4408), 
            .I3(n37532), .O(n17944[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_5 (.CI(n37532), .I0(n18208[2]), .I1(n329_adj_4408), 
            .CO(n37533));
    SB_LUT4 add_5996_4_lut (.I0(GND_net), .I1(n18208[1]), .I2(n256_adj_4407), 
            .I3(n37531), .O(n17944[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_4 (.CI(n37531), .I0(n18208[1]), .I1(n256_adj_4407), 
            .CO(n37532));
    SB_LUT4 add_5996_3_lut (.I0(GND_net), .I1(n18208[0]), .I2(n183_adj_4406), 
            .I3(n37530), .O(n17944[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_11 (.CI(n38100), .I0(n15535[8]), .I1(n746), .CO(n38101));
    SB_CARRY add_711_24 (.CI(n37328), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n3616[22]), .CO(n37329));
    SB_LUT4 add_711_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n3616[21]), .I3(n37327), .O(\PID_CONTROLLER.integral_23__N_3572 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_3 (.CI(n37530), .I0(n18208[0]), .I1(n183_adj_4406), 
            .CO(n37531));
    SB_LUT4 add_5996_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n17944[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5996_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5996_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n37530));
    SB_CARRY add_711_23 (.CI(n37327), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n3616[21]), .CO(n37328));
    SB_LUT4 add_6017_11_lut (.I0(GND_net), .I1(n18428[8]), .I2(n770), 
            .I3(n37529), .O(n18208[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6017_10_lut (.I0(GND_net), .I1(n18428[7]), .I2(n697), 
            .I3(n37528), .O(n18208[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6017_10 (.CI(n37528), .I0(n18428[7]), .I1(n697), .CO(n37529));
    SB_LUT4 add_6017_9_lut (.I0(GND_net), .I1(n18428[6]), .I2(n624), .I3(n37527), 
            .O(n18208[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_711_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n3616[20]), .I3(n37326), .O(\PID_CONTROLLER.integral_23__N_3572 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5811_10_lut (.I0(GND_net), .I1(n15535[7]), .I2(n673), 
            .I3(n38099), .O(n14888[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6017_9 (.CI(n37527), .I0(n18428[6]), .I1(n624), .CO(n37528));
    SB_CARRY add_711_22 (.CI(n37326), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n3616[20]), .CO(n37327));
    SB_LUT4 add_6017_8_lut (.I0(GND_net), .I1(n18428[5]), .I2(n551), .I3(n37526), 
            .O(n18208[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6017_8 (.CI(n37526), .I0(n18428[5]), .I1(n551), .CO(n37527));
    SB_LUT4 add_6017_7_lut (.I0(GND_net), .I1(n18428[4]), .I2(n478), .I3(n37525), 
            .O(n18208[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_10 (.CI(n38099), .I0(n15535[7]), .I1(n673), .CO(n38100));
    SB_CARRY add_6017_7 (.CI(n37525), .I0(n18428[4]), .I1(n478), .CO(n37526));
    SB_LUT4 add_6017_6_lut (.I0(GND_net), .I1(n18428[3]), .I2(n405), .I3(n37524), 
            .O(n18208[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6017_6 (.CI(n37524), .I0(n18428[3]), .I1(n405), .CO(n37525));
    SB_LUT4 add_711_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n3616[19]), .I3(n37325), .O(\PID_CONTROLLER.integral_23__N_3572 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5811_9_lut (.I0(GND_net), .I1(n15535[6]), .I2(n600), .I3(n38098), 
            .O(n14888[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6017_5_lut (.I0(GND_net), .I1(n18428[2]), .I2(n332), .I3(n37523), 
            .O(n18208[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_21 (.CI(n37325), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n3616[19]), .CO(n37326));
    SB_CARRY add_6017_5 (.CI(n37523), .I0(n18428[2]), .I1(n332), .CO(n37524));
    SB_LUT4 add_6017_4_lut (.I0(GND_net), .I1(n18428[1]), .I2(n259_adj_4401), 
            .I3(n37522), .O(n18208[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6017_4 (.CI(n37522), .I0(n18428[1]), .I1(n259_adj_4401), 
            .CO(n37523));
    SB_LUT4 add_6017_3_lut (.I0(GND_net), .I1(n18428[0]), .I2(n186), .I3(n37521), 
            .O(n18208[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6017_3 (.CI(n37521), .I0(n18428[0]), .I1(n186), .CO(n37522));
    SB_LUT4 add_6017_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n18208[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6017_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6017_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n37521));
    SB_CARRY add_5811_9 (.CI(n38098), .I0(n15535[6]), .I1(n600), .CO(n38099));
    SB_LUT4 add_5811_8_lut (.I0(GND_net), .I1(n15535[5]), .I2(n527), .I3(n38097), 
            .O(n14888[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6036_10_lut (.I0(GND_net), .I1(n18608[7]), .I2(n700), 
            .I3(n37520), .O(n18428[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6036_9_lut (.I0(GND_net), .I1(n18608[6]), .I2(n627), .I3(n37519), 
            .O(n18428[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6036_9 (.CI(n37519), .I0(n18608[6]), .I1(n627), .CO(n37520));
    SB_LUT4 add_711_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n3616[18]), .I3(n37324), .O(\PID_CONTROLLER.integral_23__N_3572 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6036_8_lut (.I0(GND_net), .I1(n18608[5]), .I2(n554), .I3(n37518), 
            .O(n18428[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6036_8 (.CI(n37518), .I0(n18608[5]), .I1(n554), .CO(n37519));
    SB_LUT4 add_6036_7_lut (.I0(GND_net), .I1(n18608[4]), .I2(n481), .I3(n37517), 
            .O(n18428[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_8 (.CI(n38097), .I0(n15535[5]), .I1(n527), .CO(n38098));
    SB_LUT4 add_5811_7_lut (.I0(GND_net), .I1(n15535[4]), .I2(n454), .I3(n38096), 
            .O(n14888[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6036_7 (.CI(n37517), .I0(n18608[4]), .I1(n481), .CO(n37518));
    SB_LUT4 add_6036_6_lut (.I0(GND_net), .I1(n18608[3]), .I2(n408), .I3(n37516), 
            .O(n18428[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_20 (.CI(n37324), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n3616[18]), .CO(n37325));
    SB_CARRY add_6036_6 (.CI(n37516), .I0(n18608[3]), .I1(n408), .CO(n37517));
    SB_LUT4 add_711_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n3616[17]), .I3(n37323), .O(\PID_CONTROLLER.integral_23__N_3572 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6036_5_lut (.I0(GND_net), .I1(n18608[2]), .I2(n335), .I3(n37515), 
            .O(n18428[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6036_5 (.CI(n37515), .I0(n18608[2]), .I1(n335), .CO(n37516));
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4771));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5811_7 (.CI(n38096), .I0(n15535[4]), .I1(n454), .CO(n38097));
    SB_LUT4 add_6036_4_lut (.I0(GND_net), .I1(n18608[1]), .I2(n262), .I3(n37514), 
            .O(n18428[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6036_4 (.CI(n37514), .I0(n18608[1]), .I1(n262), .CO(n37515));
    SB_LUT4 add_6036_3_lut (.I0(GND_net), .I1(n18608[0]), .I2(n189), .I3(n37513), 
            .O(n18428[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6036_3 (.CI(n37513), .I0(n18608[0]), .I1(n189), .CO(n37514));
    SB_LUT4 add_6036_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n18428[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6036_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6036_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n37513));
    SB_LUT4 add_6053_9_lut (.I0(GND_net), .I1(n18752[6]), .I2(n630), .I3(n37512), 
            .O(n18608[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6053_8_lut (.I0(GND_net), .I1(n18752[5]), .I2(n557_adj_4785), 
            .I3(n37511), .O(n18608[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6053_8 (.CI(n37511), .I0(n18752[5]), .I1(n557_adj_4785), 
            .CO(n37512));
    SB_LUT4 add_6053_7_lut (.I0(GND_net), .I1(n18752[4]), .I2(n484_adj_4786), 
            .I3(n37510), .O(n18608[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6053_7 (.CI(n37510), .I0(n18752[4]), .I1(n484_adj_4786), 
            .CO(n37511));
    SB_LUT4 add_6053_6_lut (.I0(GND_net), .I1(n18752[3]), .I2(n411_adj_4787), 
            .I3(n37509), .O(n18608[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6053_6 (.CI(n37509), .I0(n18752[3]), .I1(n411_adj_4787), 
            .CO(n37510));
    SB_LUT4 add_6053_5_lut (.I0(GND_net), .I1(n18752[2]), .I2(n338_adj_4788), 
            .I3(n37508), .O(n18608[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6053_5 (.CI(n37508), .I0(n18752[2]), .I1(n338_adj_4788), 
            .CO(n37509));
    SB_LUT4 add_6053_4_lut (.I0(GND_net), .I1(n18752[1]), .I2(n265_adj_4789), 
            .I3(n37507), .O(n18608[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6053_4 (.CI(n37507), .I0(n18752[1]), .I1(n265_adj_4789), 
            .CO(n37508));
    SB_LUT4 add_6053_3_lut (.I0(GND_net), .I1(n18752[0]), .I2(n192_adj_4790), 
            .I3(n37506), .O(n18608[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6053_3 (.CI(n37506), .I0(n18752[0]), .I1(n192_adj_4790), 
            .CO(n37507));
    SB_LUT4 add_6053_2_lut (.I0(GND_net), .I1(n50_adj_4791), .I2(n119_adj_4792), 
            .I3(GND_net), .O(n18608[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6053_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6053_2 (.CI(GND_net), .I0(n50_adj_4791), .I1(n119_adj_4792), 
            .CO(n37506));
    SB_LUT4 add_6068_8_lut (.I0(GND_net), .I1(n18864[5]), .I2(n560_adj_4793), 
            .I3(n37505), .O(n18752[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6068_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6068_7_lut (.I0(GND_net), .I1(n18864[4]), .I2(n487_adj_4794), 
            .I3(n37504), .O(n18752[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6068_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6068_7 (.CI(n37504), .I0(n18864[4]), .I1(n487_adj_4794), 
            .CO(n37505));
    SB_LUT4 add_6068_6_lut (.I0(GND_net), .I1(n18864[3]), .I2(n414_adj_4795), 
            .I3(n37503), .O(n18752[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6068_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6068_6 (.CI(n37503), .I0(n18864[3]), .I1(n414_adj_4795), 
            .CO(n37504));
    SB_LUT4 add_6068_5_lut (.I0(GND_net), .I1(n18864[2]), .I2(n341_adj_4796), 
            .I3(n37502), .O(n18752[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6068_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6068_5 (.CI(n37502), .I0(n18864[2]), .I1(n341_adj_4796), 
            .CO(n37503));
    SB_LUT4 add_6068_4_lut (.I0(GND_net), .I1(n18864[1]), .I2(n268_adj_4797), 
            .I3(n37501), .O(n18752[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6068_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6068_4 (.CI(n37501), .I0(n18864[1]), .I1(n268_adj_4797), 
            .CO(n37502));
    SB_LUT4 add_6068_3_lut (.I0(GND_net), .I1(n18864[0]), .I2(n195_adj_4798), 
            .I3(n37500), .O(n18752[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6068_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6068_3 (.CI(n37500), .I0(n18864[0]), .I1(n195_adj_4798), 
            .CO(n37501));
    SB_LUT4 add_6068_2_lut (.I0(GND_net), .I1(n53_adj_4799), .I2(n122_adj_4800), 
            .I3(GND_net), .O(n18752[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6068_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6068_2 (.CI(GND_net), .I0(n53_adj_4799), .I1(n122_adj_4800), 
            .CO(n37500));
    SB_LUT4 add_6081_7_lut (.I0(GND_net), .I1(n43558), .I2(n490_adj_4801), 
            .I3(n37499), .O(n18864[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6081_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6081_6_lut (.I0(GND_net), .I1(n18948[3]), .I2(n417_adj_4802), 
            .I3(n37498), .O(n18864[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6081_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6081_6 (.CI(n37498), .I0(n18948[3]), .I1(n417_adj_4802), 
            .CO(n37499));
    SB_LUT4 add_6081_5_lut (.I0(GND_net), .I1(n18948[2]), .I2(n344_adj_4803), 
            .I3(n37497), .O(n18864[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6081_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6081_5 (.CI(n37497), .I0(n18948[2]), .I1(n344_adj_4803), 
            .CO(n37498));
    SB_LUT4 add_6081_4_lut (.I0(GND_net), .I1(n18948[1]), .I2(n271_adj_4804), 
            .I3(n37496), .O(n18864[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6081_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6081_4 (.CI(n37496), .I0(n18948[1]), .I1(n271_adj_4804), 
            .CO(n37497));
    SB_LUT4 add_6081_3_lut (.I0(GND_net), .I1(n18948[0]), .I2(n198_adj_4805), 
            .I3(n37495), .O(n18864[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6081_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6081_3 (.CI(n37495), .I0(n18948[0]), .I1(n198_adj_4805), 
            .CO(n37496));
    SB_LUT4 add_6081_2_lut (.I0(GND_net), .I1(n56_adj_4806), .I2(n125_adj_4807), 
            .I3(GND_net), .O(n18864[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6081_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6081_2 (.CI(GND_net), .I0(n56_adj_4806), .I1(n125_adj_4807), 
            .CO(n37495));
    SB_LUT4 add_5811_6_lut (.I0(GND_net), .I1(n15535[3]), .I2(n381_adj_4808), 
            .I3(n38095), .O(n14888[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_6 (.CI(n38095), .I0(n15535[3]), .I1(n381_adj_4808), 
            .CO(n38096));
    SB_LUT4 add_5811_5_lut (.I0(GND_net), .I1(n15535[2]), .I2(n308_adj_4809), 
            .I3(n38094), .O(n14888[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_5 (.CI(n38094), .I0(n15535[2]), .I1(n308_adj_4809), 
            .CO(n38095));
    SB_CARRY add_711_19 (.CI(n37323), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n3616[17]), .CO(n37324));
    SB_LUT4 add_5811_4_lut (.I0(GND_net), .I1(n15535[1]), .I2(n235_adj_4810), 
            .I3(n38093), .O(n14888[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_711_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n3616[16]), .I3(n37322), .O(\PID_CONTROLLER.integral_23__N_3572 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_4 (.CI(n38093), .I0(n15535[1]), .I1(n235_adj_4810), 
            .CO(n38094));
    SB_LUT4 add_5811_3_lut (.I0(GND_net), .I1(n15535[0]), .I2(n162_adj_4811), 
            .I3(n38092), .O(n14888[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_18 (.CI(n37322), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n3616[16]), .CO(n37323));
    SB_CARRY add_5811_3 (.CI(n38092), .I0(n15535[0]), .I1(n162_adj_4811), 
            .CO(n38093));
    SB_LUT4 add_5811_2_lut (.I0(GND_net), .I1(n20_adj_4812), .I2(n89_adj_4813), 
            .I3(GND_net), .O(n14888[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5811_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_711_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n3616[15]), .I3(n37321), .O(\PID_CONTROLLER.integral_23__N_3572 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5811_2 (.CI(GND_net), .I0(n20_adj_4812), .I1(n89_adj_4813), 
            .CO(n38092));
    SB_CARRY add_711_17 (.CI(n37321), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n3616[15]), .CO(n37322));
    SB_LUT4 add_711_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n3616[14]), .I3(n37320), .O(\PID_CONTROLLER.integral_23__N_3572 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_16 (.CI(n37320), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n3616[14]), .CO(n37321));
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4762));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_711_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n3616[13]), .I3(n37319), .O(\PID_CONTROLLER.integral_23__N_3572 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_15 (.CI(n37319), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n3616[13]), .CO(n37320));
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_711_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n3616[12]), .I3(n37318), .O(\PID_CONTROLLER.integral_23__N_3572 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4760));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_711_14 (.CI(n37318), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n3616[12]), .CO(n37319));
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4759));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4758));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4757));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[23]), 
            .I3(n37449), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_711_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n3616[11]), .I3(n37317), .O(\PID_CONTROLLER.integral_23__N_3572 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[22]), 
            .I3(n37448), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n37448), .I0(GND_net), .I1(n1_adj_4822[22]), 
            .CO(n37449));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[21]), 
            .I3(n37447), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n37447), .I0(GND_net), .I1(n1_adj_4822[21]), 
            .CO(n37448));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[20]), 
            .I3(n37446), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4756));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n37446), .I0(GND_net), .I1(n1_adj_4822[20]), 
            .CO(n37447));
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[19]), 
            .I3(n37445), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4754));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4753));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n37445), .I0(GND_net), .I1(n1_adj_4822[19]), 
            .CO(n37446));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[18]), 
            .I3(n37444), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n37444), .I0(GND_net), .I1(n1_adj_4822[18]), 
            .CO(n37445));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[17]), 
            .I3(n37443), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n37443), .I0(GND_net), .I1(n1_adj_4822[17]), 
            .CO(n37444));
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[16]), 
            .I3(n37442), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n37442), .I0(GND_net), .I1(n1_adj_4822[16]), 
            .CO(n37443));
    SB_CARRY add_711_13 (.CI(n37317), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n3616[11]), .CO(n37318));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[15]), 
            .I3(n37441), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n37441), .I0(GND_net), .I1(n1_adj_4822[15]), 
            .CO(n37442));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[14]), 
            .I3(n37440), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n37440), .I0(GND_net), .I1(n1_adj_4822[14]), 
            .CO(n37441));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[13]), 
            .I3(n37439), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n37439), .I0(GND_net), .I1(n1_adj_4822[13]), 
            .CO(n37440));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[12]), 
            .I3(n37438), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n37438), .I0(GND_net), .I1(n1_adj_4822[12]), 
            .CO(n37439));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[11]), 
            .I3(n37437), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n37437), .I0(GND_net), .I1(n1_adj_4822[11]), 
            .CO(n37438));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[10]), 
            .I3(n37436), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n37436), .I0(GND_net), .I1(n1_adj_4822[10]), 
            .CO(n37437));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[9]), 
            .I3(n37435), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n37435), .I0(GND_net), .I1(n1_adj_4822[9]), 
            .CO(n37436));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[8]), 
            .I3(n37434), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n37434), .I0(GND_net), .I1(n1_adj_4822[8]), 
            .CO(n37435));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[7]), 
            .I3(n37433), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n37433), .I0(GND_net), .I1(n1_adj_4822[7]), 
            .CO(n37434));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[6]), 
            .I3(n37432), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n37432), .I0(GND_net), .I1(n1_adj_4822[6]), 
            .CO(n37433));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[5]), 
            .I3(n37431), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n37431), .I0(GND_net), .I1(n1_adj_4822[5]), 
            .CO(n37432));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[4]), 
            .I3(n37430), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n37430), .I0(GND_net), .I1(n1_adj_4822[4]), 
            .CO(n37431));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[3]), 
            .I3(n37429), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n37429), .I0(GND_net), .I1(n1_adj_4822[3]), 
            .CO(n37430));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[2]), 
            .I3(n37428), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n37428), .I0(GND_net), .I1(n1_adj_4822[2]), 
            .CO(n37429));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[1]), 
            .I3(n37427), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n37427), .I0(GND_net), .I1(n1_adj_4822[1]), 
            .CO(n37428));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4822[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4822[0]), 
            .CO(n37427));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4821[23]), 
            .I3(n37426), .O(\PID_CONTROLLER.integral_23__N_3623 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_711_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n3616[10]), .I3(n37316), .O(\PID_CONTROLLER.integral_23__N_3572 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4821[22]), .I3(n37425), .O(n45_adj_4575)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n37425), .I0(GND_net), .I1(n1_adj_4821[22]), 
            .CO(n37426));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4821[21]), .I3(n37424), .O(n43_adj_4572)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n37424), .I0(GND_net), .I1(n1_adj_4821[21]), 
            .CO(n37425));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4821[20]), .I3(n37423), .O(n41_adj_4620)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n37423), .I0(GND_net), .I1(n1_adj_4821[20]), 
            .CO(n37424));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4821[19]), .I3(n37422), .O(n39_adj_4611)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n37422), .I0(GND_net), .I1(n1_adj_4821[19]), 
            .CO(n37423));
    SB_CARRY add_711_12 (.CI(n37316), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n3616[10]), .CO(n37317));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4821[18]), .I3(n37421), .O(n37_adj_4583)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n37421), .I0(GND_net), .I1(n1_adj_4821[18]), 
            .CO(n37422));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4821[17]), .I3(n37420), .O(n35_adj_4584)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n37420), .I0(GND_net), .I1(n1_adj_4821[17]), 
            .CO(n37421));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4821[16]), .I3(n37419), .O(n33_adj_4585)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n37419), .I0(GND_net), .I1(n1_adj_4821[16]), 
            .CO(n37420));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4821[15]), .I3(n37418), .O(n31_adj_4581)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n37418), .I0(GND_net), .I1(n1_adj_4821[15]), 
            .CO(n37419));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4821[14]), .I3(n37417), .O(n29_adj_4582)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n37417), .I0(GND_net), .I1(n1_adj_4821[14]), 
            .CO(n37418));
    SB_LUT4 add_711_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n3616[9]), .I3(n37315), .O(\PID_CONTROLLER.integral_23__N_3572 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4821[13]), .I3(n37416), .O(n27_adj_4564)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n37416), .I0(GND_net), .I1(n1_adj_4821[13]), 
            .CO(n37417));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4821[12]), .I3(n37415), .O(n25_adj_4579)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n37415), .I0(GND_net), .I1(n1_adj_4821[12]), 
            .CO(n37416));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4821[11]), .I3(n37414), .O(n23_adj_4580)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n37414), .I0(GND_net), .I1(n1_adj_4821[11]), 
            .CO(n37415));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4821[10]), .I3(n37413), .O(n21_adj_4568)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n37413), .I0(GND_net), .I1(n1_adj_4821[10]), 
            .CO(n37414));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4821[9]), .I3(n37412), .O(n19_adj_4569)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n37412), .I0(GND_net), .I1(n1_adj_4821[9]), 
            .CO(n37413));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4821[8]), .I3(n37411), .O(n17_adj_4570)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n37411), .I0(GND_net), .I1(n1_adj_4821[8]), 
            .CO(n37412));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4821[7]), .I3(n37410), .O(n15_adj_4565)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n37410), .I0(GND_net), .I1(n1_adj_4821[7]), 
            .CO(n37411));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4821[6]), .I3(n37409), .O(n13_adj_4566)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n37409), .I0(GND_net), .I1(n1_adj_4821[6]), 
            .CO(n37410));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4821[5]), .I3(n37408), .O(n11_adj_4567)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n37408), .I0(GND_net), .I1(n1_adj_4821[5]), 
            .CO(n37409));
    SB_CARRY add_711_11 (.CI(n37315), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n3616[9]), .CO(n37316));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4821[4]), .I3(n37407), .O(n9_adj_4571)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n37407), .I0(GND_net), .I1(n1_adj_4821[4]), 
            .CO(n37408));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4821[3]), .I3(n37406), .O(n7_adj_4577)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n37406), .I0(GND_net), .I1(n1_adj_4821[3]), 
            .CO(n37407));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4821[2]), .I3(n37405), .O(n5_adj_4578)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n37405), .I0(GND_net), .I1(n1_adj_4821[2]), 
            .CO(n37406));
    SB_LUT4 add_711_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n3616[8]), .I3(n37314), .O(\PID_CONTROLLER.integral_23__N_3572 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4821[1]), .I3(n37404), .O(n3_adj_4596)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n37404), .I0(GND_net), .I1(n1_adj_4821[1]), 
            .CO(n37405));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4821[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3623 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4821[0]), 
            .CO(n37404));
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n37403), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n37402), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n37402), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n37403));
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n37401), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_711_10 (.CI(n37314), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n3616[8]), .CO(n37315));
    SB_CARRY sub_3_add_2_23 (.CI(n37401), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n37402));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n37400), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_22 (.CI(n37400), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n37401));
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n37399), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n37399), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n37400));
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n37398), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n37398), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n37399));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n37397), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_711_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n3616[7]), .I3(n37313), .O(\PID_CONTROLLER.integral_23__N_3572 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_711_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n37397), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n37398));
    SB_CARRY add_711_9 (.CI(n37313), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n3616[7]), .CO(n37314));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n37396), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4750));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4744));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4742));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4741));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4740));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4736));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4735));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4733));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32902_3_lut_4_lut (.I0(duty_23__N_3672[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3672[2]), .O(n47855));   // verilog/motorControl.v(38[19:35])
    defparam i32902_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3672[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4466));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i32937_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3672[3]), 
            .I2(duty_23__N_3672[2]), .I3(PWMLimit[2]), .O(n47890));   // verilog/motorControl.v(36[10:25])
    defparam i32937_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_832_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3672[3]), 
            .I2(duty_23__N_3672[2]), .I3(GND_net), .O(n6_adj_4436));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4732));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4730));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4728));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4727));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4726));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4725));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4723));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4722));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4721));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4720));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4719));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4711));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4710));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4708));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4707));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20636_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20636_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20635_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20635_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20634_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20634_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4595));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i20633_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20633_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4812));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4811));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20632_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20632_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4696));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4695));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34295_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49248));   // verilog/motorControl.v(29[14] 48[8])
    defparam i34295_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4809));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4684));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4681));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4677));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24103_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4814), 
            .I3(n19032[1]), .O(n6_adj_4416));   // verilog/motorControl.v(34[16:22])
    defparam i24103_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4675));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1519 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n19032[1]), 
            .I3(n4_adj_4814), .O(n18983[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1519.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4674));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1520 (.I0(\Kp[2] ), .I1(n1[19]), .I2(n19063[0]), 
            .I3(n37072), .O(n19032[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1520.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4672));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4671));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4669));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4667));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4666));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4665));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24064_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n37072), 
            .I3(n19063[0]), .O(n4_adj_4417));   // verilog/motorControl.v(34[16:22])
    defparam i24064_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4657));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24051_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n19032[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24051_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24053_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n37072));   // verilog/motorControl.v(34[16:22])
    defparam i24053_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4642));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4641));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4640));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4639));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4638));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4808));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4637));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4636));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24041_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n37047), 
            .I3(n19080[0]), .O(n4_adj_4423));   // verilog/motorControl.v(34[16:22])
    defparam i24041_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4635));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1521 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n19080[0]), 
            .I3(n37047), .O(n19063[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1521.LUT_INIT = 16'h8778;
    SB_LUT4 i24030_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n37047));   // verilog/motorControl.v(34[16:22])
    defparam i24030_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4633));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24028_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n19063[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24028_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4632));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4806));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4805));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4631));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4628));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4626));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4625));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4803));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1522 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n19032[0]), 
            .I3(n37106), .O(n18983[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1522.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4802));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1523 (.I0(n6_adj_4782), .I1(\Ki[4] ), .I2(n19008[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [18]), .O(n18948[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1523.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4614));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32868_2_lut_4_lut (.I0(duty_23__N_3672[21]), .I1(n257[21]), 
            .I2(duty_23__N_3672[9]), .I3(n257[9]), .O(n47821));
    defparam i32868_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32879_2_lut_4_lut (.I0(duty_23__N_3672[16]), .I1(n257[16]), 
            .I2(duty_23__N_3672[7]), .I3(n257[7]), .O(n47832));
    defparam i32879_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i24095_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n37106), 
            .I3(n19032[0]), .O(n4_adj_4814));   // verilog/motorControl.v(34[16:22])
    defparam i24095_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i32905_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3672[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3672[9]), .O(n47858));
    defparam i32905_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32915_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3672[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3672[7]), .O(n47868));
    defparam i32915_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i24082_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n18983[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24082_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24084_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n37106));   // verilog/motorControl.v(34[16:22])
    defparam i24084_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i23905_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [21]), .O(n19072[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23905_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4607));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1524 (.I0(n4_adj_4779), .I1(\Ki[3] ), .I2(n19048[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [19]), .O(n19008[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1524.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4801));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1525 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [20]), .O(n12_adj_4815));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1525.LUT_INIT = 16'h9c50;
    SB_LUT4 i24018_4_lut (.I0(n19008[2]), .I1(\Ki[4] ), .I2(n6_adj_4782), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [18]), .O(n8_adj_4816));   // verilog/motorControl.v(34[25:36])
    defparam i24018_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3672[1]), .I1(n257[1]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1526 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [21]), .O(n11_adj_4817));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut_adj_1526.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23979_4_lut (.I0(n19048[1]), .I1(\Ki[3] ), .I2(n4_adj_4779), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [19]), .O(n6_adj_4818));   // verilog/motorControl.v(34[25:36])
    defparam i23979_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3647[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3672[2]), .I1(n257[2]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23907_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [21]), .O(n36913));   // verilog/motorControl.v(34[25:36])
    defparam i23907_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1527 (.I0(n6_adj_4818), .I1(n11_adj_4817), .I2(n8_adj_4816), 
            .I3(n12_adj_4815), .O(n18_adj_4819));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1528 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [22]), .O(n13_adj_4820));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut_adj_1528.LUT_INIT = 16'h6ca0;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3647[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1529 (.I0(n13_adj_4820), .I1(n18_adj_4819), .I2(n36913), 
            .I3(n4_adj_4778), .O(n43558));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3672[3]), .I1(n257[3]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3647[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3672[4]), .I1(n257[4]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3647[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3672[5]), .I1(n257[5]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3647[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3672[6]), .I1(n257[6]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3647[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3672[7]), .I1(n257[7]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3647[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3672[8]), .I1(n257[8]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3647[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3672[9]), .I1(n257[9]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4800));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3647[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4799));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3672[10]), .I1(n257[10]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3647[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3672[11]), .I1(n257[11]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3647[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3672[12]), .I1(n257[12]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4798));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4797));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4796));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3647[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4795));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4794));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3672[13]), .I1(n257[13]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3647[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4793));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4792));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3672[14]), .I1(n257[14]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3647[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3672[15]), .I1(n257[15]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4791));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4790));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3647[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3672[16]), .I1(n257[16]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3647[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3672[17]), .I1(n257[17]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4789));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4788));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4787));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3647[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3672[18]), .I1(n257[18]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3647[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3672[19]), .I1(n257[19]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3647[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4786));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4785));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (\a_new[1] , ENCODER1_B_N_keep, n1188, 
            ENCODER1_A_N_keep, b_prev, n28216, n1193, direction_N_3807, 
            encoder1_position, GND_net, VCC_net) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    input ENCODER1_B_N_keep;
    input n1188;
    input ENCODER1_A_N_keep;
    output b_prev;
    input n28216;
    output n1193;
    output direction_N_3807;
    output [31:0]encoder1_position;
    input GND_net;
    input VCC_net;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire a_prev_N_3813, debounce_cnt, n28217;
    wire [31:0]n133;
    
    wire n28196, a_prev, direction_N_3806, n38597, n38596, n38595, 
        n38594, n38593, n38592, n38591, n38590, n38589, n38588, 
        n38587, n38586, n38585, n38584, n38583, n38582, n38581, 
        n38580, n38579, n38578, n38577, n38576, n38575, n38574, 
        n38573, n38572, n38571, n38570, n38569, n38568, n38567, 
        direction_N_3810;
    
    SB_LUT4 i33563_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i33563_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1188), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1188), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1188), .D(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1188), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1188), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1188), .D(n28217));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1193), .C(n1188), .D(n28216));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_1549__i0 (.Q(encoder1_position[0]), .C(n1188), .E(direction_N_3807), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1188), .D(n28196));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i15158_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(b_new[1]), 
            .I3(b_prev), .O(n28217));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15158_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15137_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n28196));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15137_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE position_1549__i1 (.Q(encoder1_position[1]), .C(n1188), .E(direction_N_3807), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i2 (.Q(encoder1_position[2]), .C(n1188), .E(direction_N_3807), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i3 (.Q(encoder1_position[3]), .C(n1188), .E(direction_N_3807), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i4 (.Q(encoder1_position[4]), .C(n1188), .E(direction_N_3807), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i5 (.Q(encoder1_position[5]), .C(n1188), .E(direction_N_3807), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i6 (.Q(encoder1_position[6]), .C(n1188), .E(direction_N_3807), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i7 (.Q(encoder1_position[7]), .C(n1188), .E(direction_N_3807), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i8 (.Q(encoder1_position[8]), .C(n1188), .E(direction_N_3807), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i9 (.Q(encoder1_position[9]), .C(n1188), .E(direction_N_3807), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i10 (.Q(encoder1_position[10]), .C(n1188), .E(direction_N_3807), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i11 (.Q(encoder1_position[11]), .C(n1188), .E(direction_N_3807), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i12 (.Q(encoder1_position[12]), .C(n1188), .E(direction_N_3807), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i13 (.Q(encoder1_position[13]), .C(n1188), .E(direction_N_3807), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i14 (.Q(encoder1_position[14]), .C(n1188), .E(direction_N_3807), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i15 (.Q(encoder1_position[15]), .C(n1188), .E(direction_N_3807), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i16 (.Q(encoder1_position[16]), .C(n1188), .E(direction_N_3807), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i17 (.Q(encoder1_position[17]), .C(n1188), .E(direction_N_3807), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i18 (.Q(encoder1_position[18]), .C(n1188), .E(direction_N_3807), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i19 (.Q(encoder1_position[19]), .C(n1188), .E(direction_N_3807), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i20 (.Q(encoder1_position[20]), .C(n1188), .E(direction_N_3807), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i21 (.Q(encoder1_position[21]), .C(n1188), .E(direction_N_3807), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i22 (.Q(encoder1_position[22]), .C(n1188), .E(direction_N_3807), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i23 (.Q(encoder1_position[23]), .C(n1188), .E(direction_N_3807), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i24 (.Q(encoder1_position[24]), .C(n1188), .E(direction_N_3807), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i25 (.Q(encoder1_position[25]), .C(n1188), .E(direction_N_3807), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i26 (.Q(encoder1_position[26]), .C(n1188), .E(direction_N_3807), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i27 (.Q(encoder1_position[27]), .C(n1188), .E(direction_N_3807), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i28 (.Q(encoder1_position[28]), .C(n1188), .E(direction_N_3807), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i29 (.Q(encoder1_position[29]), .C(n1188), .E(direction_N_3807), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i30 (.Q(encoder1_position[30]), .C(n1188), .E(direction_N_3807), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1549__i31 (.Q(encoder1_position[31]), .C(n1188), .E(direction_N_3807), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_1549_add_4_33_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[31]), .I3(n38597), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1549_add_4_32_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[30]), .I3(n38596), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_32 (.CI(n38596), .I0(direction_N_3806), 
            .I1(encoder1_position[30]), .CO(n38597));
    SB_LUT4 position_1549_add_4_31_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[29]), .I3(n38595), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_31 (.CI(n38595), .I0(direction_N_3806), 
            .I1(encoder1_position[29]), .CO(n38596));
    SB_LUT4 position_1549_add_4_30_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[28]), .I3(n38594), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_30 (.CI(n38594), .I0(direction_N_3806), 
            .I1(encoder1_position[28]), .CO(n38595));
    SB_LUT4 position_1549_add_4_29_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[27]), .I3(n38593), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_29 (.CI(n38593), .I0(direction_N_3806), 
            .I1(encoder1_position[27]), .CO(n38594));
    SB_LUT4 position_1549_add_4_28_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[26]), .I3(n38592), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_28 (.CI(n38592), .I0(direction_N_3806), 
            .I1(encoder1_position[26]), .CO(n38593));
    SB_LUT4 position_1549_add_4_27_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[25]), .I3(n38591), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_27 (.CI(n38591), .I0(direction_N_3806), 
            .I1(encoder1_position[25]), .CO(n38592));
    SB_LUT4 position_1549_add_4_26_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[24]), .I3(n38590), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_26 (.CI(n38590), .I0(direction_N_3806), 
            .I1(encoder1_position[24]), .CO(n38591));
    SB_LUT4 position_1549_add_4_25_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[23]), .I3(n38589), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_25 (.CI(n38589), .I0(direction_N_3806), 
            .I1(encoder1_position[23]), .CO(n38590));
    SB_LUT4 position_1549_add_4_24_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[22]), .I3(n38588), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_24 (.CI(n38588), .I0(direction_N_3806), 
            .I1(encoder1_position[22]), .CO(n38589));
    SB_LUT4 position_1549_add_4_23_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[21]), .I3(n38587), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_23 (.CI(n38587), .I0(direction_N_3806), 
            .I1(encoder1_position[21]), .CO(n38588));
    SB_LUT4 position_1549_add_4_22_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[20]), .I3(n38586), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_22 (.CI(n38586), .I0(direction_N_3806), 
            .I1(encoder1_position[20]), .CO(n38587));
    SB_LUT4 position_1549_add_4_21_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[19]), .I3(n38585), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_21 (.CI(n38585), .I0(direction_N_3806), 
            .I1(encoder1_position[19]), .CO(n38586));
    SB_LUT4 position_1549_add_4_20_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[18]), .I3(n38584), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_20 (.CI(n38584), .I0(direction_N_3806), 
            .I1(encoder1_position[18]), .CO(n38585));
    SB_LUT4 position_1549_add_4_19_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[17]), .I3(n38583), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_19 (.CI(n38583), .I0(direction_N_3806), 
            .I1(encoder1_position[17]), .CO(n38584));
    SB_LUT4 position_1549_add_4_18_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[16]), .I3(n38582), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_18 (.CI(n38582), .I0(direction_N_3806), 
            .I1(encoder1_position[16]), .CO(n38583));
    SB_LUT4 position_1549_add_4_17_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[15]), .I3(n38581), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_17 (.CI(n38581), .I0(direction_N_3806), 
            .I1(encoder1_position[15]), .CO(n38582));
    SB_LUT4 position_1549_add_4_16_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[14]), .I3(n38580), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_16 (.CI(n38580), .I0(direction_N_3806), 
            .I1(encoder1_position[14]), .CO(n38581));
    SB_LUT4 position_1549_add_4_15_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[13]), .I3(n38579), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_15 (.CI(n38579), .I0(direction_N_3806), 
            .I1(encoder1_position[13]), .CO(n38580));
    SB_LUT4 position_1549_add_4_14_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[12]), .I3(n38578), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_14 (.CI(n38578), .I0(direction_N_3806), 
            .I1(encoder1_position[12]), .CO(n38579));
    SB_LUT4 position_1549_add_4_13_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[11]), .I3(n38577), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_13 (.CI(n38577), .I0(direction_N_3806), 
            .I1(encoder1_position[11]), .CO(n38578));
    SB_LUT4 position_1549_add_4_12_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[10]), .I3(n38576), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_12 (.CI(n38576), .I0(direction_N_3806), 
            .I1(encoder1_position[10]), .CO(n38577));
    SB_LUT4 position_1549_add_4_11_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[9]), .I3(n38575), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_11 (.CI(n38575), .I0(direction_N_3806), 
            .I1(encoder1_position[9]), .CO(n38576));
    SB_LUT4 position_1549_add_4_10_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[8]), .I3(n38574), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_10 (.CI(n38574), .I0(direction_N_3806), 
            .I1(encoder1_position[8]), .CO(n38575));
    SB_LUT4 position_1549_add_4_9_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[7]), .I3(n38573), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_9 (.CI(n38573), .I0(direction_N_3806), 
            .I1(encoder1_position[7]), .CO(n38574));
    SB_LUT4 position_1549_add_4_8_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[6]), .I3(n38572), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_8 (.CI(n38572), .I0(direction_N_3806), 
            .I1(encoder1_position[6]), .CO(n38573));
    SB_LUT4 position_1549_add_4_7_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[5]), .I3(n38571), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_7 (.CI(n38571), .I0(direction_N_3806), 
            .I1(encoder1_position[5]), .CO(n38572));
    SB_LUT4 position_1549_add_4_6_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[4]), .I3(n38570), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_6 (.CI(n38570), .I0(direction_N_3806), 
            .I1(encoder1_position[4]), .CO(n38571));
    SB_LUT4 position_1549_add_4_5_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[3]), .I3(n38569), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_5 (.CI(n38569), .I0(direction_N_3806), 
            .I1(encoder1_position[3]), .CO(n38570));
    SB_LUT4 position_1549_add_4_4_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[2]), .I3(n38568), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_4 (.CI(n38568), .I0(direction_N_3806), 
            .I1(encoder1_position[2]), .CO(n38569));
    SB_LUT4 position_1549_add_4_3_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[1]), .I3(n38567), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_3 (.CI(n38567), .I0(direction_N_3806), 
            .I1(encoder1_position[1]), .CO(n38568));
    SB_LUT4 position_1549_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1549_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1549_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n38567));
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3810));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3810), 
            .I3(\a_new[1] ), .O(direction_N_3807));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3806));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module coms
//

module coms (CLK_c, n28292, control_mode, n28291, n28290, n28289, 
            n28288, GND_net, \data_in_frame[3] , n28287, \data_in_frame[2] , 
            n28286, \data_in_frame[1] , n28285, PWMLimit, n28284, 
            \data_in_frame[8] , \data_in_frame[6] , n23943, \data_in_frame[13] , 
            \data_in_frame[12] , \data_in_frame[10] , byte_transmit_counter, 
            n28283, n28282, n28281, n28280, \data_in_frame[0] , \data_in_frame[5] , 
            \data_in_frame[4] , n28279, n28278, n28277, n28276, rx_data_ready, 
            setpoint, \data_in_frame[11] , n28275, n28274, \data_in[3] , 
            \data_in[1] , \data_in[0] , \data_in[2] , n28273, n28272, 
            \data_in_frame[9] , \byte_transmit_counter[0] , \data_out_frame[8] , 
            \data_out_frame[9] , n28271, \data_out_frame[10] , \data_out_frame[11] , 
            n28270, n28269, \data_out_frame[14] , \data_out_frame[15] , 
            \data_out_frame[12] , \data_out_frame[13] , n28268, n28267, 
            n28266, n28265, n28264, n28263, \data_out_frame[16] , 
            \data_out_frame[17] , \data_out_frame[18] , \data_out_frame[19] , 
            \data_out_frame[23] , \data_out_frame[20] , DE_c, tx_active, 
            \data_out_frame[6] , \data_out_frame[7] , \data_out_frame[4] , 
            \data_out_frame[5] , n49368, n46660, ID, n43603, n42551, 
            n27752, \data_out_frame[24] , n47614, \data_out_frame[25] , 
            n42541, n42790, LED_c, n49422, n28189, n43610, n27554, 
            n28188, n42897, \data_out_frame[18][6] , n40598, n28187, 
            n28186, neopxl_color, n28185, \Ki[0] , n28184, \Kp[0] , 
            n28183, n28738, IntegralLimit, n28737, n28736, n28735, 
            n28734, n28733, n28732, n28731, n28730, n28729, n28728, 
            n28727, n28726, n28725, n28724, n28723, n28722, n28721, 
            n28720, n28719, n28718, n28717, n28716, n28715, n28714, 
            n28713, n28712, n28711, n28710, n28709, n28708, n28707, 
            n28706, n28705, n28704, n28703, n28702, n28701, n28700, 
            n28698, n28697, n28696, n28695, n28694, n28693, n28692, 
            n28691, n28690, n28689, n28688, n28687, n28686, n28685, 
            n28684, n28683, \Kp[1] , n28682, \Kp[2] , n28681, \Kp[3] , 
            n28680, \Kp[4] , n28679, \Kp[5] , n28678, \Kp[6] , n28677, 
            \Kp[7] , n28676, \Kp[8] , n28675, \Kp[9] , n28674, \Kp[10] , 
            n28673, \Kp[11] , n28672, \Kp[12] , n28671, \Kp[13] , 
            n28670, \Kp[14] , n28669, \Kp[15] , n28668, \Ki[1] , 
            n28667, \Ki[2] , n28666, \Ki[3] , n28665, \Ki[4] , n28664, 
            \Ki[5] , n28663, \Ki[6] , n28662, \Ki[7] , n28661, \Ki[8] , 
            n28660, \Ki[9] , n28659, \Ki[10] , n28658, \Ki[11] , 
            n28657, \Ki[12] , n28656, \Ki[13] , n28655, \Ki[14] , 
            n28654, \Ki[15] , n28653, n28652, n28651, n28650, n28649, 
            n28648, n28647, n28646, n28645, n28644, n28643, n28642, 
            n28641, n28640, n28639, n28638, n28637, n28636, n28635, 
            n28634, n28633, n28632, n28631, n28630, n28629, n28628, 
            n28627, n28626, n28625, n28624, n28623, n28622, n28621, 
            n28620, n28619, n28618, n28617, n28616, n28615, n28614, 
            n28613, n28612, n28611, n28610, n28609, n28608, n28607, 
            n28606, n28605, n28604, n28603, n28602, n28601, n28600, 
            n28599, n28598, n28597, n28596, n28595, n28594, n28593, 
            n28592, n28591, n28590, n28589, n28588, n28587, n28586, 
            n28585, n28584, n28583, n28582, rx_data, n28581, n28580, 
            n28579, n28578, n28577, n28576, n28575, n28574, n28573, 
            n28572, n28571, n28570, n28569, n28568, n28567, n28566, 
            n28565, n28564, n28563, n28562, n28561, n28560, n28559, 
            n28558, n28557, n28556, n28555, n28554, n28553, n28552, 
            n28551, n28550, n28549, n28548, n28547, n28546, n28545, 
            n28544, n28543, n28542, n28541, n28539, n28538, n28537, 
            n28536, n28535, n28534, n28533, n28532, n28531, n28530, 
            n28529, n28528, n28527, n28526, n28525, n28524, n28523, 
            n28522, n28521, n28520, n28519, n28518, n28517, n28516, 
            n28515, n28514, n28513, n28512, n28511, n28510, n28509, 
            n28508, n28507, n28164, n28506, n28505, n28504, n28503, 
            n28502, n28501, n28500, n28499, n28498, n28497, n28496, 
            n28495, n28494, n28493, n28492, n28491, n28490, n28489, 
            n28488, n28487, n28486, n28485, n28484, n28483, n28482, 
            n28481, n28480, n28479, n28478, n28477, n28476, n28475, 
            n28474, n28473, n28472, n28471, n28470, n28469, n28468, 
            n28467, n28466, n28465, n28464, n28405, n28403, n28402, 
            n28401, n28400, n28399, n28398, n28397, n4, \state[0] , 
            \state[2] , \state[3] , n6014, \displacement[17] , n27753, 
            n42230, n42229, \r_SM_Main_2__N_3513[1] , r_SM_Main, \r_Bit_Index[0] , 
            n42123, n27820, tx_o, n19247, n49552, n28192, n4_adj_6, 
            n28212, VCC_net, tx_enable, n4_adj_7, r_SM_Main_adj_14, 
            r_Rx_Data, \r_SM_Main_2__N_3442[2] , n27824, \r_Bit_Index[0]_adj_11 , 
            n26628, n33696, RX_N_10, n42126, n41813, n28224, n28182, 
            n28181, n28180, n27784, n28179, n28178, n28177, n28176, 
            n42185, n28215, n26633, n4_adj_12, n4_adj_13) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    input n28292;
    output [7:0]control_mode;
    input n28291;
    input n28290;
    input n28289;
    input n28288;
    input GND_net;
    output [7:0]\data_in_frame[3] ;
    input n28287;
    output [7:0]\data_in_frame[2] ;
    input n28286;
    output [7:0]\data_in_frame[1] ;
    input n28285;
    output [23:0]PWMLimit;
    input n28284;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[6] ;
    output n23943;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]byte_transmit_counter;
    input n28283;
    input n28282;
    input n28281;
    input n28280;
    output [7:0]\data_in_frame[0] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[4] ;
    input n28279;
    input n28278;
    input n28277;
    input n28276;
    output rx_data_ready;
    output [23:0]setpoint;
    output [7:0]\data_in_frame[11] ;
    input n28275;
    input n28274;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[2] ;
    input n28273;
    input n28272;
    output [7:0]\data_in_frame[9] ;
    output \byte_transmit_counter[0] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[9] ;
    input n28271;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    input n28270;
    input n28269;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    input n28268;
    input n28267;
    input n28266;
    input n28265;
    input n28264;
    input n28263;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[20] ;
    output DE_c;
    output tx_active;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    input n49368;
    input n46660;
    input [7:0]ID;
    input n43603;
    output n42551;
    output n27752;
    output [7:0]\data_out_frame[24] ;
    input n47614;
    output [7:0]\data_out_frame[25] ;
    input n42541;
    input n42790;
    output LED_c;
    output n49422;
    input n28189;
    output n43610;
    output n27554;
    input n28188;
    output n42897;
    output \data_out_frame[18][6] ;
    output n40598;
    input n28187;
    input n28186;
    output [23:0]neopxl_color;
    input n28185;
    output \Ki[0] ;
    input n28184;
    output \Kp[0] ;
    input n28183;
    input n28738;
    output [23:0]IntegralLimit;
    input n28737;
    input n28736;
    input n28735;
    input n28734;
    input n28733;
    input n28732;
    input n28731;
    input n28730;
    input n28729;
    input n28728;
    input n28727;
    input n28726;
    input n28725;
    input n28724;
    input n28723;
    input n28722;
    input n28721;
    input n28720;
    input n28719;
    input n28718;
    input n28717;
    input n28716;
    input n28715;
    input n28714;
    input n28713;
    input n28712;
    input n28711;
    input n28710;
    input n28709;
    input n28708;
    input n28707;
    input n28706;
    input n28705;
    input n28704;
    input n28703;
    input n28702;
    input n28701;
    input n28700;
    input n28698;
    input n28697;
    input n28696;
    input n28695;
    input n28694;
    input n28693;
    input n28692;
    input n28691;
    input n28690;
    input n28689;
    input n28688;
    input n28687;
    input n28686;
    input n28685;
    input n28684;
    input n28683;
    output \Kp[1] ;
    input n28682;
    output \Kp[2] ;
    input n28681;
    output \Kp[3] ;
    input n28680;
    output \Kp[4] ;
    input n28679;
    output \Kp[5] ;
    input n28678;
    output \Kp[6] ;
    input n28677;
    output \Kp[7] ;
    input n28676;
    output \Kp[8] ;
    input n28675;
    output \Kp[9] ;
    input n28674;
    output \Kp[10] ;
    input n28673;
    output \Kp[11] ;
    input n28672;
    output \Kp[12] ;
    input n28671;
    output \Kp[13] ;
    input n28670;
    output \Kp[14] ;
    input n28669;
    output \Kp[15] ;
    input n28668;
    output \Ki[1] ;
    input n28667;
    output \Ki[2] ;
    input n28666;
    output \Ki[3] ;
    input n28665;
    output \Ki[4] ;
    input n28664;
    output \Ki[5] ;
    input n28663;
    output \Ki[6] ;
    input n28662;
    output \Ki[7] ;
    input n28661;
    output \Ki[8] ;
    input n28660;
    output \Ki[9] ;
    input n28659;
    output \Ki[10] ;
    input n28658;
    output \Ki[11] ;
    input n28657;
    output \Ki[12] ;
    input n28656;
    output \Ki[13] ;
    input n28655;
    output \Ki[14] ;
    input n28654;
    output \Ki[15] ;
    input n28653;
    input n28652;
    input n28651;
    input n28650;
    input n28649;
    input n28648;
    input n28647;
    input n28646;
    input n28645;
    input n28644;
    input n28643;
    input n28642;
    input n28641;
    input n28640;
    input n28639;
    input n28638;
    input n28637;
    input n28636;
    input n28635;
    input n28634;
    input n28633;
    input n28632;
    input n28631;
    input n28630;
    input n28629;
    input n28628;
    input n28627;
    input n28626;
    input n28625;
    input n28624;
    input n28623;
    input n28622;
    input n28621;
    input n28620;
    input n28619;
    input n28618;
    input n28617;
    input n28616;
    input n28615;
    input n28614;
    input n28613;
    input n28612;
    input n28611;
    input n28610;
    input n28609;
    input n28608;
    input n28607;
    input n28606;
    input n28605;
    input n28604;
    input n28603;
    input n28602;
    input n28601;
    input n28600;
    input n28599;
    input n28598;
    input n28597;
    input n28596;
    input n28595;
    input n28594;
    input n28593;
    input n28592;
    input n28591;
    input n28590;
    input n28589;
    input n28588;
    input n28587;
    input n28586;
    input n28585;
    input n28584;
    input n28583;
    input n28582;
    output [7:0]rx_data;
    input n28581;
    input n28580;
    input n28579;
    input n28578;
    input n28577;
    input n28576;
    input n28575;
    input n28574;
    input n28573;
    input n28572;
    input n28571;
    input n28570;
    input n28569;
    input n28568;
    input n28567;
    input n28566;
    input n28565;
    input n28564;
    input n28563;
    input n28562;
    input n28561;
    input n28560;
    input n28559;
    input n28558;
    input n28557;
    input n28556;
    input n28555;
    input n28554;
    input n28553;
    input n28552;
    input n28551;
    input n28550;
    input n28549;
    input n28548;
    input n28547;
    input n28546;
    input n28545;
    input n28544;
    input n28543;
    input n28542;
    input n28541;
    input n28539;
    input n28538;
    input n28537;
    input n28536;
    input n28535;
    input n28534;
    input n28533;
    input n28532;
    input n28531;
    input n28530;
    input n28529;
    input n28528;
    input n28527;
    input n28526;
    input n28525;
    input n28524;
    input n28523;
    input n28522;
    input n28521;
    input n28520;
    input n28519;
    input n28518;
    input n28517;
    input n28516;
    input n28515;
    input n28514;
    input n28513;
    input n28512;
    input n28511;
    input n28510;
    input n28509;
    input n28508;
    input n28507;
    input n28164;
    input n28506;
    input n28505;
    input n28504;
    input n28503;
    input n28502;
    input n28501;
    input n28500;
    input n28499;
    input n28498;
    input n28497;
    input n28496;
    input n28495;
    input n28494;
    input n28493;
    input n28492;
    input n28491;
    input n28490;
    input n28489;
    input n28488;
    input n28487;
    input n28486;
    input n28485;
    input n28484;
    input n28483;
    input n28482;
    input n28481;
    input n28480;
    input n28479;
    input n28478;
    input n28477;
    input n28476;
    input n28475;
    input n28474;
    input n28473;
    input n28472;
    input n28471;
    input n28470;
    input n28469;
    input n28468;
    input n28467;
    input n28466;
    input n28465;
    input n28464;
    input n28405;
    input n28403;
    input n28402;
    input n28401;
    input n28400;
    input n28399;
    input n28398;
    input n28397;
    output n4;
    input \state[0] ;
    input \state[2] ;
    input \state[3] ;
    output n6014;
    input \displacement[17] ;
    output n27753;
    output n42230;
    output n42229;
    output \r_SM_Main_2__N_3513[1] ;
    output [2:0]r_SM_Main;
    output \r_Bit_Index[0] ;
    output n42123;
    output n27820;
    output tx_o;
    output n19247;
    input n49552;
    input n28192;
    output n4_adj_6;
    input n28212;
    input VCC_net;
    output tx_enable;
    output n4_adj_7;
    output [2:0]r_SM_Main_adj_14;
    output r_Rx_Data;
    output \r_SM_Main_2__N_3442[2] ;
    output n27824;
    output \r_Bit_Index[0]_adj_11 ;
    output n26628;
    output n33696;
    input RX_N_10;
    output n42126;
    input n41813;
    input n28224;
    input n28182;
    input n28181;
    input n28180;
    output n27784;
    input n28179;
    input n28178;
    input n28177;
    input n28176;
    input n42185;
    input n28215;
    output n26633;
    output n4_adj_12;
    output n4_adj_13;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n28295;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n28294, n28293;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n8, n5785, n5787, n5788, n5789, n7, n37247;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n37248, n5790, n5791, n5792, n5793;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n5794, n5795, n2, n3, n5796, n5797, n5798, n5799, n5800, 
        n5801;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, 
        Kp_23__N_761, n2482, n26617, n84, n3_adj_4109, n3_adj_4110, 
        Kp_23__N_993, n42388, n27427, n3_adj_4111;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n8_adj_4112;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n6, n3_adj_4113, n42654;
    wire [7:0]n8825;
    
    wire n27768, n36013;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(102[12:33])
    
    wire n3_adj_4114, n3_adj_4115, n3_adj_4116, n3_adj_4117, n3_adj_4118, 
        n18, n2_adj_4119, n37246, n3_adj_4120, n42416, n27200, n42422, 
        n42443, n27066, n6_adj_4121, n42353, n42548;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n42747, n40241, n42483, Kp_23__N_830, n42883, n6_adj_4122, 
        n42738, n42566, n26819, n42246, n6_adj_4123, Kp_23__N_869, 
        n27534, n42255, n12, n26903, n42360, n42721, n6_adj_4124, 
        Kp_23__N_996, n16, n27360, n42724, n42391, n22, n24, n42295, 
        n20, n27660, n40132, n42404, Kp_23__N_1095, n42265, n23, 
        n42410, n12_adj_4125, n42413, Kp_23__N_836, n44642, n3_adj_4126, 
        n27381, n27417, n10, n26999, n26, n26969, n40128, n8_adj_4127, 
        n27, n27061, n25, n28, n31, n24130, n31_adj_4128, n1, 
        n5786, n3_adj_4129, n161, n44461, n10_adj_4130;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n6_adj_4131, n3_adj_4132, n3_adj_4133;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n26861, n42538, n3_adj_4134, n3_adj_4135, n46778;
    wire [2:0]r_SM_Main_2__N_3516;
    
    wire n43085, n3_adj_4136, n3_adj_4137, n3_adj_4138, n3_adj_4139, 
        \FRAME_MATCHER.rx_data_ready_prev , n41663, n41655, n42249, 
        n10_adj_4140, n27762, n40257, n3_adj_4141, n3_adj_4142, n42797, 
        Kp_23__N_1210, n24_adj_4143, n8_adj_4144, n26688, n4452, n42918, 
        n42252, n36017, n49, n33593, n3183, n14, n26691, n15, 
        n26519, n10_adj_4145, n10_adj_4146, n14_adj_4147, n26694, 
        n16_adj_4148, n17, n26625, n16_adj_4149, n17_adj_4150, n63, 
        n42289, n18_adj_4151, n20_adj_4152, n15_adj_4153, n63_adj_4154, 
        n10_adj_4155, n42677, n27594, n40606, n42900, n14_adj_4156, 
        n10_adj_4157, n40578, n20_adj_4158, n19, n46542, n63_adj_4159, 
        n23831;
    wire [31:0]\FRAME_MATCHER.state_31__N_2560 ;
    
    wire n5, n771, n44, n42, n43, n41, n40, n39, n50, n45, 
        n26494, n8_adj_4160, n3303, n52, n42940, n42938, n4_c, 
        n81, n33940, n6_adj_4161, n26646, n26622, n34511, n359, 
        n59, n46777, n46776, n42837, n42619, n10_adj_4162, n46641, 
        n46642, n46633, n46632, n42591, n42753, n42471, n42741, 
        n42357, n42269, n27414, n40544, n42665, n47620, n38;
    wire [31:0]\FRAME_MATCHER.state_31__N_2624 ;
    
    wire n43623, n43490, n6_adj_4163, n27469, n42894, n12_adj_4164, 
        Kp_23__N_1206, n10_adj_4165, n42434, n42813, n42437, n42687, 
        n42258, n42298, n10_adj_4166, n42690, n26858, Kp_23__N_1402, 
        n16_adj_4167, n17_adj_4168, n47594, n47593, n42323, n42400, 
        n22_adj_4169, n42335, n42367, n26_adj_4170, n42880, n42385, 
        Kp_23__N_1466, n41649, n41721, n6_adj_4171, n43097, n44935, 
        n26924, Kp_23__N_990, Kp_23__N_1182, n42705, n27054, n42850, 
        n42662, n13, n11, n1475, n78, n10_adj_4172, n5_adj_4173, 
        n26482, n39630, n42657, n42633, n26870, n46730, n46728, 
        n49308, n49302, n14_adj_4174, n49266, n47592, n46721, n46719, 
        n49278, n49272, n14_adj_4175, n10_adj_4176, n25058, n26838, 
        n48074, n49529, n49530, n26942, n26981, n40506, n10_adj_4177, 
        n6_adj_4178, n42744, n42594, n42426, n26_adj_4179, n42449, 
        n24_adj_4180, n27639, n25_adj_4181, n23_adj_4182, n39681, 
        n10_adj_4183, n27347, n39699, n42844, n14_adj_4184, n10_adj_4185, 
        n44467, n7_adj_4186, n42906, n42636, n46714, n27041, n26223, 
        n46715, n46713, n42500, n12_adj_4187, n87, n10_adj_4188, 
        n11_adj_4189, n9, n49338, n49332, n14_adj_4190, n49428, 
        n47595, n46675, n49398, n48080, n46708, n10_adj_4191, Kp_23__N_1233, 
        n27438, n42506, n6_adj_4192, n40198, n42480, n10_adj_4193, 
        n44382, n12_adj_4194, n8_adj_4195, n6_adj_4196, n42786, n18_adj_4197, 
        n20_adj_4198, n42756, n16_adj_4199, n42584, n44495, n42580, 
        n40652, n42865, n10_adj_4200, n40524, n40570, n42825;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n4_adj_4201, n46709, n46707, n8_adj_4202, n42613, n43997, 
        n43562, n42525, n40504, n44626, n43581, n49326, n49416, 
        n14_adj_4203, n42491, n44122, n39733, n44455, n6_adj_4204, 
        n49434, n47601, n40629, n50_adj_4205, n46672, n43998, n44475, 
        n49392, n48086, n46702, n46703, n46701, n41717, n41769, 
        n49320, n49458, n14_adj_4206, n49440, n47604, n46669, n7_adj_4207, 
        n8_adj_4208, n41715, n41771, n41713, n41773, n41711, n41775, 
        n41709, n41729, n41707, n41725, n41705, n41777, n7_adj_4209, 
        n41779, n41703, n41781, n41701, n41783, n43666, n49386, 
        n48092, n46696, n41699, n41785, n41697, n41787, n41695, 
        n41789, n41693, n41791, n41691, n41793, n41689, n41743, 
        n41687, n41795, n41685, n41797, n41683, n41799, n41681, 
        n41741, n41679, n41801, n41677, n41803, n7_adj_4210, n41739, 
        n41675, n41737, n41673, n41805, n41671, n41669, n41665, 
        n41733, n46697, n46695, n40235, n44775, n44445, n7_adj_4211, 
        n40502, n43715, n18_adj_4212, n46540, n44001, n42768, n46427, 
        n43504, n23_adj_4213, n27_adj_4214, n29, n42915, n42732, 
        n48, n49314, n49482, n14_adj_4215, n49446, n47607, n46666, 
        n49380, n48096, n49_adj_4216, n46688, n46686, n49452, n47611, 
        n46663, n49374, n48100, n46684, n46685, n46683, n49290, 
        n49284, n14_adj_4217, n49464, n47617, n46657, n49362, n48104, 
        n44563, n27893;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n42407, n47, n43_adj_4218, n42611, n43933, n42625, n44321, 
        n43986, n42627, n42905, n44856;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n43837, n43664, n43918, n44471, n43527, n43931, n42604, 
        n40634, n42649, n14_adj_4219, n10_adj_4220, n42497, n27210, 
        n39632, n46, n48_adj_4221, n46_adj_4222, n47_adj_4223, n45_adj_4224, 
        n54, n49515, n7_adj_4225;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n49_adj_4226, n49509, n26951, n42458, n45_adj_4227, n44027, 
        n42616, n49404, n7_adj_4228, n44_adj_4229, n49503, n7_adj_4230, 
        n49497, n7_adj_4231, n49491, n7_adj_4232, n49485, n7_adj_4233, 
        n49479, n49473, n7_adj_4234, n49260, n49467, n7_adj_4235, 
        n49461, n49455, n49449, n42607, n27239, n14_adj_4236, n2_adj_4237, 
        n2_adj_4238, n2_adj_4239, n2_adj_4240, n2_adj_4241, n2_adj_4242, 
        n2_adj_4243, n2_adj_4244, n2_adj_4245, n2_adj_4246, n2_adj_4247, 
        n2_adj_4248, n2_adj_4249, n2_adj_4250, n2_adj_4251, n2_adj_4252, 
        n2_adj_4253, n2_adj_4254, n2_adj_4255, n2_adj_4256, n2_adj_4257, 
        n2_adj_4258, n2_adj_4259, n3_adj_4260, n2_adj_4261, n3_adj_4262, 
        n2_adj_4263, n3_adj_4264, n2_adj_4265, n3_adj_4266, n2_adj_4267, 
        n3_adj_4268, n2_adj_4269, n3_adj_4270, n2_adj_4271, n3_adj_4272, 
        n2_adj_4273, n3_adj_4274, n3_adj_4275, n10_adj_4276, n40554, 
        n56, \FRAME_MATCHER.i_31__N_2524 , n85, n49443, n49437, n49431, 
        n30, n51, n42535, n39689, n42903, n16_adj_4277, n27196, 
        n19_adj_4278, n44066, n49425, n22_adj_4279, n40073, n42834, 
        n43940, n40668, n40114, n42645, n42646, n17_adj_4280, n40586, 
        n42801, n40283, n42780, n6_adj_4281, n26238, n42648, n27181, 
        n42550, n12_adj_4282, n27679, n42759, n50_adj_4283, n40658, 
        n42774, n48_adj_4284, n42886, n26258, n49_adj_4285, n42312, 
        n42503, n47_adj_4286, n39650, n42771, n30_adj_4287, n42588, 
        n46_adj_4288, n42486, n45_adj_4289, n56_adj_4290, n42522, 
        n51_adj_4291, n27998, n43465, n42519, n40517, n6_adj_4292, 
        n33507, n42206, n49419, n49413, n49401, n49395, n49389, 
        n49383, n49377, n2206, n44460, n27517, n39761, n26774, 
        n6_adj_4293, n40052, n40673, n42513, n42840, n42699, n42601, 
        n26235, n42378, n42735, n40033, n27223, n27569, n23_adj_4294;
    wire [7:0]\data_out_frame[18]_c ;   // verilog/coms.v(97[12:26])
    
    wire n49371, n1794, n27321, n22_adj_4295, n20_adj_4296, n40582, 
        n26_adj_4297, n49359, n49335, n49329, n49323, n40512, n40576, 
        n42783, n42553, n42241, n39724, n24914, n27337, n27340, 
        n12_adj_4298, n37283, n37282, n37281, n2063, n39642, n37280, 
        n42777, n6_adj_4299, n27113, n48504, n48508, n37279, n6_adj_4300, 
        n42274, n6_adj_4301, n42462, n37278, n6_adj_4302, n43813, 
        n37277, n42639, n6_adj_4303, n42804, n42831, tx_transmit_N_3413, 
        n10_adj_4304, n16_adj_4305, n42816, n12_adj_4306, n37276, 
        n42559, n1673, n42762, n10_adj_4307, n1516, n1513, n37275, 
        n42610, n37274, n1_adj_4308, n1_adj_4309, n37273, n37272, 
        n42455, n42765, n18_adj_4310, n42909, n20_adj_4311, n42847, 
        n16_adj_4312, n42598, n42494, n42286, n6_adj_4313, n27128, 
        n42465, n37271, n42877, n37270, n37269, n42674, n27705, 
        n14_adj_4314, n10_adj_4315, n27215, n42277, n16_adj_4316, 
        n42668, n17_adj_4317, n27547, n42874, n26939, n14_adj_4318, 
        n10_adj_4319, n27492, n42718, n12_adj_4320, n27627, n42793, 
        n42622, n27121, n42338, n6_adj_4321, n37268, n49317, n49311, 
        n42856, n42912, n40604, n42853, n10_adj_4322, n42452, n1519, 
        n9_adj_4323, n49305, n27666, n42331, n6_adj_4324, n1668, 
        n42364, n42711, n10_adj_4325, n27498, n12_adj_4326, n1522, 
        n42238, n42708, n10_adj_4327, n36, n34, n42431, n42243, 
        n39_adj_4328, n42468, n38_adj_4329, n42510, n42302, n37, 
        n49299, n27278, n40530, n41_adj_4330, n26822, n43_adj_4331, 
        n44221, n36_adj_4332, n42822, n42642, n34_adj_4333, n26_adj_4334, 
        n40_adj_4335, n38_adj_4336, n42_adj_4337, n37_adj_4338, n42576, 
        n42819, n12_adj_4339, n42807, n42868, n42394, n42696, n27406, 
        n26702, n1191, n42262, n6_adj_4340, n42488, n42544, n2_adj_4341, 
        n4_adj_4342, n7_adj_4343, n2_adj_4344, n5_adj_4345, n37267, 
        n37266, n40542, n36_adj_4346, n37265, n34_adj_4347, n37264, 
        n37263;
    wire [31:0]n92;
    
    wire n27_adj_4348, n37262, n39_adj_4349, n42862, n38_adj_4350, 
        n42563, n37_adj_4351, n42572, n41_adj_4352, n42810, n42397, 
        n43_adj_4353, n42750, n10_adj_4354, n40112, n42680, n10_adj_4355, 
        n42859, n42651, n14_adj_4356, n42235, n27324, n40347, n42528, 
        n42292, n6_adj_4357, n27026, n27461, n42344, n6_adj_4358, 
        n42891, n42556, n42727, n6_adj_4359, n14_adj_4360, n26217, 
        n1510, n27103, n42671, n26725, n6_adj_4361, n26771, n27287, 
        n6_adj_4362, n8_adj_4363, n42216, n6_adj_4364, n26762, n10_adj_4365, 
        n14_adj_4366, n42673, n42871, n10_adj_4367, n2122, n6_adj_4368, 
        n40662, n10_adj_4369, n42231, n10_adj_4370, n42225, n28456, 
        n28457, n37261, n29941, n7_adj_4371, n28458, n28459, n28460, 
        n8_adj_4372, n42219, n37260, n28461, n28462, n28463, n42222, 
        n28448, n28449, n28450, n28451, n28452, n28453, n37259, 
        n28454, n28455, n37258, n8_adj_4373, n8_adj_4374, n37257, 
        n42693, n42213, n37256, n28440, n37255, \FRAME_MATCHER.i_31__N_2523 , 
        n28441, n28442, n28443, n28540, n28296, n28444, n28445, 
        n28446, n28447, n28432, n28433, n28434, n28435, n28436, 
        n28437, n28438, n28439, n28431, n28430, n28429, n28428, 
        n28427, n28426, n28425, n28424, n28423, n28422, n28421, 
        n28420, n28419, n28418, n28417, n28416, n28415, n28414, 
        n28413, n28410, n28409, n28408, n28407, n28406, n28396, 
        n28395, n28394, n28393, n28392, n28391, n28390, n28389, 
        n28388, n28387, n28386, n28385, n28384, n28383, n28382, 
        n28381, n28380, n28379, n28378, n28377, n28376, n28375, 
        n28374, n28373, n28372, n28371, n28370, n28369, n28368, 
        n28367, n28366, n28365, n28364, n28363, n28362, n28361, 
        n28360, n28359, n28358, n28357, n28356, n28355, n28354, 
        n28353, n28352, n28351, n28350, n28349, n28348, n28347, 
        n28346, n28345, n28344, n28343, n28342, n28341, n28340, 
        n28339, n28338, n28337, n28336, n28335, n28334, n28333, 
        n28332, n28331, n28330, n28329, n28328, n28327, n28326, 
        n28325, n28324, n28323, n28322, Kp_23__N_1221, n28321, n28320, 
        n28319, n28318, n28317, n28316, n28315, n28314, n28313, 
        n28312, n28311, n28310, n28309, n28308, n28307, n28306, 
        n28305, n43987, n37254, n26_adj_4375, n30_adj_4376, n23_adj_4377, 
        n46425, n32, n5_adj_4378, n28304, n27_adj_4379, n28303, 
        n28302, n22_adj_4380, n8_adj_4381, n37253, n28301, n28300, 
        n28299, n12_adj_4382, n28298, n28297, n42203, n37252, n37251, 
        n37250, n37249, n49287, n43891, n8_adj_4384, n39_adj_4385, 
        n1_adj_4386, n10_adj_4387, n5_adj_4388, n6_adj_4389;
    wire [31:0]\FRAME_MATCHER.state_31__N_2720 ;
    
    wire n5_adj_4390, n10_adj_4391, n49281, n49275, n49269, n49263, 
        n49257;
    
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n28295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n28294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n28293));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n28292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n28291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n28290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n28289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n28288));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n8));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1362_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n5785), .I3(GND_net), .O(n5787));
    defparam mux_1362_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n5785), .I3(GND_net), .O(n5788));
    defparam mux_1362_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n5785), .I3(GND_net), .O(n5789));
    defparam mux_1362_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n28287));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_43_4 (.CI(n37247), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n37248));
    SB_LUT4 mux_1362_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n5785), .I3(GND_net), .O(n5790));
    defparam mux_1362_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n5785), .I3(GND_net), .O(n5791));
    defparam mux_1362_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n5785), .I3(GND_net), .O(n5792));
    defparam mux_1362_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n5785), .I3(GND_net), .O(n5793));
    defparam mux_1362_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n5785), .I3(GND_net), .O(n5794));
    defparam mux_1362_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n5785), .I3(GND_net), .O(n5795));
    defparam mux_1362_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1362_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n5785), .I3(GND_net), .O(n5796));
    defparam mux_1362_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n5785), .I3(GND_net), .O(n5797));
    defparam mux_1362_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n5785), .I3(GND_net), .O(n5798));
    defparam mux_1362_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n28286));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1362_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n5785), .I3(GND_net), .O(n5799));
    defparam mux_1362_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n5785), .I3(GND_net), .O(n5800));
    defparam mux_1362_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n5785), .I3(GND_net), .O(n5801));
    defparam mux_1362_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n5785), .I3(GND_net), .O(n5802));
    defparam mux_1362_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n5785), .I3(GND_net), .O(n5803));
    defparam mux_1362_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n5785), .I3(GND_net), .O(n5804));
    defparam mux_1362_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n28285));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n28284));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1362_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n5785), .I3(GND_net), .O(n5805));
    defparam mux_1362_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n5785), .I3(GND_net), .O(n5806));
    defparam mux_1362_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n5785), .I3(GND_net), .O(n5807));
    defparam mux_1362_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n5785), .I3(GND_net), .O(n5808));
    defparam mux_1362_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1362_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n5785), .I3(GND_net), .O(n5809));
    defparam mux_1362_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[19] [1]), .I1(n7), .I2(\data_in_frame[19] [7]), 
            .I3(n8), .O(Kp_23__N_761));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_428_Select_10_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4109));
    defparam select_428_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_11_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4110));
    defparam select_428_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[8] [5]), .I1(Kp_23__N_993), .I2(\data_in_frame[6] [3]), 
            .I3(n42388), .O(n27427));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_428_Select_12_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4111));
    defparam select_428_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i4_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n8_adj_4112), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n23943));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut.LUT_INIT = 16'h0440;
    SB_LUT4 i1_2_lut_adj_851 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_851.LUT_INIT = 16'h6666;
    SB_LUT4 select_428_Select_13_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4113));
    defparam select_428_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i4_4_lut_adj_852 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[10] [6]), .I3(n6), .O(n42654));
    defparam i4_4_lut_adj_852.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n27768), .D(n8825[1]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
            .E(n27768), .D(n8825[2]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), 
            .C(CLK_c), .E(n27768), .D(n8825[3]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), 
            .C(CLK_c), .E(n27768), .D(n8825[4]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(CLK_c), .E(n27768), .D(n8825[5]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(CLK_c), .E(n27768), .D(n8825[6]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(CLK_c), .E(n27768), .D(n8825[7]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n28283));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_428_Select_14_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4114));
    defparam select_428_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_15_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4115));
    defparam select_428_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_16_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4116));
    defparam select_428_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n28282));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_428_Select_17_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4117));
    defparam select_428_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_18_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4118));
    defparam select_428_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i4_2_lut (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n18));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n28281));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_3_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n37246), .O(n2_adj_4119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n28280));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_428_Select_19_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4120));
    defparam select_428_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_CARRY add_43_3 (.CI(n37246), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n37247));
    SB_LUT4 i1_2_lut_adj_853 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42416));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_853.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_854 (.I0(\data_in_frame[5] [3]), .I1(n27200), .I2(GND_net), 
            .I3(GND_net), .O(n42422));
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(n42443), .I1(n27066), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_4121));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[5] [6]), 
            .I2(n6_adj_4121), .I3(n42353), .O(n42548));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_855 (.I0(\data_in_frame[7] [5]), .I1(n42747), .I2(n42422), 
            .I3(\data_in_frame[5] [4]), .O(n40241));
    defparam i3_4_lut_adj_855.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_856 (.I0(\data_in_frame[6] [7]), .I1(n42483), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_830));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_856.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_857 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42883));
    defparam i1_2_lut_adj_857.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_858 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[1] [4]), .I3(GND_net), .O(n42353));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_858.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_859 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4122));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_859.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_860 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[3] [6]), .I3(n6_adj_4122), .O(n42738));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_860.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_861 (.I0(\data_in_frame[5] [5]), .I1(n42566), .I2(GND_net), 
            .I3(GND_net), .O(n26819));
    defparam i1_2_lut_adj_861.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_862 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(n42246), .I3(n6_adj_4123), .O(Kp_23__N_869));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_863 (.I0(n27534), .I1(\data_in_frame[5] [1]), .I2(n42255), 
            .I3(\data_in_frame[2] [7]), .O(n12));   // verilog/coms.v(77[16:27])
    defparam i5_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(n26903), .I1(n12), .I2(\data_in_frame[4] [6]), 
            .I3(n42360), .O(n42721));   // verilog/coms.v(77[16:27])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_864 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[4] [2]), .I3(n6_adj_4124), .O(Kp_23__N_996));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_864.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut (.I0(n42721), .I1(Kp_23__N_869), .I2(GND_net), .I3(GND_net), 
            .O(n16));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut (.I0(n27360), .I1(n42724), .I2(n42747), .I3(n42391), 
            .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(n42353), .I1(n22), .I2(n16), .I3(n42883), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n42295), .I1(n24), .I2(n20), .I3(n27660), 
            .O(n40132));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_865 (.I0(n40132), .I1(Kp_23__N_830), .I2(n42404), 
            .I3(\data_in_frame[6] [0]), .O(n42443));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_865.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n28279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n28278));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut (.I0(Kp_23__N_1095), .I1(n42265), .I2(\data_in_frame[8] [6]), 
            .I3(n42443), .O(n23));
    defparam i7_4_lut.LUT_INIT = 16'hde7b;
    SB_LUT4 i5_4_lut_adj_866 (.I0(\data_in_frame[8] [1]), .I1(n42410), .I2(n40132), 
            .I3(Kp_23__N_996), .O(n12_adj_4125));
    defparam i5_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_867 (.I0(Kp_23__N_830), .I1(n12_adj_4125), .I2(n42413), 
            .I3(Kp_23__N_836), .O(n44642));
    defparam i6_4_lut_adj_867.LUT_INIT = 16'h6996;
    SB_LUT4 select_428_Select_20_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4126));
    defparam select_428_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i10_4_lut (.I0(n27381), .I1(n27417), .I2(n10), .I3(n26999), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_868 (.I0(n26969), .I1(n44642), .I2(n40128), 
            .I3(n8_adj_4127), .O(n27));
    defparam i11_4_lut_adj_868.LUT_INIT = 16'hffef;
    SB_LUT4 i9_4_lut_adj_869 (.I0(n40241), .I1(n42548), .I2(n27061), .I3(n27427), 
            .O(n25));
    defparam i9_4_lut_adj_869.LUT_INIT = 16'hfffb;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n31));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20513_4_lut (.I0(n24130), .I1(n31_adj_4128), .I2(n31), .I3(\FRAME_MATCHER.state [1]), 
            .O(n1));
    defparam i20513_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 mux_1362_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n5785), .I3(GND_net), .O(n5786));
    defparam mux_1362_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n28277));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_428_Select_21_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4129));
    defparam select_428_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 add_43_2_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_870 (.I0(\data_in_frame[10] [1]), .I1(n26999), 
            .I2(n44461), .I3(n27381), .O(n10_adj_4130));
    defparam i4_4_lut_adj_870.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_871 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[12] [6]), 
            .I2(n10_adj_4130), .I3(\data_in_frame[17] [1]), .O(n6_adj_4131));
    defparam i1_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n37246));
    SB_LUT4 select_428_Select_22_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4132));
    defparam select_428_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_23_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4133));
    defparam select_428_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i4_4_lut_adj_872 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[14] [5]), 
            .I2(n26861), .I3(n6_adj_4131), .O(n42538));
    defparam i4_4_lut_adj_872.LUT_INIT = 16'h6996;
    SB_LUT4 select_428_Select_24_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4134));
    defparam select_428_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_25_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4135));
    defparam select_428_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n28276));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3516[0]), .C(CLK_c), .D(n46778), 
            .R(n43085));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_428_Select_26_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4136));
    defparam select_428_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_27_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4137));
    defparam select_428_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_28_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4138));
    defparam select_428_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_29_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4139));
    defparam select_428_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(CLK_c), 
            .D(n41663), .S(n41655));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_873 (.I0(n42249), .I1(n27381), .I2(\data_in_frame[17] [2]), 
            .I3(n42654), .O(n10_adj_4140));
    defparam i4_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n27762), .D(n5786));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[12] [7]), .I1(n10_adj_4140), .I2(n27427), 
            .I3(GND_net), .O(n40257));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_428_Select_30_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4141));
    defparam select_428_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_31_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4142));
    defparam select_428_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i10_4_lut_adj_874 (.I0(n42797), .I1(\data_in_frame[1] [6]), 
            .I2(Kp_23__N_1210), .I3(\data_in_frame[8] [3]), .O(n24_adj_4143));
    defparam i10_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_LUT4 select_428_Select_0_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_428_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i20785_4_lut (.I0(n8_adj_4144), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n26688), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i20785_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_875 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42918));
    defparam i1_2_lut_adj_875.LUT_INIT = 16'h6666;
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n28275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n28274));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[1] [1]), .I1(n42252), .I2(\data_in_frame[3] [2]), 
            .I3(\data_in_frame[5] [4]), .O(n42566));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_876 (.I0(n36017), .I1(n49), .I2(n33593), .I3(n2482), 
            .O(n3183));
    defparam i3_4_lut_adj_876.LUT_INIT = 16'h0020;
    SB_LUT4 i5_3_lut_adj_877 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14));
    defparam i5_3_lut_adj_877.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_878 (.I0(\data_in[0] [6]), .I1(n26691), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15));
    defparam i6_4_lut_adj_878.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(\data_in[2] [2]), .I2(n14), .I3(\data_in[0] [3]), 
            .O(n26519));
    defparam i8_4_lut.LUT_INIT = 16'hfbff;
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n28273));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_879 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4145));
    defparam i4_4_lut_adj_879.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_880 (.I0(\data_in[3] [4]), .I1(n10_adj_4145), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n26691));
    defparam i5_3_lut_adj_880.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut_adj_881 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4146));
    defparam i2_2_lut_adj_881.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_882 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4147));
    defparam i6_4_lut_adj_882.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_883 (.I0(\data_in[3] [6]), .I1(n14_adj_4147), .I2(n10_adj_4146), 
            .I3(\data_in[2] [1]), .O(n26694));
    defparam i7_4_lut_adj_883.LUT_INIT = 16'hfffd;
    SB_LUT4 i6_4_lut_adj_884 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4148));
    defparam i6_4_lut_adj_884.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_885 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut_adj_885.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_886 (.I0(n17), .I1(\data_in[1] [6]), .I2(n16_adj_4148), 
            .I3(\data_in[3] [7]), .O(n26625));
    defparam i9_4_lut_adj_886.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_887 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n26519), .O(n16_adj_4149));
    defparam i6_4_lut_adj_887.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_888 (.I0(n26625), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4150));
    defparam i7_4_lut_adj_888.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_889 (.I0(n17_adj_4150), .I1(\data_in[3] [5]), .I2(n16_adj_4149), 
            .I3(\data_in[3] [3]), .O(n63));
    defparam i9_4_lut_adj_889.LUT_INIT = 16'hfbff;
    SB_LUT4 i3_4_lut_adj_890 (.I0(\data_in_frame[12] [6]), .I1(n42918), 
            .I2(\data_in_frame[8] [6]), .I3(Kp_23__N_1095), .O(n42289));
    defparam i3_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_891 (.I0(\data_in[2] [4]), .I1(n26694), .I2(\data_in[1] [5]), 
            .I3(n26691), .O(n18_adj_4151));
    defparam i7_4_lut_adj_891.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_892 (.I0(\data_in[0] [6]), .I1(n18_adj_4151), .I2(\data_in[3] [0]), 
            .I3(n26625), .O(n20_adj_4152));
    defparam i9_4_lut_adj_892.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_893 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4153));
    defparam i4_2_lut_adj_893.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_894 (.I0(n15_adj_4153), .I1(n20_adj_4152), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_4154));
    defparam i10_4_lut_adj_894.LUT_INIT = 16'hfeff;
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n28272));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[17] [3]), .I3(GND_net), .O(n10_adj_4155));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_895 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42677));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_896 (.I0(n40128), .I1(\data_in_frame[9] [0]), .I2(n27594), 
            .I3(n40606), .O(n42900));
    defparam i3_4_lut_adj_896.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_897 (.I0(n42900), .I1(n27061), .I2(n42677), .I3(\data_in_frame[13] [0]), 
            .O(n14_adj_4156));
    defparam i6_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_898 (.I0(\data_in_frame[17] [4]), .I1(n14_adj_4156), 
            .I2(n10_adj_4157), .I3(n42289), .O(n40578));
    defparam i7_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_899 (.I0(n26694), .I1(\data_in[1] [3]), .I2(n26519), 
            .I3(\data_in[2] [0]), .O(n20_adj_4158));
    defparam i8_4_lut_adj_899.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_900 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19));
    defparam i7_4_lut_adj_900.LUT_INIT = 16'hfeff;
    SB_LUT4 i31663_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [5]), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [2]), .O(n46542));
    defparam i31663_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n46542), .I1(n19), .I2(n20_adj_4158), .I3(GND_net), 
            .O(n63_adj_4159));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\FRAME_MATCHER.state [0]), .I1(n23831), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2560 [0]));
    defparam i1_2_lut_adj_901.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20778_4_lut (.I0(n5), .I1(\FRAME_MATCHER.i [31]), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i20778_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_902 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut_adj_902.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n26688));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_903 (.I0(\FRAME_MATCHER.i [4]), .I1(n26688), .I2(GND_net), 
            .I3(GND_net), .O(n26494));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_903.LUT_INIT = 16'heeee;
    SB_LUT4 i20784_4_lut (.I0(n8_adj_4160), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n26494), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i20784_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i28068_2_lut (.I0(n52), .I1(n4452), .I2(GND_net), .I3(GND_net), 
            .O(n42940));
    defparam i28068_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_904 (.I0(n36013), .I1(n42938), .I2(\FRAME_MATCHER.state_31__N_2560 [0]), 
            .I3(n4_c), .O(n41655));
    defparam i1_4_lut_adj_904.LUT_INIT = 16'hfaba;
    SB_LUT4 i2_3_lut_adj_905 (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[6]), 
            .I2(byte_transmit_counter_c[7]), .I3(GND_net), .O(n81));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_adj_905.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_906 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n33940));
    defparam i2_3_lut_adj_906.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_907 (.I0(n81), .I1(\FRAME_MATCHER.state [0]), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n6_adj_4161), .O(n26646));
    defparam i4_4_lut_adj_907.LUT_INIT = 16'hffbf;
    SB_LUT4 i21462_2_lut (.I0(n33940), .I1(n26622), .I2(GND_net), .I3(GND_net), 
            .O(n34511));
    defparam i21462_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut (.I0(\byte_transmit_counter[0] ), .I1(byte_transmit_counter[2]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n359));   // verilog/coms.v(102[12:33])
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i28210_4_lut (.I0(n26622), .I1(\FRAME_MATCHER.state [3]), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n84), .O(n43085));
    defparam i28210_4_lut.LUT_INIT = 16'heaee;
    SB_LUT4 i31824_3_lut (.I0(n59), .I1(n34511), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n46777));
    defparam i31824_3_lut.LUT_INIT = 16'h8b8b;
    SB_LUT4 i31823_3_lut (.I0(n26646), .I1(n34511), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n46776));
    defparam i31823_3_lut.LUT_INIT = 16'h8b8b;
    SB_LUT4 i31825_3_lut (.I0(n46776), .I1(n46777), .I2(n359), .I3(GND_net), 
            .O(n46778));
    defparam i31825_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_3_lut_adj_908 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[11] [1]), 
            .I2(n26999), .I3(GND_net), .O(n42837));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_908.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_909 (.I0(\data_in_frame[13] [1]), .I1(n42619), 
            .I2(\data_in_frame[15] [3]), .I3(n42837), .O(n10_adj_4162));
    defparam i4_4_lut_adj_909.LUT_INIT = 16'h6996;
    SB_LUT4 i31688_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46641));
    defparam i31688_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n28271));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31689_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46642));
    defparam i31689_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n28270));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n28269));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31680_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46633));
    defparam i31680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31679_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46632));
    defparam i31679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_910 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [7]), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n42591));
    defparam i2_3_lut_adj_910.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_911 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[11] [5]), 
            .I2(\data_in_frame[12] [0]), .I3(GND_net), .O(n42753));
    defparam i2_3_lut_adj_911.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_912 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[13] [6]), 
            .I2(n40606), .I3(n42471), .O(n42741));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_912.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42357));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_914 (.I0(n27381), .I1(n42269), .I2(n27414), .I3(n40544), 
            .O(n42665));
    defparam i3_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_915 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42471));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_916 (.I0(n43085), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n47620), .I3(n34511), .O(n38));
    defparam i1_4_lut_adj_916.LUT_INIT = 16'h5011;
    SB_LUT4 i3_4_lut_adj_917 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state_31__N_2624 [3]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n43623));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_917.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_3_lut_adj_918 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n1), .I3(GND_net), .O(n43490));
    defparam i2_3_lut_adj_918.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [6]), .I3(GND_net), .O(n6_adj_4123));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_919 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(n42548), .I3(n6_adj_4163), .O(n40544));
    defparam i4_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27469));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_921 (.I0(\data_in_frame[7] [6]), .I1(n40544), .I2(\data_in_frame[7] [7]), 
            .I3(GND_net), .O(n42894));
    defparam i2_3_lut_adj_921.LUT_INIT = 16'h6969;
    SB_LUT4 i33920_4_lut (.I0(n38), .I1(n34511), .I2(n43490), .I3(n43623), 
            .O(n12_adj_4164));
    defparam i33920_4_lut.LUT_INIT = 16'h2a22;
    SB_LUT4 i4_4_lut_adj_922 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[14] [4]), 
            .I2(\data_in_frame[12] [2]), .I3(Kp_23__N_1206), .O(n10_adj_4165));
    defparam i4_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_923 (.I0(n42434), .I1(n10_adj_4165), .I2(\data_in_frame[10] [0]), 
            .I3(GND_net), .O(n42813));
    defparam i5_3_lut_adj_923.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_924 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42437));
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h6666;
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n28268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n28267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n28266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n28265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n28264));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_925 (.I0(\data_in_frame[12] [1]), .I1(n40128), 
            .I2(GND_net), .I3(GND_net), .O(n42687));
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_926 (.I0(n42258), .I1(\data_in_frame[3] [5]), .I2(\data_in_frame[1] [4]), 
            .I3(n42298), .O(n10_adj_4166));
    defparam i4_4_lut_adj_926.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_927 (.I0(\data_in_frame[7] [7]), .I1(n10_adj_4166), 
            .I2(\data_in_frame[8] [0]), .I3(GND_net), .O(n42690));
    defparam i5_3_lut_adj_927.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_928 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26858));
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_16__7__I_0_3896_2_lut (.I0(\data_in_frame[16] [7]), 
            .I1(\data_in_frame[16] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1402));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_16__7__I_0_3896_2_lut.LUT_INIT = 16'h6666;
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n28263));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n16_adj_4167));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n17_adj_4168));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32840_2_lut (.I0(\data_out_frame[23] [7]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n47594));
    defparam i32840_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32842_2_lut (.I0(\data_out_frame[20] [7]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n47593));
    defparam i32842_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_929 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[5] [0]), .O(n42360));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut_adj_929.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_930 (.I0(\data_in_frame[6] [1]), .I1(Kp_23__N_836), 
            .I2(GND_net), .I3(GND_net), .O(n42323));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_930.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_931 (.I0(n42400), .I1(\data_in_frame[8] [4]), .I2(\data_in_frame[9] [7]), 
            .I3(\data_in_frame[9] [2]), .O(n22_adj_4169));
    defparam i8_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n27762), .D(n5809));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_932 (.I0(n26969), .I1(n10), .I2(\data_in_frame[9] [2]), 
            .I3(GND_net), .O(n42335));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_932.LUT_INIT = 16'h9696;
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n27762), .D(n5808));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n27762), .D(n5807));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n27762), .D(n5806));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n27762), .D(n5805));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n27762), .D(n5804));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n27762), .D(n5803));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n27762), .D(n5802));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n27762), .D(n5801));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n27762), .D(n5800));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_933 (.I0(n26969), .I1(n24_adj_4143), .I2(n18), 
            .I3(n42367), .O(n26_adj_4170));
    defparam i12_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n27762), .D(n5799));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n27762), .D(n5798));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n27762), .D(n5797));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n27762), .D(n5796));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n27762), .D(n5795));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[9] [0]), .I1(n26_adj_4170), .I2(n22_adj_4169), 
            .I3(\data_in_frame[8] [0]), .O(n42880));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n27762), .D(n5794));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n27762), .D(n5793));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n27762), .D(n5792));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n27762), .D(n5791));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n27762), .D(n5790));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n27762), .D(n5789));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n27762), .D(n5788));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n27762), .D(n5787));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_in_frame[11] [4]), .I1(n42385), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1466));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(CLK_c), 
            .D(n41649), .S(n41721));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n26969), .I1(n10), .I2(n27417), 
            .I3(n40128), .O(n40606));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(CLK_c), .E(n27768), .D(n8825[0]), .R(n36013));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_935 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(n27360), .I3(GND_net), .O(n6_adj_4124));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_935.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_936 (.I0(n27660), .I1(\data_in_frame[8] [2]), .I2(n27469), 
            .I3(n6_adj_4171), .O(n27061));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(CLK_c), .E(n43097), .D(n84), 
            .R(n44935));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_937 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26924));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_938 (.I0(\data_in_frame[8] [3]), .I1(n42323), .I2(Kp_23__N_990), 
            .I3(\data_in_frame[6] [2]), .O(n26999));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_939 (.I0(n26999), .I1(n27061), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1182));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_939.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_940 (.I0(n42335), .I1(n42705), .I2(\data_in_frame[11] [3]), 
            .I3(GND_net), .O(n27054));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_940.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_941 (.I0(n27427), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42850));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_942 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [4]), .I3(n42738), .O(Kp_23__N_990));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_943 (.I0(n27414), .I1(\data_in_frame[9] [1]), .I2(\data_in_frame[11] [2]), 
            .I3(\data_in_frame[13] [3]), .O(n42662));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_944 (.I0(n42894), .I1(n26819), .I2(\data_in_frame[12] [4]), 
            .I3(\data_in_frame[14] [6]), .O(n13));
    defparam i5_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_945 (.I0(n13), .I1(n11), .I2(\data_in_frame[12] [5]), 
            .I3(n27066), .O(n42249));
    defparam i7_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_946 (.I0(r_SM_Main_2__N_3516[0]), .I1(tx_active), 
            .I2(GND_net), .I3(GND_net), .O(n1475));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_946.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_947 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n78));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_947.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_948 (.I0(n42662), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[15] [5]), .I3(n42850), .O(n10_adj_4172));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i33915_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n5_adj_4173), 
            .I2(GND_net), .I3(GND_net), .O(n36013));
    defparam i33915_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n78), .I1(n36013), .I2(n26482), .I3(n1475), 
            .O(n27768));
    defparam i1_4_lut_adj_949.LUT_INIT = 16'hccce;
    SB_LUT4 i5_3_lut_adj_950 (.I0(n42269), .I1(n10_adj_4172), .I2(n27054), 
            .I3(GND_net), .O(n39630));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_950.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_951 (.I0(n42657), .I1(\data_in_frame[17] [0]), 
            .I2(n42249), .I3(GND_net), .O(n42633));
    defparam i2_3_lut_adj_951.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_952 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n26870));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_952.LUT_INIT = 16'h9696;
    SB_LUT4 i31777_4_lut (.I0(\data_out_frame[6] [7]), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n46730));
    defparam i31777_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i31775_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46728));
    defparam i31775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2171647_i1_3_lut (.I0(n49308), .I1(n49302), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4174));
    defparam i2171647_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32827_2_lut (.I0(n49266), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47592));
    defparam i32827_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31768_4_lut (.I0(\data_out_frame[6] [6]), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n46721));
    defparam i31768_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i31766_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46719));
    defparam i31766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_953 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n27066));
    defparam i1_2_lut_3_lut_adj_953.LUT_INIT = 16'h9696;
    SB_LUT4 i2172250_i1_3_lut (.I0(n49278), .I1(n49272), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4175));
    defparam i2172250_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[6] [1]), .I3(n10_adj_4176), .O(n25058));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_954 (.I0(n26838), .I1(n42721), .I2(\data_in_frame[7] [2]), 
            .I3(GND_net), .O(n27417));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_954.LUT_INIT = 16'h9696;
    SB_LUT4 i33121_3_lut (.I0(n49368), .I1(n46660), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48074));
    defparam i33121_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(CLK_c), 
           .D(n49529));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(CLK_c), 
           .D(n49530));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_955 (.I0(\data_in_frame[6] [1]), .I1(n26942), .I2(\data_in_frame[6] [4]), 
            .I3(n26981), .O(n42483));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_956 (.I0(Kp_23__N_1182), .I1(n40506), .I2(\data_in_frame[9] [0]), 
            .I3(n42665), .O(n10_adj_4177));
    defparam i4_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_957 (.I0(n27534), .I1(\data_in_frame[7] [4]), .I2(\data_in_frame[3] [2]), 
            .I3(n6_adj_4178), .O(n42744));
    defparam i4_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42594));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_959 (.I0(n42426), .I1(\data_in_frame[7] [1]), 
            .I2(\data_in_frame[6] [0]), .I3(n40132), .O(n26_adj_4179));
    defparam i11_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_960 (.I0(n42449), .I1(n42687), .I2(\data_in_frame[12] [0]), 
            .I3(\data_in_frame[11] [6]), .O(n24_adj_4180));
    defparam i9_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_961 (.I0(\data_in_frame[9] [6]), .I1(n42744), 
            .I2(n27639), .I3(n42483), .O(n25_adj_4181));
    defparam i10_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(\data_in_frame[10] [0]), .I1(n42880), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n23_adj_4182));
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut_adj_962 (.I0(n23_adj_4182), .I1(n25_adj_4181), .I2(n24_adj_4180), 
            .I3(n26_adj_4179), .O(n39681));
    defparam i14_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42252));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_964 (.I0(n42813), .I1(n42443), .I2(\data_in_frame[12] [3]), 
            .I3(n42894), .O(n10_adj_4183));
    defparam i4_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_965 (.I0(n42566), .I1(n10_adj_4183), .I2(n27347), 
            .I3(GND_net), .O(n39699));
    defparam i5_3_lut_adj_965.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[18] [6]), 
            .I2(n39681), .I3(n42594), .O(n42844));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1206));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_966 (.I0(n42690), .I1(n40241), .I2(n42437), .I3(\data_in_frame[9] [7]), 
            .O(n44461));
    defparam i3_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_967 (.I0(n42690), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[10] [1]), .O(n14_adj_4184));
    defparam i6_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_968 (.I0(\data_in_frame[14] [3]), .I1(n14_adj_4184), 
            .I2(n10_adj_4185), .I3(Kp_23__N_1206), .O(n44467));
    defparam i7_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_969 (.I0(n25058), .I1(n26858), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4186));
    defparam i2_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_970 (.I0(n7_adj_4186), .I1(n44467), .I2(\data_in_frame[18] [7]), 
            .I3(n44461), .O(n42906));
    defparam i4_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_971 (.I0(\data_in_frame[16] [6]), .I1(n42906), 
            .I2(GND_net), .I3(GND_net), .O(n42636));
    defparam i1_2_lut_adj_971.LUT_INIT = 16'h6666;
    SB_LUT4 i31761_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46714));
    defparam i31761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_972 (.I0(\data_in_frame[16] [5]), .I1(n42636), 
            .I2(\data_in_frame[14] [5]), .I3(n27041), .O(n26223));
    defparam i3_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i31762_4_lut (.I0(n46714), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n46715));
    defparam i31762_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i31760_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46713));
    defparam i31760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_973 (.I0(\data_in_frame[19] [1]), .I1(n26223), 
            .I2(GND_net), .I3(GND_net), .O(n42500));
    defparam i1_2_lut_adj_973.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_974 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4187));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_974.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_adj_975 (.I0(\FRAME_MATCHER.state [0]), .I1(n26622), 
            .I2(GND_net), .I3(GND_net), .O(n87));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_975.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_976 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4188));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_976.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_977 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4189));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_977.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_978 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_978.LUT_INIT = 16'h7bde;
    SB_LUT4 i2172853_i1_3_lut (.I0(n49338), .I1(n49332), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4190));
    defparam i2172853_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_979 (.I0(n9), .I1(n11_adj_4189), .I2(n10_adj_4188), 
            .I3(n12_adj_4187), .O(n24130));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i32841_2_lut (.I0(n49428), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47595));
    defparam i32841_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31722_4_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n46675));
    defparam i31722_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i33127_3_lut (.I0(n49398), .I1(n46675), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48080));
    defparam i33127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31755_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46708));
    defparam i31755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_980 (.I0(n42360), .I1(\data_in_frame[6] [7]), .I2(\data_in_frame[2] [6]), 
            .I3(\data_in_frame[4] [7]), .O(n10_adj_4191));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_981 (.I0(n42404), .I1(n10_adj_4191), .I2(\data_in_frame[7] [1]), 
            .I3(GND_net), .O(n10));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_982 (.I0(n10), .I1(n27417), .I2(GND_net), .I3(GND_net), 
            .O(Kp_23__N_1233));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_983 (.I0(n27438), .I1(\data_in_frame[11] [4]), 
            .I2(n42506), .I3(n6_adj_4192), .O(n40198));
    defparam i4_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42480));
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_985 (.I0(n40241), .I1(n27639), .I2(\data_in_frame[13] [7]), 
            .I3(n42449), .O(n10_adj_4193));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_986 (.I0(n42753), .I1(n42880), .I2(n44382), .I3(n42443), 
            .O(n12_adj_4194));
    defparam i5_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_987 (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[9] [1]), 
            .I2(n12_adj_4194), .I3(n8_adj_4195), .O(n42506));
    defparam i1_4_lut_adj_987.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4196));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_989 (.I0(\data_in_frame[16] [3]), .I1(n44467), 
            .I2(n42506), .I3(n6_adj_4196), .O(n42786));
    defparam i4_4_lut_adj_989.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_990 (.I0(n42357), .I1(n27438), .I2(\data_in_frame[16] [2]), 
            .I3(n40198), .O(n18_adj_4197));
    defparam i7_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_991 (.I0(\data_in_frame[11] [5]), .I1(n18_adj_4197), 
            .I2(\data_in_frame[18] [3]), .I3(\data_in_frame[14] [0]), .O(n20_adj_4198));
    defparam i9_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_992 (.I0(n42756), .I1(n20_adj_4198), .I2(n16_adj_4199), 
            .I3(\data_in_frame[13] [7]), .O(n42584));
    defparam i10_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_993 (.I0(n39681), .I1(n42506), .I2(\data_in_frame[14] [2]), 
            .I3(GND_net), .O(n44495));
    defparam i2_3_lut_adj_993.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_994 (.I0(\data_in_frame[18] [4]), .I1(n44495), 
            .I2(n42480), .I3(n40198), .O(n42580));
    defparam i3_4_lut_adj_994.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_995 (.I0(n42741), .I1(\data_in_frame[15] [6]), 
            .I2(n40652), .I3(n42865), .O(n10_adj_4200));
    defparam i4_4_lut_adj_995.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_996 (.I0(n42591), .I1(n10_adj_4200), .I2(n40524), 
            .I3(GND_net), .O(n40570));
    defparam i5_3_lut_adj_996.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_997 (.I0(n42825), .I1(\data_in_frame[20] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4201));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h6666;
    SB_LUT4 i31756_4_lut (.I0(n46708), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n46709));
    defparam i31756_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i31754_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46707));
    defparam i31754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[20] [7]), .I1(n40570), .I2(n42786), 
            .I3(GND_net), .O(n8_adj_4202));
    defparam i3_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_998 (.I0(Kp_23__N_761), .I1(n42613), .I2(n40570), 
            .I3(\data_in_frame[21] [1]), .O(n43997));
    defparam i3_4_lut_adj_998.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_999 (.I0(n40652), .I1(n8_adj_4202), .I2(\data_in_frame[19] [0]), 
            .I3(Kp_23__N_761), .O(n43562));
    defparam i4_4_lut_adj_999.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1000 (.I0(\data_in_frame[21] [5]), .I1(n42525), 
            .I2(n40504), .I3(\data_in_frame[19] [4]), .O(n44626));
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1001 (.I0(n42580), .I1(n42786), .I2(\data_in_frame[20] [6]), 
            .I3(GND_net), .O(n43581));
    defparam i2_3_lut_adj_1001.LUT_INIT = 16'h9696;
    SB_LUT4 i2173456_i1_3_lut (.I0(n49326), .I1(n49416), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4203));
    defparam i2173456_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1002 (.I0(\data_in_frame[20] [0]), .I1(n42491), 
            .I2(n44122), .I3(n39733), .O(n44455));
    defparam i3_4_lut_adj_1002.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1003 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[21] [6]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n6_adj_4204));
    defparam i2_3_lut_adj_1003.LUT_INIT = 16'h9696;
    SB_LUT4 i32835_2_lut (.I0(n49434), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47601));
    defparam i32835_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i21_4_lut (.I0(n42437), .I1(n40241), .I2(n40629), .I3(\data_in_frame[11] [2]), 
            .O(n50_adj_4205));
    defparam i21_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i31719_4_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n46672));
    defparam i31719_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i3_4_lut_adj_1004 (.I0(\data_in_frame[21] [2]), .I1(n42500), 
            .I2(n43998), .I3(\data_in_frame[19] [0]), .O(n44475));
    defparam i3_4_lut_adj_1004.LUT_INIT = 16'h9669;
    SB_LUT4 i33133_3_lut (.I0(n49392), .I1(n46672), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48086));
    defparam i33133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31749_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46702));
    defparam i31749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31750_4_lut (.I0(n46702), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n46703));
    defparam i31750_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i31748_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46701));
    defparam i31748_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(CLK_c), 
            .D(n41717), .S(n41769));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2174059_i1_3_lut (.I0(n49320), .I1(n49458), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4206));
    defparam i2174059_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32832_2_lut (.I0(n49440), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47604));
    defparam i32832_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31716_4_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n46669));
    defparam i31716_4_lut.LUT_INIT = 16'hc00a;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(CLK_c), 
            .D(n7_adj_4207), .S(n8_adj_4208));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(CLK_c), 
            .D(n41715), .S(n41771));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(CLK_c), 
            .D(n41713), .S(n41773));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(CLK_c), 
            .D(n41711), .S(n41775));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(CLK_c), 
            .D(n41709), .S(n41729));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(CLK_c), 
            .D(n41707), .S(n41725));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(CLK_c), 
            .D(n41705), .S(n41777));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(CLK_c), 
            .D(n7_adj_4209), .S(n41779));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(CLK_c), 
            .D(n41703), .S(n41781));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(CLK_c), 
            .D(n41701), .S(n41783));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1005 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[20] [2]), 
            .I2(n44122), .I3(GND_net), .O(n43666));
    defparam i2_3_lut_adj_1005.LUT_INIT = 16'h6969;
    SB_LUT4 i33139_3_lut (.I0(n49386), .I1(n46669), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48092));
    defparam i33139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31743_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46696));
    defparam i31743_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(CLK_c), 
            .D(n41699), .S(n41785));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(CLK_c), 
            .D(n41697), .S(n41787));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(CLK_c), 
            .D(n41695), .S(n41789));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(CLK_c), 
            .D(n41693), .S(n41791));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(CLK_c), 
            .D(n41691), .S(n41793));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(CLK_c), 
            .D(n41689), .S(n41743));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(CLK_c), 
            .D(n41687), .S(n41795));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(CLK_c), 
            .D(n41685), .S(n41797));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(CLK_c), 
            .D(n41683), .S(n41799));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(CLK_c), 
            .D(n41681), .S(n41741));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(CLK_c), 
            .D(n41679), .S(n41801));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(CLK_c), 
            .D(n41677), .S(n41803));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(CLK_c), 
            .D(n7_adj_4210), .S(n41739));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(CLK_c), 
            .D(n41675), .S(n41737));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(CLK_c), 
            .D(n41673), .S(n41805));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(CLK_c), 
            .D(n41671), .S(n41669));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n41665), .S(n41733));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31744_4_lut (.I0(n46696), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n46697));
    defparam i31744_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i31742_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46695));
    defparam i31742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1006 (.I0(n40235), .I1(\data_in_frame[18] [1]), 
            .I2(\data_in_frame[20] [3]), .I3(n42825), .O(n44775));
    defparam i2_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1007 (.I0(n40235), .I1(n42491), .I2(\data_in_frame[20] [1]), 
            .I3(GND_net), .O(n44445));
    defparam i2_3_lut_adj_1007.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1008 (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[19] [0]), 
            .I2(Kp_23__N_761), .I3(GND_net), .O(n7_adj_4211));
    defparam i2_3_lut_adj_1008.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1009 (.I0(n40502), .I1(\data_in_frame[19] [5]), 
            .I2(n39733), .I3(\data_in_frame[21] [7]), .O(n43715));
    defparam i3_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1010 (.I0(n42584), .I1(\data_in_frame[20] [5]), 
            .I2(n4_adj_4201), .I3(n42580), .O(n18_adj_4212));
    defparam i2_4_lut_adj_1010.LUT_INIT = 16'h7edb;
    SB_LUT4 i31661_4_lut (.I0(n43581), .I1(n44626), .I2(n43562), .I3(n43997), 
            .O(n46540));
    defparam i31661_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut_adj_1011 (.I0(n7_adj_4211), .I1(n43998), .I2(n40570), 
            .I3(n42613), .O(n44001));
    defparam i4_4_lut_adj_1011.LUT_INIT = 16'h9669;
    SB_LUT4 i31549_4_lut (.I0(n44455), .I1(n42525), .I2(n42768), .I3(\data_in_frame[21] [4]), 
            .O(n46427));
    defparam i31549_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_4_lut_adj_1012 (.I0(n43504), .I1(n40578), .I2(n6_adj_4204), 
            .I3(n40257), .O(n23_adj_4213));
    defparam i7_4_lut_adj_1012.LUT_INIT = 16'hbeeb;
    SB_LUT4 i11_4_lut_adj_1013 (.I0(n44445), .I1(n44775), .I2(n43666), 
            .I3(n44475), .O(n27_adj_4214));
    defparam i11_4_lut_adj_1013.LUT_INIT = 16'hfffb;
    SB_LUT4 i13_4_lut_adj_1014 (.I0(n44001), .I1(n46540), .I2(n18_adj_4212), 
            .I3(n43715), .O(n29));
    defparam i13_4_lut_adj_1014.LUT_INIT = 16'hfff7;
    SB_LUT4 i15_4_lut_adj_1015 (.I0(n29), .I1(n27_adj_4214), .I2(n23_adj_4213), 
            .I3(n46427), .O(n31_adj_4128));
    defparam i15_4_lut_adj_1015.LUT_INIT = 16'hfeff;
    SB_LUT4 i19_4_lut_adj_1016 (.I0(\data_in_frame[16] [5]), .I1(n42813), 
            .I2(n42915), .I3(n42732), .O(n48));
    defparam i19_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i2174662_i1_3_lut (.I0(n49314), .I1(n49482), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4215));
    defparam i2174662_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32830_2_lut (.I0(n49446), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47607));
    defparam i32830_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31713_4_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n46666));
    defparam i31713_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i33143_3_lut (.I0(n49380), .I1(n46666), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48096));
    defparam i33143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20_4_lut (.I0(n42677), .I1(n42594), .I2(n42657), .I3(n42480), 
            .O(n49_adj_4216));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31735_4_lut (.I0(\data_out_frame[6] [1]), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n46688));
    defparam i31735_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i31733_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46686));
    defparam i31733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32878_2_lut (.I0(n49452), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47611));
    defparam i32878_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31710_4_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n46663));
    defparam i31710_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i33147_3_lut (.I0(n49374), .I1(n46663), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48100));
    defparam i33147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31731_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46684));
    defparam i31731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31732_4_lut (.I0(n46684), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n46685));
    defparam i31732_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i31730_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n46683));
    defparam i31730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2176471_i1_3_lut (.I0(n49290), .I1(n49284), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4217));
    defparam i2176471_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32838_2_lut (.I0(n49464), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47617));
    defparam i32838_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31704_4_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n46657));
    defparam i31704_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i33151_3_lut (.I0(n49362), .I1(n46657), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48104));
    defparam i33151_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n27893), .D(n44563));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1017 (.I0(\data_in_frame[1] [4]), .I1(n26924), 
            .I2(n26870), .I3(\data_in_frame[1] [3]), .O(n42407));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1018 (.I0(n42591), .I1(n26858), .I2(\data_in_frame[14] [6]), 
            .I3(\data_in_frame[9] [3]), .O(n47));
    defparam i18_4_lut_adj_1018.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1019 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [10]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n43_adj_4218));   // verilog/coms.v(231[5:23])
    defparam i15_4_lut_adj_1019.LUT_INIT = 16'hfffe;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n27893), .D(n42611));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n27893), .D(n43933));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n27893), .D(n42625));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n27893), .D(n44321));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n27893), .D(n43986));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(CLK_c), 
            .E(n27893), .D(n42627));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(CLK_c), 
            .E(n27893), .D(n42905));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n27893), .D(n44856));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n27893), .D(n43837));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n27893), .D(n43664));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n27893), .D(n43918));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n27893), .D(n44471));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n27893), .D(n43603));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n27893), .D(n43527));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n27893), .D(n43931));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1020 (.I0(\data_out_frame[23] [6]), .I1(n42604), 
            .I2(n40634), .I3(GND_net), .O(n43931));
    defparam i2_3_lut_adj_1020.LUT_INIT = 16'h6969;
    SB_LUT4 i7_4_lut_adj_1021 (.I0(n42649), .I1(n14_adj_4219), .I2(n10_adj_4220), 
            .I3(n42497), .O(n43527));
    defparam i7_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1022 (.I0(n27210), .I1(n42551), .I2(\data_out_frame[23] [7]), 
            .I3(n39632), .O(n42497));
    defparam i3_4_lut_adj_1022.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_1023 (.I0(\data_in_frame[12] [1]), .I1(n42753), 
            .I2(n42918), .I3(n42665), .O(n46));
    defparam i17_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1024 (.I0(n31_adj_4128), .I1(n24130), .I2(n49), 
            .I3(GND_net), .O(n27752));
    defparam i2_3_lut_adj_1024.LUT_INIT = 16'h1010;
    SB_LUT4 i20_4_lut_adj_1025 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [7]), .I3(\FRAME_MATCHER.state [20]), 
            .O(n48_adj_4221));   // verilog/coms.v(231[5:23])
    defparam i20_4_lut_adj_1025.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1026 (.I0(\FRAME_MATCHER.state [11]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(\FRAME_MATCHER.state [26]), .I3(\FRAME_MATCHER.state [17]), 
            .O(n46_adj_4222));   // verilog/coms.v(231[5:23])
    defparam i18_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1027 (.I0(\FRAME_MATCHER.state [19]), .I1(\FRAME_MATCHER.state [24]), 
            .I2(\FRAME_MATCHER.state [9]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n47_adj_4223));   // verilog/coms.v(231[5:23])
    defparam i19_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1028 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [21]), 
            .I2(\FRAME_MATCHER.state [18]), .I3(\FRAME_MATCHER.state [8]), 
            .O(n45_adj_4224));   // verilog/coms.v(231[5:23])
    defparam i17_4_lut_adj_1028.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45_adj_4224), .I1(n47_adj_4223), .I2(n46_adj_4222), 
            .I3(n48_adj_4221), .O(n54));   // verilog/coms.v(231[5:23])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter_c[3]), 
            .I1(n48104), .I2(n47617), .I3(byte_transmit_counter_c[4]), 
            .O(n49515));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49515_bdd_4_lut (.I0(n49515), .I1(n14_adj_4217), .I2(n7_adj_4225), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[0]));
    defparam n49515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i21_4_lut_adj_1029 (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(\FRAME_MATCHER.state [29]), .I3(\FRAME_MATCHER.state [12]), 
            .O(n49_adj_4226));   // verilog/coms.v(231[5:23])
    defparam i21_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_34515 (.I0(byte_transmit_counter_c[3]), 
            .I1(n48100), .I2(n47611), .I3(byte_transmit_counter_c[4]), 
            .O(n49509));
    defparam byte_transmit_counter_3__bdd_4_lut_34515.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1030 (.I0(n40634), .I1(n42497), .I2(n26951), 
            .I3(GND_net), .O(n44471));
    defparam i2_3_lut_adj_1030.LUT_INIT = 16'h6969;
    SB_LUT4 i16_4_lut_adj_1031 (.I0(n42654), .I1(n26861), .I2(Kp_23__N_1402), 
            .I3(n42458), .O(n45_adj_4227));
    defparam i16_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1032 (.I0(n39632), .I1(\data_out_frame[24] [2]), 
            .I2(n44027), .I3(GND_net), .O(n43918));
    defparam i2_3_lut_adj_1032.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1033 (.I0(n27210), .I1(n42616), .I2(\data_out_frame[24] [3]), 
            .I3(GND_net), .O(n44027));
    defparam i2_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 n49509_bdd_4_lut (.I0(n49509), .I1(n49404), .I2(n7_adj_4228), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[1]));
    defparam n49509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4226), .I1(n54), .I2(n43_adj_4218), 
            .I3(n44_adj_4229), .O(n26622));   // verilog/coms.v(231[5:23])
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_34510 (.I0(byte_transmit_counter_c[3]), 
            .I1(n48096), .I2(n47607), .I3(byte_transmit_counter_c[4]), 
            .O(n49503));
    defparam byte_transmit_counter_3__bdd_4_lut_34510.LUT_INIT = 16'he4aa;
    SB_LUT4 n49503_bdd_4_lut (.I0(n49503), .I1(n14_adj_4215), .I2(n7_adj_4230), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[2]));
    defparam n49503_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_34505 (.I0(byte_transmit_counter_c[3]), 
            .I1(n48092), .I2(n47604), .I3(byte_transmit_counter_c[4]), 
            .O(n49497));
    defparam byte_transmit_counter_3__bdd_4_lut_34505.LUT_INIT = 16'he4aa;
    SB_LUT4 n49497_bdd_4_lut (.I0(n49497), .I1(n14_adj_4206), .I2(n7_adj_4231), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[3]));
    defparam n49497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_34500 (.I0(byte_transmit_counter_c[3]), 
            .I1(n48086), .I2(n47601), .I3(byte_transmit_counter_c[4]), 
            .O(n49491));
    defparam byte_transmit_counter_3__bdd_4_lut_34500.LUT_INIT = 16'he4aa;
    SB_LUT4 n49491_bdd_4_lut (.I0(n49491), .I1(n14_adj_4203), .I2(n7_adj_4232), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[4]));
    defparam n49491_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i33685_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n84));
    defparam i33685_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_34495 (.I0(byte_transmit_counter_c[3]), 
            .I1(n48080), .I2(n47595), .I3(byte_transmit_counter_c[4]), 
            .O(n49485));
    defparam byte_transmit_counter_3__bdd_4_lut_34495.LUT_INIT = 16'he4aa;
    SB_LUT4 n49485_bdd_4_lut (.I0(n49485), .I1(n14_adj_4190), .I2(n7_adj_4233), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[5]));
    defparam n49485_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1034 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n26622), .I3(GND_net), .O(n26482));
    defparam i2_3_lut_adj_1034.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n49479));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49479_bdd_4_lut (.I0(n49479), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n49482));
    defparam n49479_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_34490 (.I0(byte_transmit_counter_c[3]), 
            .I1(n48074), .I2(n47614), .I3(byte_transmit_counter_c[4]), 
            .O(n49473));
    defparam byte_transmit_counter_3__bdd_4_lut_34490.LUT_INIT = 16'he4aa;
    SB_LUT4 n49473_bdd_4_lut (.I0(n49473), .I1(n14_adj_4175), .I2(n7_adj_4234), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[6]));
    defparam n49473_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_34480 (.I0(byte_transmit_counter_c[3]), 
            .I1(n49260), .I2(n47592), .I3(byte_transmit_counter_c[4]), 
            .O(n49467));
    defparam byte_transmit_counter_3__bdd_4_lut_34480.LUT_INIT = 16'he4aa;
    SB_LUT4 n49467_bdd_4_lut (.I0(n49467), .I1(n14_adj_4174), .I2(n7_adj_4235), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[7]));
    defparam n49467_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34485 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n49461));
    defparam byte_transmit_counter_0__bdd_4_lut_34485.LUT_INIT = 16'he4aa;
    SB_LUT4 n49461_bdd_4_lut (.I0(n49461), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n49464));
    defparam n49461_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34471 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n49455));
    defparam byte_transmit_counter_0__bdd_4_lut_34471.LUT_INIT = 16'he4aa;
    SB_LUT4 n49455_bdd_4_lut (.I0(n49455), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n49458));
    defparam n49455_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34466 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n49449));
    defparam byte_transmit_counter_0__bdd_4_lut_34466.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_1035 (.I0(n42607), .I1(n27239), .I2(\data_out_frame[13] [4]), 
            .I3(\data_out_frame[19] [6]), .O(n14_adj_4236));
    defparam i6_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_4237), .S(n3_adj_4142));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4238), .S(n3_adj_4141));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4239), .S(n3_adj_4139));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4240), .S(n3_adj_4138));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_4241), .S(n3_adj_4137));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_4242), .S(n3_adj_4136));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_4243), .S(n3_adj_4135));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_4244), .S(n3_adj_4134));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_4245), .S(n3_adj_4133));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_4246), .S(n3_adj_4132));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_4247), .S(n3_adj_4129));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_4248), .S(n3_adj_4126));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_4249), .S(n3_adj_4120));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_4250), .S(n3_adj_4118));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_4251), .S(n3_adj_4117));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_4252), .S(n3_adj_4116));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_4253), .S(n3_adj_4115));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_4254), .S(n3_adj_4114));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_4255), .S(n3_adj_4113));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_4256), .S(n3_adj_4111));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_4257), .S(n3_adj_4110));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_4258), .S(n3_adj_4109));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_4259), .S(n3_adj_4260));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_4261), .S(n3_adj_4262));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4263), .S(n3_adj_4264));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4265), .S(n3_adj_4266));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4267), .S(n3_adj_4268));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4269), .S(n3_adj_4270));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_4271), .S(n3_adj_4272));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4273), .S(n3_adj_4274));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4119), .S(n3_adj_4275));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1036 (.I0(\data_out_frame[20] [0]), .I1(n14_adj_4236), 
            .I2(n10_adj_4276), .I3(n40554), .O(n27210));
    defparam i7_4_lut_adj_1036.LUT_INIT = 16'h9669;
    SB_LUT4 i27_4_lut_adj_1037 (.I0(n47), .I1(n49_adj_4216), .I2(n48), 
            .I3(n50_adj_4205), .O(n56));
    defparam i27_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 n49449_bdd_4_lut (.I0(n49449), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n49452));
    defparam n49449_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1038 (.I0(n52), .I1(\FRAME_MATCHER.i_31__N_2524 ), 
            .I2(n85), .I3(GND_net), .O(n2482));
    defparam i2_3_lut_adj_1038.LUT_INIT = 16'hdfdf;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34461 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n49443));
    defparam byte_transmit_counter_0__bdd_4_lut_34461.LUT_INIT = 16'he4aa;
    SB_LUT4 n49443_bdd_4_lut (.I0(n49443), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n49446));
    defparam n49443_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34456 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n49437));
    defparam byte_transmit_counter_0__bdd_4_lut_34456.LUT_INIT = 16'he4aa;
    SB_LUT4 n49437_bdd_4_lut (.I0(n49437), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n49440));
    defparam n49437_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34451 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n49431));
    defparam byte_transmit_counter_0__bdd_4_lut_34451.LUT_INIT = 16'he4aa;
    SB_LUT4 i22_4_lut (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[15] [4]), .I3(n30), .O(n51));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(\data_in_frame[18] [1]), .I1(n42825), 
            .I2(GND_net), .I3(GND_net), .O(n42535));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1040 (.I0(n42649), .I1(\data_out_frame[24] [5]), 
            .I2(n39689), .I3(n42903), .O(n44856));
    defparam i3_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 n49431_bdd_4_lut (.I0(n49431), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n49434));
    defparam n49431_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(\data_out_frame[24] [6]), .I1(n42903), 
            .I2(GND_net), .I3(GND_net), .O(n42905));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h6666;
    SB_LUT4 i4_3_lut (.I0(n42906), .I1(n42580), .I2(n42584), .I3(GND_net), 
            .O(n16_adj_4277));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1042 (.I0(n42786), .I1(n42535), .I2(n27196), 
            .I3(n42844), .O(n19_adj_4278));
    defparam i7_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n51), .I1(n56), .I2(n45_adj_4227), .I3(n46), 
            .O(n44066));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34446 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n49425));
    defparam byte_transmit_counter_0__bdd_4_lut_34446.LUT_INIT = 16'he4aa;
    SB_LUT4 i10_4_lut_adj_1043 (.I0(n19_adj_4278), .I1(n42633), .I2(n16_adj_4277), 
            .I3(n39630), .O(n22_adj_4279));
    defparam i10_4_lut_adj_1043.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1044 (.I0(n40073), .I1(n42834), .I2(\data_out_frame[25] [7]), 
            .I3(GND_net), .O(n42604));
    defparam i2_3_lut_adj_1044.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(n43940), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40668));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(n40114), .I1(n42645), .I2(GND_net), 
            .I3(GND_net), .O(n42646));
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26951));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1048 (.I0(n17_adj_4280), .I1(n22_adj_4279), .I2(\data_in_frame[16] [7]), 
            .I3(n44066), .O(n40524));
    defparam i11_4_lut_adj_1048.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(n40586), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42801));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h6666;
    SB_LUT4 n49425_bdd_4_lut (.I0(n49425), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n49428));
    defparam n49425_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1050 (.I0(n40283), .I1(\data_out_frame[19] [7]), 
            .I2(n42780), .I3(n6_adj_4281), .O(n26238));
    defparam i4_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(\data_out_frame[20] [1]), .I1(n26238), 
            .I2(GND_net), .I3(GND_net), .O(n42648));
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27181));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1053 (.I0(\data_out_frame[20] [1]), .I1(n42645), 
            .I2(\data_out_frame[20] [5]), .I3(GND_net), .O(n42550));
    defparam i2_3_lut_adj_1053.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1054 (.I0(n42541), .I1(n42550), .I2(\data_out_frame[17] [5]), 
            .I3(\data_out_frame[15] [4]), .O(n12_adj_4282));
    defparam i5_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1055 (.I0(n43940), .I1(n12_adj_4282), .I2(n42801), 
            .I3(n27679), .O(n40114));
    defparam i6_4_lut_adj_1055.LUT_INIT = 16'h9669;
    SB_LUT4 i21_4_lut_adj_1056 (.I0(n40114), .I1(n42790), .I2(\data_out_frame[23] [3]), 
            .I3(n42759), .O(n50_adj_4283));
    defparam i21_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1057 (.I0(n40658), .I1(n27181), .I2(\data_out_frame[24] [7]), 
            .I3(n42774), .O(n48_adj_4284));
    defparam i19_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1058 (.I0(\data_out_frame[23] [7]), .I1(n42886), 
            .I2(n26258), .I3(n42648), .O(n49_adj_4285));
    defparam i20_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1059 (.I0(n42312), .I1(n39689), .I2(n26951), 
            .I3(n42503), .O(n47_adj_4286));
    defparam i18_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(n39650), .I1(n42771), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_4287));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut_adj_1061 (.I0(n42588), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[25] [1]), .I3(\data_out_frame[24] [6]), 
            .O(n46_adj_4288));
    defparam i17_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1062 (.I0(n42486), .I1(\data_out_frame[24] [3]), 
            .I2(n42604), .I3(n42625), .O(n45_adj_4289));
    defparam i16_4_lut_adj_1062.LUT_INIT = 16'h9669;
    SB_LUT4 i27_4_lut_adj_1063 (.I0(n47_adj_4286), .I1(n49_adj_4285), .I2(n48_adj_4284), 
            .I3(n50_adj_4283), .O(n56_adj_4290));
    defparam i27_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1064 (.I0(n42522), .I1(n42646), .I2(n40668), 
            .I3(n30_adj_4287), .O(n51_adj_4291));
    defparam i22_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut_adj_1065 (.I0(n51_adj_4291), .I1(n56_adj_4290), .I2(n45_adj_4289), 
            .I3(n46_adj_4288), .O(n42627));
    defparam i28_4_lut_adj_1065.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1066 (.I0(n40524), .I1(n40570), .I2(\data_in_frame[19] [7]), 
            .I3(GND_net), .O(n42491));
    defparam i2_3_lut_adj_1066.LUT_INIT = 16'h6969;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(CLK_c), .E(n12_adj_4164), .D(n27998), 
            .R(n43465));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1067 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n42519));
    defparam i2_3_lut_adj_1067.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1068 (.I0(n40517), .I1(\data_out_frame[15] [4]), 
            .I2(n42519), .I3(n6_adj_4292), .O(n26258));
    defparam i4_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1069 (.I0(n33507), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n42206));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1069.LUT_INIT = 16'hffdf;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34441 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n49419));
    defparam byte_transmit_counter_0__bdd_4_lut_34441.LUT_INIT = 16'he4aa;
    SB_LUT4 n49419_bdd_4_lut (.I0(n49419), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n49422));
    defparam n49419_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34436 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n49413));
    defparam byte_transmit_counter_0__bdd_4_lut_34436.LUT_INIT = 16'he4aa;
    SB_LUT4 n49413_bdd_4_lut (.I0(n49413), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n49416));
    defparam n49413_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n46632), .I2(n46633), .I3(byte_transmit_counter[2]), .O(n49401));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49401_bdd_4_lut (.I0(n49401), .I1(n46642), .I2(n46641), .I3(byte_transmit_counter[2]), 
            .O(n49404));
    defparam n49401_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34431 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n49395));
    defparam byte_transmit_counter_0__bdd_4_lut_34431.LUT_INIT = 16'he4aa;
    SB_LUT4 n49395_bdd_4_lut (.I0(n49395), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n49398));
    defparam n49395_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34416 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n49389));
    defparam byte_transmit_counter_0__bdd_4_lut_34416.LUT_INIT = 16'he4aa;
    SB_LUT4 n49389_bdd_4_lut (.I0(n49389), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n49392));
    defparam n49389_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34411 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n49383));
    defparam byte_transmit_counter_0__bdd_4_lut_34411.LUT_INIT = 16'he4aa;
    SB_LUT4 n49383_bdd_4_lut (.I0(n49383), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n49386));
    defparam n49383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34406 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n49377));
    defparam byte_transmit_counter_0__bdd_4_lut_34406.LUT_INIT = 16'he4aa;
    SB_LUT4 n49377_bdd_4_lut (.I0(n49377), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n49380));
    defparam n49377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_out_frame[20] [2]), .I1(n26258), 
            .I2(GND_net), .I3(GND_net), .O(n42312));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 i1418_2_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2206));   // verilog/coms.v(78[16:27])
    defparam i1418_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1071 (.I0(n44460), .I1(n27517), .I2(n2206), .I3(n39761), 
            .O(n42774));
    defparam i3_4_lut_adj_1071.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1072 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n26774));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_out_frame[23] [0]), .I1(n42774), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4293));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1074 (.I0(n40052), .I1(n40673), .I2(n42513), 
            .I3(n6_adj_4293), .O(n39650));
    defparam i4_4_lut_adj_1074.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1075 (.I0(n39650), .I1(n42840), .I2(n42699), 
            .I3(\data_out_frame[24] [6]), .O(n43986));
    defparam i3_4_lut_adj_1075.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1076 (.I0(\data_out_frame[24] [7]), .I1(n42601), 
            .I2(GND_net), .I3(GND_net), .O(n40052));
    defparam i1_2_lut_adj_1076.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(n26235), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42378));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1078 (.I0(n42735), .I1(n40033), .I2(n27223), 
            .I3(n27569), .O(n23_adj_4294));
    defparam i9_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34401 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18]_c [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n49371));
    defparam byte_transmit_counter_0__bdd_4_lut_34401.LUT_INIT = 16'he4aa;
    SB_LUT4 n49371_bdd_4_lut (.I0(n49371), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n49374));
    defparam n49371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_1079 (.I0(\data_out_frame[18]_c [1]), .I1(n1794), 
            .I2(n27321), .I3(n27679), .O(n22_adj_4295));
    defparam i8_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1080 (.I0(n23_adj_4294), .I1(n42378), .I2(n20_adj_4296), 
            .I3(n40582), .O(n26_adj_4297));
    defparam i12_4_lut_adj_1080.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34391 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n49359));
    defparam byte_transmit_counter_0__bdd_4_lut_34391.LUT_INIT = 16'he4aa;
    SB_LUT4 n49359_bdd_4_lut (.I0(n49359), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n49362));
    defparam n49359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34386 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n49335));
    defparam byte_transmit_counter_0__bdd_4_lut_34386.LUT_INIT = 16'he4aa;
    SB_LUT4 n49335_bdd_4_lut (.I0(n49335), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n49338));
    defparam n49335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34367 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n49329));
    defparam byte_transmit_counter_0__bdd_4_lut_34367.LUT_INIT = 16'he4aa;
    SB_LUT4 n49329_bdd_4_lut (.I0(n49329), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n49332));
    defparam n49329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34362 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n49323));
    defparam byte_transmit_counter_0__bdd_4_lut_34362.LUT_INIT = 16'he4aa;
    SB_LUT4 i13_4_lut_adj_1081 (.I0(n40512), .I1(n26_adj_4297), .I2(n22_adj_4295), 
            .I3(n40576), .O(n42783));
    defparam i13_4_lut_adj_1081.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1082 (.I0(\data_out_frame[18] [2]), .I1(n42783), 
            .I2(n42553), .I3(n42241), .O(n39724));
    defparam i3_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42246));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_LUT4 n49323_bdd_4_lut (.I0(n49323), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n49326));
    defparam n49323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(n39724), .I1(n24914), .I2(GND_net), 
            .I3(GND_net), .O(n42522));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1085 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[4] [6]), 
            .I2(n27337), .I3(n27340), .O(n12_adj_4298));   // verilog/coms.v(236[9:81])
    defparam i5_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n37283), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n37282), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_8 (.CI(n37282), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n37283));
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n37281), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1086 (.I0(\data_in_frame[7] [0]), .I1(n12_adj_4298), 
            .I2(n26774), .I3(\data_in_frame[6] [7]), .O(n26969));   // verilog/coms.v(236[9:81])
    defparam i6_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1087 (.I0(n2063), .I1(n39642), .I2(\data_out_frame[23] [1]), 
            .I3(GND_net), .O(n42886));
    defparam i2_3_lut_adj_1087.LUT_INIT = 16'h9696;
    SB_CARRY add_3971_7 (.CI(n37281), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n37282));
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter_c[4]), 
            .I2(GND_net), .I3(n37280), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1088 (.I0(\data_out_frame[25] [2]), .I1(n39761), 
            .I2(n42777), .I3(n6_adj_4299), .O(n44321));
    defparam i4_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1089 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[16] [0]), .I3(GND_net), .O(n27569));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1089.LUT_INIT = 16'h9696;
    SB_LUT4 i33551_2_lut (.I0(n27113), .I1(\data_out_frame[13] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n48504));   // verilog/coms.v(97[12:26])
    defparam i33551_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3971_6 (.CI(n37280), .I0(byte_transmit_counter_c[4]), .I1(GND_net), 
            .CO(n37281));
    SB_LUT4 i3_4_lut_adj_1090 (.I0(n26235), .I1(n27569), .I2(\data_out_frame[13] [6]), 
            .I3(n48504), .O(n42241));
    defparam i3_4_lut_adj_1090.LUT_INIT = 16'h9669;
    SB_LUT4 i33555_3_lut (.I0(n42241), .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[16] [2]), 
            .I3(GND_net), .O(n48508));
    defparam i33555_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(n37279), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1091 (.I0(\data_out_frame[18] [2]), .I1(n40582), 
            .I2(n48508), .I3(n6_adj_4300), .O(n24914));
    defparam i3_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1092 (.I0(n44460), .I1(\data_out_frame[20] [4]), 
            .I2(n42274), .I3(n6_adj_4301), .O(n42462));
    defparam i4_4_lut_adj_1092.LUT_INIT = 16'h9669;
    SB_CARRY add_3971_5 (.CI(n37279), .I0(byte_transmit_counter_c[3]), .I1(GND_net), 
            .CO(n37280));
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n37278), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1093 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42759));
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4302));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1095 (.I0(n42759), .I1(n42462), .I2(n43813), 
            .I3(n6_adj_4302), .O(n42625));
    defparam i4_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_4 (.CI(n37278), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n37279));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n37277), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1096 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(n42639), .I3(n6_adj_4303), .O(n40512));
    defparam i4_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_out_frame[16] [1]), .I1(n40512), 
            .I2(GND_net), .I3(GND_net), .O(n42553));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_out_frame[20] [6]), .I1(n43813), 
            .I2(GND_net), .I3(GND_net), .O(n42274));
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1099 (.I0(\data_out_frame[18] [4]), .I1(n42804), 
            .I2(n42553), .I3(n40576), .O(n2063));
    defparam i3_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_3 (.CI(n37277), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n37278));
    SB_LUT4 i3_4_lut_adj_1100 (.I0(\data_out_frame[25] [3]), .I1(n42831), 
            .I2(n42601), .I3(\data_out_frame[23] [1]), .O(n43933));
    defparam i3_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1101 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n26838));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1101.LUT_INIT = 16'h9696;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3413), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut_adj_1102 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[11] [6]), .I3(n10_adj_4304), .O(n16_adj_4305));
    defparam i7_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3413), .CO(n37277));
    SB_LUT4 i8_4_lut_adj_1103 (.I0(n42816), .I1(n16_adj_4305), .I2(n12_adj_4306), 
            .I3(\data_out_frame[5] [2]), .O(n6_adj_4300));
    defparam i8_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_33_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n37276), .O(n2_adj_4237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1104 (.I0(n42559), .I1(n1673), .I2(\data_out_frame[13] [6]), 
            .I3(n42762), .O(n10_adj_4307));
    defparam i4_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1105 (.I0(n1516), .I1(n10_adj_4307), .I2(n1513), 
            .I3(GND_net), .O(n40582));
    defparam i5_3_lut_adj_1105.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_out_frame[20] [6]), .I1(n42513), 
            .I2(GND_net), .I3(GND_net), .O(n42777));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_32_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n37275), .O(n2_adj_4238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1107 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n27360));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1107.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1108 (.I0(n27360), .I1(\data_in_frame[4] [4]), 
            .I2(n26838), .I3(GND_net), .O(n27337));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1108.LUT_INIT = 16'h9696;
    SB_CARRY add_43_32 (.CI(n37275), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n37276));
    SB_LUT4 i1_2_lut_adj_1109 (.I0(n42486), .I1(n42610), .I2(GND_net), 
            .I3(GND_net), .O(n42611));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h9999;
    SB_LUT4 add_43_31_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n37274), .O(n2_adj_4239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1110 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [4]), .I3(GND_net), .O(n41671));
    defparam i1_2_lut_3_lut_adj_1110.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1111 (.I0(\data_in_frame[2] [1]), .I1(n27340), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[4] [4]), .O(n42724));   // verilog/coms.v(70[16:69])
    defparam i3_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1112 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [5]), .I3(GND_net), .O(n41673));
    defparam i1_2_lut_3_lut_adj_1112.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_31 (.CI(n37274), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n37275));
    SB_LUT4 add_43_30_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n37273), .O(n2_adj_4240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1113 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [6]), .I3(GND_net), .O(n41675));
    defparam i1_2_lut_3_lut_adj_1113.LUT_INIT = 16'he0e0;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n28189));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_30 (.CI(n37273), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n37274));
    SB_LUT4 add_43_29_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n37272), .O(n2_adj_4241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1114 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [7]), .I3(GND_net), .O(n7_adj_4210));
    defparam i1_2_lut_3_lut_adj_1114.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1115 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [8]), .I3(GND_net), .O(n41677));
    defparam i1_2_lut_3_lut_adj_1115.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42455));
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1117 (.I0(\data_out_frame[8] [2]), .I1(n42455), 
            .I2(n42765), .I3(\data_out_frame[8] [1]), .O(n18_adj_4310));
    defparam i7_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1118 (.I0(\data_out_frame[10] [3]), .I1(n18_adj_4310), 
            .I2(n42559), .I3(n42909), .O(n20_adj_4311));
    defparam i9_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1119 (.I0(n42847), .I1(n20_adj_4311), .I2(n16_adj_4312), 
            .I3(n42598), .O(n40576));
    defparam i10_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1120 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[18] [5]), .I3(\data_out_frame[18] [4]), 
            .O(n42494));
    defparam i3_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1121 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n42735));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1122 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42804));
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1123 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n42607));
    defparam i2_3_lut_adj_1123.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1124 (.I0(n43610), .I1(n42607), .I2(n27554), 
            .I3(n40554), .O(n43940));
    defparam i3_4_lut_adj_1124.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1125 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [9]), .I3(GND_net), .O(n41679));
    defparam i1_2_lut_3_lut_adj_1125.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(n40586), .I1(n42286), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4313));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1127 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(n6_adj_4313), .O(n43610));
    defparam i4_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1128 (.I0(\data_out_frame[19] [4]), .I1(n27128), 
            .I2(n43610), .I3(GND_net), .O(n42465));
    defparam i1_3_lut_adj_1128.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1129 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [10]), .I3(GND_net), .O(n41681));
    defparam i1_2_lut_3_lut_adj_1129.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n27239));
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_CARRY add_43_29 (.CI(n37272), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n37273));
    SB_LUT4 i1_2_lut_3_lut_adj_1131 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [11]), .I3(GND_net), .O(n41683));
    defparam i1_2_lut_3_lut_adj_1131.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_28_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n37271), .O(n2_adj_4242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1132 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[11] [5]), 
            .I2(n42877), .I3(n40283), .O(n42639));
    defparam i1_4_lut_adj_1132.LUT_INIT = 16'h9669;
    SB_CARRY add_43_28 (.CI(n37271), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n37272));
    SB_LUT4 i1_2_lut_3_lut_adj_1133 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [12]), .I3(GND_net), .O(n41685));
    defparam i1_2_lut_3_lut_adj_1133.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_27_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n37270), .O(n2_adj_4243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_27 (.CI(n37270), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n37271));
    SB_LUT4 i1_2_lut_3_lut_adj_1134 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [13]), .I3(GND_net), .O(n41687));
    defparam i1_2_lut_3_lut_adj_1134.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1135 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [14]), .I3(GND_net), .O(n41689));
    defparam i1_2_lut_3_lut_adj_1135.LUT_INIT = 16'he0e0;
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n28188));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_26_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n37269), .O(n2_adj_4244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1136 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [15]), .I3(GND_net), .O(n41691));
    defparam i1_2_lut_3_lut_adj_1136.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1137 (.I0(n42674), .I1(n27705), .I2(\data_out_frame[12] [7]), 
            .I3(\data_out_frame[8] [4]), .O(n14_adj_4314));
    defparam i6_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1138 (.I0(\data_out_frame[13] [1]), .I1(n14_adj_4314), 
            .I2(n10_adj_4315), .I3(n27215), .O(n40586));
    defparam i7_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1139 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n42897));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1139.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1140 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[13] [2]), 
            .I2(n42277), .I3(\data_out_frame[8] [6]), .O(n16_adj_4316));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42367));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1142 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(n42668), .I3(\data_out_frame[10] [6]), .O(n17_adj_4317));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1143 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [16]), .I3(GND_net), .O(n41693));
    defparam i1_2_lut_3_lut_adj_1143.LUT_INIT = 16'he0e0;
    SB_LUT4 i9_4_lut_adj_1144 (.I0(n17_adj_4317), .I1(\data_out_frame[8] [5]), 
            .I2(n16_adj_4316), .I3(n27547), .O(n27554));   // verilog/coms.v(74[16:43])
    defparam i9_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1145 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [17]), .I3(GND_net), .O(n41695));
    defparam i1_2_lut_3_lut_adj_1145.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1146 (.I0(n42874), .I1(\data_out_frame[9] [1]), 
            .I2(n26939), .I3(\data_out_frame[9] [3]), .O(n14_adj_4318));
    defparam i6_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1147 (.I0(\data_out_frame[13] [5]), .I1(n14_adj_4318), 
            .I2(n10_adj_4319), .I3(\data_out_frame[5] [1]), .O(n40283));
    defparam i7_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1148 (.I0(n27492), .I1(n42718), .I2(\data_out_frame[13] [3]), 
            .I3(\data_out_frame[9] [1]), .O(n12_adj_4320));
    defparam i5_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1149 (.I0(n27627), .I1(n12_adj_4320), .I2(n42793), 
            .I3(n27705), .O(n27679));
    defparam i6_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(n40283), .I1(n27554), .I2(GND_net), 
            .I3(GND_net), .O(n42622));
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1151 (.I0(\data_out_frame[11] [5]), .I1(n27121), 
            .I2(n42338), .I3(n6_adj_4321), .O(n27113));
    defparam i4_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1152 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [18]), .I3(GND_net), .O(n41697));
    defparam i1_2_lut_3_lut_adj_1152.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_26 (.CI(n37269), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n37270));
    SB_LUT4 add_43_25_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n37268), .O(n2_adj_4245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34357 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n49317));
    defparam byte_transmit_counter_0__bdd_4_lut_34357.LUT_INIT = 16'he4aa;
    SB_LUT4 n49317_bdd_4_lut (.I0(n49317), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n49320));
    defparam n49317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34352 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n49311));
    defparam byte_transmit_counter_0__bdd_4_lut_34352.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1153 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [19]), .I3(GND_net), .O(n41699));
    defparam i1_2_lut_3_lut_adj_1153.LUT_INIT = 16'he0e0;
    SB_LUT4 n49311_bdd_4_lut (.I0(n49311), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n49314));
    defparam n49311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1154 (.I0(n42856), .I1(n42912), .I2(\data_out_frame[11] [0]), 
            .I3(GND_net), .O(n42674));
    defparam i2_3_lut_adj_1154.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1155 (.I0(n42674), .I1(n40604), .I2(\data_out_frame[11] [5]), 
            .I3(n42853), .O(n10_adj_4322));
    defparam i4_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1156 (.I0(n42452), .I1(n1519), .I2(n9_adj_4323), 
            .I3(n10_adj_4322), .O(n42559));
    defparam i2_4_lut_adj_1156.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1157 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [20]), .I3(GND_net), .O(n41701));
    defparam i1_2_lut_3_lut_adj_1157.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34347 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n49305));
    defparam byte_transmit_counter_0__bdd_4_lut_34347.LUT_INIT = 16'he4aa;
    SB_LUT4 n49305_bdd_4_lut (.I0(n49305), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n49308));
    defparam n49305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_out_frame[8] [7]), .I1(n27666), 
            .I2(GND_net), .I3(GND_net), .O(n42718));
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1159 (.I0(n42331), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n42338));   // verilog/coms.v(71[16:62])
    defparam i2_3_lut_adj_1159.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27627));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4324));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1162 (.I0(\data_out_frame[12] [4]), .I1(n1668), 
            .I2(\data_out_frame[12] [5]), .I3(n6_adj_4324), .O(n42364));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_out_frame[12] [1]), .I1(n42364), 
            .I2(GND_net), .I3(GND_net), .O(n1673));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1164 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(n42711), .I3(n27492), .O(n10_adj_4325));   // verilog/coms.v(73[16:34])
    defparam i4_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1165 (.I0(n27498), .I1(n42877), .I2(n40604), 
            .I3(\data_out_frame[11] [0]), .O(n12_adj_4326));   // verilog/coms.v(75[16:43])
    defparam i5_4_lut_adj_1165.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1166 (.I0(n1673), .I1(n12_adj_4326), .I2(n1522), 
            .I3(n42853), .O(n42452));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1167 (.I0(n42238), .I1(n27705), .I2(\data_out_frame[6] [6]), 
            .I3(n42708), .O(n10_adj_4327));
    defparam i4_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1168 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [21]), .I3(GND_net), .O(n41703));
    defparam i1_2_lut_3_lut_adj_1168.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1169 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [22]), .I3(GND_net), .O(n7_adj_4209));
    defparam i1_2_lut_3_lut_adj_1169.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_adj_1170 (.I0(n27547), .I1(n10_adj_4327), .I2(\data_out_frame[11] [2]), 
            .I3(GND_net), .O(n26235));
    defparam i5_3_lut_adj_1170.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut_adj_1171 (.I0(n26235), .I1(\data_out_frame[12] [7]), 
            .I2(n42452), .I3(\data_out_frame[14] [2]), .O(n36));
    defparam i13_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1172 (.I0(n40517), .I1(n27113), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[13] [6]), .O(n34));
    defparam i11_4_lut_adj_1172.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_1173 (.I0(n42431), .I1(\data_out_frame[12] [5]), 
            .I2(n42243), .I3(\data_out_frame[12] [0]), .O(n39_adj_4328));
    defparam i16_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1174 (.I0(\data_out_frame[14] [6]), .I1(n42559), 
            .I2(\data_out_frame[14] [7]), .I3(n42468), .O(n38_adj_4329));
    defparam i15_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1175 (.I0(n42510), .I1(\data_out_frame[14] [1]), 
            .I2(n42302), .I3(n40586), .O(n37));
    defparam i14_4_lut_adj_1175.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34342 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n49299));
    defparam byte_transmit_counter_0__bdd_4_lut_34342.LUT_INIT = 16'he4aa;
    SB_LUT4 n49299_bdd_4_lut (.I0(n49299), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n49302));
    defparam n49299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i18_4_lut_adj_1176 (.I0(n27278), .I1(n36), .I2(n40530), .I3(n42639), 
            .O(n41_adj_4330));
    defparam i18_4_lut_adj_1176.LUT_INIT = 16'h9669;
    SB_LUT4 i20_4_lut_adj_1177 (.I0(n39_adj_4328), .I1(\data_out_frame[13] [0]), 
            .I2(n34), .I3(n26822), .O(n43_adj_4331));
    defparam i20_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1178 (.I0(n43_adj_4331), .I1(n41_adj_4330), .I2(n37), 
            .I3(n38_adj_4329), .O(n44221));
    defparam i22_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_996), 
            .I2(GND_net), .I3(GND_net), .O(n42388));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1180 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [23]), .I3(GND_net), .O(n41705));
    defparam i1_2_lut_3_lut_adj_1180.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1181 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [24]), .I3(GND_net), .O(n41707));
    defparam i1_2_lut_3_lut_adj_1181.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1182 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [25]), .I3(GND_net), .O(n41709));
    defparam i1_2_lut_3_lut_adj_1182.LUT_INIT = 16'he0e0;
    SB_LUT4 i14_4_lut_adj_1183 (.I0(\data_out_frame[18]_c [1]), .I1(n44221), 
            .I2(\data_out_frame[18] [2]), .I3(n42897), .O(n36_adj_4332));
    defparam i14_4_lut_adj_1183.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1184 (.I0(n42465), .I1(\data_out_frame[19] [2]), 
            .I2(n42822), .I3(n42642), .O(n34_adj_4333));
    defparam i12_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1185 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [26]), .I3(GND_net), .O(n41711));
    defparam i1_2_lut_3_lut_adj_1185.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1186 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [27]), .I3(GND_net), .O(n41713));
    defparam i1_2_lut_3_lut_adj_1186.LUT_INIT = 16'he0e0;
    SB_LUT4 i18_4_lut_adj_1187 (.I0(\data_out_frame[16] [1]), .I1(n36_adj_4332), 
            .I2(n26_adj_4334), .I3(n43940), .O(n40_adj_4335));
    defparam i18_4_lut_adj_1187.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_1188 (.I0(n42302), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[19] [3]), .I3(\data_out_frame[19] [6]), 
            .O(n38_adj_4336));
    defparam i16_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1189 (.I0(\data_out_frame[16] [0]), .I1(n40_adj_4335), 
            .I2(n34_adj_4333), .I3(\data_out_frame[18] [0]), .O(n42_adj_4337));
    defparam i20_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1190 (.I0(n42804), .I1(n42622), .I2(n42735), 
            .I3(n42494), .O(n37_adj_4338));
    defparam i15_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1191 (.I0(n37_adj_4338), .I1(n42576), .I2(n42_adj_4337), 
            .I3(n38_adj_4336), .O(n42819));
    defparam i1_4_lut_adj_1191.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1192 (.I0(n40033), .I1(n42819), .I2(\data_out_frame[16] [5]), 
            .I3(GND_net), .O(n27517));
    defparam i2_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1193 (.I0(n40576), .I1(n27321), .I2(\data_out_frame[18][6] ), 
            .I3(n42513), .O(n12_adj_4339));
    defparam i5_4_lut_adj_1193.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1194 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [28]), .I3(GND_net), .O(n41715));
    defparam i1_2_lut_3_lut_adj_1194.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1195 (.I0(\data_out_frame[16] [3]), .I1(n12_adj_4339), 
            .I2(n42819), .I3(\data_out_frame[18] [5]), .O(n40673));
    defparam i6_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1196 (.I0(n40673), .I1(n27517), .I2(\data_out_frame[20] [7]), 
            .I3(GND_net), .O(n43813));
    defparam i2_3_lut_adj_1196.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(n43813), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42588));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1198 (.I0(n40598), .I1(n42513), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n40073));
    defparam i2_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42822));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1200 (.I0(n1794), .I1(n42807), .I2(\data_out_frame[18] [7]), 
            .I3(GND_net), .O(n42576));
    defparam i2_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(85[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1201 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [29]), .I3(GND_net), .O(n7_adj_4207));
    defparam i1_2_lut_3_lut_adj_1201.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42868));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1203 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [30]), .I3(GND_net), .O(n41717));
    defparam i1_2_lut_3_lut_adj_1203.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1204 (.I0(n42277), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n42912));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1204.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42394));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1206 (.I0(n1_adj_4308), .I1(n1_adj_4309), 
            .I2(\FRAME_MATCHER.state [31]), .I3(GND_net), .O(n41649));
    defparam i1_2_lut_3_lut_adj_1206.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42696));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1208 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n27215));
    defparam i2_3_lut_adj_1208.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1209 (.I0(\data_out_frame[4] [1]), .I1(n42394), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[6] [4]), .O(n27406));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42816));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42668));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42243));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1213 (.I0(n26702), .I1(n1191), .I2(n42243), .I3(\data_out_frame[5] [1]), 
            .O(n42331));   // verilog/coms.v(73[16:34])
    defparam i3_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_CARRY add_43_25 (.CI(n37268), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n37269));
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26981));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1215 (.I0(\data_in_frame[8] [6]), .I1(Kp_23__N_1095), 
            .I2(\data_in_frame[8] [7]), .I3(GND_net), .O(n42269));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1215.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n28187));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1216 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n42262));
    defparam i2_3_lut_adj_1216.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4340));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1218 (.I0(n42488), .I1(\data_out_frame[10] [4]), 
            .I2(\data_out_frame[10] [1]), .I3(n6_adj_4340), .O(n42544));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_out_frame[10] [7]), .I1(n27406), 
            .I2(GND_net), .I3(GND_net), .O(n42793));
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(n2_adj_4341), .I1(n4_adj_4342), .I2(n1_adj_4308), 
            .I3(\FRAME_MATCHER.state [3]), .O(n7_adj_4343));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n28186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n28185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n28184));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_4_lut (.I0(n63_adj_4159), .I1(n771), .I2(n2_adj_4344), 
            .I3(n85), .O(n5_adj_4345));   // verilog/coms.v(157[6] 159[9])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'ha0a2;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n28183));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_24_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n37267), .O(n2_adj_4246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n37267), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n37268));
    SB_LUT4 add_43_23_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n37266), .O(n2_adj_4247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n37266), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n37267));
    SB_LUT4 i3_4_lut_adj_1220 (.I0(\data_out_frame[10] [5]), .I1(n42793), 
            .I2(n42544), .I3(n40542), .O(n40604));
    defparam i3_4_lut_adj_1220.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1221 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[5] [4]), .I3(n42816), .O(n36_adj_4346));   // verilog/coms.v(75[16:27])
    defparam i13_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_22_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n37265), .O(n2_adj_4248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_22 (.CI(n37265), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n37266));
    SB_LUT4 i11_3_lut_adj_1222 (.I0(n42262), .I1(\data_out_frame[6] [6]), 
            .I2(n27492), .I3(GND_net), .O(n34_adj_4347));   // verilog/coms.v(75[16:27])
    defparam i11_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_21_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n37264), .O(n2_adj_4249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_21 (.CI(n37264), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n37265));
    SB_LUT4 add_43_20_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n37263), .O(n2_adj_4250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n37263), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n37264));
    SB_LUT4 i1_2_lut_3_lut_adj_1223 (.I0(n63_adj_4159), .I1(n771), .I2(n92[1]), 
            .I3(GND_net), .O(n27_adj_4348));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_3_lut_adj_1223.LUT_INIT = 16'hfdfd;
    SB_LUT4 add_43_19_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n37262), .O(n2_adj_4251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16_4_lut_adj_1224 (.I0(n42394), .I1(n42912), .I2(\data_out_frame[7] [1]), 
            .I3(n42868), .O(n39_adj_4349));   // verilog/coms.v(75[16:27])
    defparam i16_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1225 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [3]), 
            .I2(n27594), .I3(\data_in_frame[11] [3]), .O(n42385));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1226 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [3]), 
            .I2(Kp_23__N_1206), .I3(n10_adj_4193), .O(n44382));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1227 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [3]), 
            .I2(n42668), .I3(n42862), .O(n38_adj_4350));   // verilog/coms.v(75[16:27])
    defparam i15_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1228 (.I0(n42563), .I1(n42874), .I2(\data_out_frame[9] [1]), 
            .I3(n27406), .O(n37_adj_4351));   // verilog/coms.v(75[16:27])
    defparam i14_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1229 (.I0(\data_out_frame[8] [2]), .I1(n36_adj_4346), 
            .I2(\data_out_frame[9] [6]), .I3(n42572), .O(n41_adj_4352));   // verilog/coms.v(75[16:27])
    defparam i18_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1230 (.I0(n39_adj_4349), .I1(n42810), .I2(n34_adj_4347), 
            .I3(n42397), .O(n43_adj_4353));   // verilog/coms.v(75[16:27])
    defparam i20_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1231 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_1210), .I3(\data_in_frame[11] [2]), .O(n42705));   // verilog/coms.v(72[16:41])
    defparam i3_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42255));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1233 (.I0(n42407), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n42750));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1234 (.I0(n42426), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[7] [3]), .I3(n27200), .O(n10_adj_4354));
    defparam i4_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1235 (.I0(n43_adj_4353), .I1(n41_adj_4352), .I2(n37_adj_4351), 
            .I3(n38_adj_4350), .O(n40542));   // verilog/coms.v(75[16:27])
    defparam i22_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(n40542), .I1(n40604), .I2(GND_net), 
            .I3(GND_net), .O(n40112));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1237 (.I0(n42680), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4355));
    defparam i2_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1238 (.I0(n42859), .I1(n40112), .I2(n42651), 
            .I3(\data_out_frame[10] [7]), .O(n14_adj_4356));
    defparam i6_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1239 (.I0(n1668), .I1(n14_adj_4356), .I2(n10_adj_4355), 
            .I3(n42235), .O(n40530));
    defparam i7_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n28738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n28737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n28736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n28735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n28734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n28733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n28732));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1240 (.I0(n40530), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40554));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42302));
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1242 (.I0(\data_out_frame[17] [2]), .I1(n42302), 
            .I2(n27324), .I3(n40554), .O(n27128));
    defparam i3_4_lut_adj_1242.LUT_INIT = 16'h9669;
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n28731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n28730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n28729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n28728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n28727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n28726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n28725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n28724));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n28723));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n28722));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n28721));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n28720));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n28719));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n28718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n28717));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n28716));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n28715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n28714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n28713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n28712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n28711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n28710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n28709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n28708));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n28707));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n28706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n28705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n28704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n28703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n28702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n28701));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1243 (.I0(n27128), .I1(n40347), .I2(\data_out_frame[17] [1]), 
            .I3(GND_net), .O(n42528));
    defparam i2_3_lut_adj_1243.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1244 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n42235));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1244.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1245 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[5] [5]), 
            .I2(n42292), .I3(n6_adj_4357), .O(n1519));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(71[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42651));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42292));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(n40128), .I1(n27026), .I2(GND_net), 
            .I3(GND_net), .O(n40506));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(n40257), .I1(n27461), .I2(GND_net), 
            .I3(GND_net), .O(n40504));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42458));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1251 (.I0(n42680), .I1(n42856), .I2(n42292), 
            .I3(GND_net), .O(n1522));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1251.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_out_frame[12] [5]), .I1(n1519), 
            .I2(GND_net), .I3(GND_net), .O(n42344));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1253 (.I0(n27196), .I1(n26223), .I2(n40504), 
            .I3(n6_adj_4358), .O(n42613));
    defparam i4_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1254 (.I0(\data_out_frame[12] [6]), .I1(n42344), 
            .I2(\data_out_frame[14] [7]), .I3(n1522), .O(n42286));
    defparam i3_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_in_frame[5] [5]), .I1(n27347), 
            .I2(GND_net), .I3(GND_net), .O(n42258));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1256 (.I0(n42265), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n42797));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1256.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\data_in_frame[5] [7]), .I1(n42797), 
            .I2(GND_net), .I3(GND_net), .O(n42891));
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_out_frame[17] [1]), .I1(n27321), 
            .I2(GND_net), .I3(GND_net), .O(n42556));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1259 (.I0(\data_out_frame[16] [7]), .I1(n42286), 
            .I2(\data_out_frame[15] [0]), .I3(n27223), .O(n40347));
    defparam i3_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1260 (.I0(n27324), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n42807));
    defparam i2_3_lut_adj_1260.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42298));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1262 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n42727));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1262.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1263 (.I0(n42727), .I1(n42298), .I2(\data_in_frame[8] [2]), 
            .I3(n42891), .O(n10_adj_4176));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1264 (.I0(\data_out_frame[19] [2]), .I1(n40347), 
            .I2(n6_adj_4359), .I3(n42556), .O(n40598));
    defparam i1_4_lut_adj_1264.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\data_out_frame[19] [3]), .I1(n42528), 
            .I2(GND_net), .I3(GND_net), .O(n42503));
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42732));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26702));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1268 (.I0(n42732), .I1(\data_in_frame[10] [3]), 
            .I2(n42289), .I3(n25058), .O(n14_adj_4360));
    defparam i6_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(n26217), .I1(n1510), .I2(GND_net), 
            .I3(GND_net), .O(n42762));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1270 (.I0(n42850), .I1(n14_adj_4360), .I2(n10_adj_4155), 
            .I3(\data_in_frame[15] [1]), .O(n27461));
    defparam i7_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(n40578), .I1(n27461), .I2(GND_net), 
            .I3(GND_net), .O(n40502));
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1272 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42468));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1272.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[4] [7]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n42810));
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42563));
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1275 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[7] [6]), 
            .I2(n26702), .I3(\data_out_frame[9] [7]), .O(n42510));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1276 (.I0(\data_out_frame[11] [7]), .I1(n42510), 
            .I2(n27103), .I3(\data_out_frame[7] [5]), .O(n26217));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1277 (.I0(n42468), .I1(n42762), .I2(\data_out_frame[12] [2]), 
            .I3(GND_net), .O(n40033));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1277.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42711));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1279 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26939));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1280 (.I0(n26939), .I1(n42711), .I2(\data_out_frame[7] [2]), 
            .I3(GND_net), .O(n42671));   // verilog/coms.v(73[16:34])
    defparam i2_3_lut_adj_1280.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1281 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42431));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1281.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1282 (.I0(n26725), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[10] [1]), .I3(n6_adj_4361), .O(n1510));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42488));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26771));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42765));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42397));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut_4_lut (.I0(n43085), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n33940), .I3(n26622), .O(n43465));   // verilog/coms.v(127[12] 300[6])
    defparam i2_2_lut_4_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i4_4_lut_adj_1287 (.I0(n26771), .I1(n27287), .I2(n42488), 
            .I3(n6_adj_4362), .O(n1516));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n28700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n28698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n28697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n28696));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n28695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n28694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n28693));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n28692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n28691));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n28690));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n28689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n28688));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n28687));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n28686));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n28685));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n28684));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n28683));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n28682));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n28681));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n28680));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n28679));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n28678));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n28677));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n28676));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n28675));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n28674));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n28673));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n28672));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n28671));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n28670));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n28669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n28668));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n28667));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n28666));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n28665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n28664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n28663));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n28662));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n28661));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n28660));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n28659));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n28658));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n28657));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n28656));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n28655));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n28654));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n28653));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n28652));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n28651));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n28650));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n28649));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n28648));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n28647));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n28646));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n28645));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n28644));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n28643));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n28642));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n28641));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n28640));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n28639));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n28638));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n28637));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n28636));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n28635));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n28634));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n28633));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n28632));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n28631));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n28630));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n28629));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n28628));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n28627));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n28626));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n28625));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n28624));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n28623));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n28622));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n28621));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n28620));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n28619));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n28618));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n28617));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n28616));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n28615));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n28614));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42859));
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n28613));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n28612));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n28611));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n28610));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n28609));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n28608));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n28607));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n28606));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n28605));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n28604));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n28603));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n28602));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n28601));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n28600));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n28599));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n28598));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n28597));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n28596));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n28595));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n28594));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n28593));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n28592));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n28591));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n28590));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n28589));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n28588));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n28587));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n28586));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n28585));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n28584));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n28583));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n28582));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1289 (.I0(n33507), .I1(n8_adj_4363), .I2(GND_net), 
            .I3(GND_net), .O(n42216));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27287));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42572));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(n27287), .I1(\data_out_frame[5] [3]), 
            .I2(n42859), .I3(n6_adj_4364), .O(n1513));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(GND_net), .I3(GND_net), .O(n26762));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1294 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n26622), .O(n36017));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1294.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_1295 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(GND_net), .I3(GND_net), .O(n27278));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1295.LUT_INIT = 16'h6666;
    SB_LUT4 i28066_2_lut_3_lut_4_lut (.I0(n26482), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n771), .O(n42938));
    defparam i28066_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\data_out_frame[14] [4]), .I1(n27223), 
            .I2(GND_net), .I3(GND_net), .O(n26822));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_4_lut (.I0(n33940), .I1(n26622), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n44935));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i2_2_lut_adj_1297 (.I0(n42598), .I1(\data_out_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4365));
    defparam i2_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1298 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[4] [7]), 
            .I2(n42671), .I3(n26725), .O(n14_adj_4366));
    defparam i6_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1299 (.I0(n40033), .I1(n14_adj_4366), .I2(n10_adj_4365), 
            .I3(n26217), .O(n42673));
    defparam i7_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1300 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n42871));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1300.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut (.I0(n42335), .I1(n42705), .I2(\data_in_frame[11] [3]), 
            .I3(\data_in_frame[18] [0]), .O(n42865));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n42642));
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1302 (.I0(\data_out_frame[20] [3]), .I1(n39724), 
            .I2(\data_out_frame[20] [1]), .I3(n26238), .O(n42649));
    defparam i1_2_lut_3_lut_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1303 (.I0(\data_out_frame[19] [0]), .I1(n42642), 
            .I2(n42673), .I3(n1794), .O(n10_adj_4367));
    defparam i4_4_lut_adj_1303.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1304 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[13] [7]), .I3(GND_net), .O(n42915));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1304.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1305 (.I0(\data_out_frame[16] [4]), .I1(n10_adj_4367), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n42513));
    defparam i5_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1306 (.I0(n42576), .I1(n42822), .I2(n40033), 
            .I3(GND_net), .O(n40658));
    defparam i2_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(n40658), .I1(n42513), .I2(GND_net), 
            .I3(GND_net), .O(n2122));
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1308 (.I0(n33940), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n26622), .I3(GND_net), .O(n27893));
    defparam i3_3_lut_adj_1308.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(\data_out_frame[23] [5]), .I1(n42610), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4368));
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1310 (.I0(n42834), .I1(\data_out_frame[23] [4]), 
            .I2(n2122), .I3(n6_adj_4368), .O(n44563));
    defparam i4_4_lut_adj_1310.LUT_INIT = 16'h9669;
    SB_CARRY add_43_19 (.CI(n37262), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n37263));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1311 (.I0(\data_out_frame[24] [7]), .I1(n42601), 
            .I2(n42462), .I3(\data_out_frame[25] [1]), .O(n42699));
    defparam i1_2_lut_3_lut_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1312 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(n40662), .I3(n10_adj_4369), .O(n44122));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_4_lut_adj_1312.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1313 (.I0(n63_adj_4154), .I1(n63), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n63_adj_4159), .O(n42231));
    defparam i1_2_lut_4_lut_adj_1313.LUT_INIT = 16'h80ff;
    SB_LUT4 i15397_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n28456));
    defparam i15397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15398_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n28457));
    defparam i15398_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_18_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n37261), .O(n2_adj_4252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1314 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [4]), 
            .I2(n39724), .I3(n24914), .O(n39761));
    defparam i1_2_lut_3_lut_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1315 (.I0(n29941), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n5_adj_4173), .I3(n5_adj_4345), .O(n7_adj_4371));
    defparam i2_3_lut_4_lut_adj_1315.LUT_INIT = 16'hab03;
    SB_LUT4 i15399_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n28458));
    defparam i15399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_18 (.CI(n37261), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n37262));
    SB_LUT4 i15400_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n28459));
    defparam i15400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15401_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n28460));
    defparam i15401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(n33507), .I1(n8_adj_4372), .I2(GND_net), 
            .I3(GND_net), .O(n42219));
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'hdddd;
    SB_LUT4 add_43_17_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n37260), .O(n2_adj_4253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15402_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n28461));
    defparam i15402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15403_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n28462));
    defparam i15403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15404_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42225), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n28463));
    defparam i15404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_17 (.CI(n37260), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n37261));
    SB_LUT4 i15389_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n28448));
    defparam i15389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1317 (.I0(n44460), .I1(\data_out_frame[20] [6]), 
            .I2(n42513), .I3(n24914), .O(n6_adj_4301));
    defparam i1_2_lut_3_lut_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i15390_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n28449));
    defparam i15390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15391_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n28450));
    defparam i15391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15392_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n28451));
    defparam i15392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15393_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n28452));
    defparam i15393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15394_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n28453));
    defparam i15394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_16_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n37259), .O(n2_adj_4254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n37259), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n37260));
    SB_LUT4 i15395_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n28454));
    defparam i15395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n28581));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1318 (.I0(\data_in_frame[8] [7]), .I1(n27414), 
            .I2(n10), .I3(n27417), .O(n27594));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i15396_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42222), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n28455));
    defparam i15396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1319 (.I0(n40257), .I1(n42538), .I2(n40578), 
            .I3(n27461), .O(n27196));
    defparam i1_2_lut_3_lut_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_15_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n37258), .O(n2_adj_4255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 equal_132_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4373));   // verilog/coms.v(154[7:23])
    defparam equal_132_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_123_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4374));   // verilog/coms.v(154[7:23])
    defparam equal_123_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_CARRY add_43_15 (.CI(n37258), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n37259));
    SB_LUT4 add_43_14_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n37257), .O(n2_adj_4256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1320 (.I0(n42756), .I1(n40629), .I2(n42915), 
            .I3(GND_net), .O(n42693));
    defparam i2_3_lut_adj_1320.LUT_INIT = 16'h9696;
    SB_CARRY add_43_14 (.CI(n37257), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n37258));
    SB_LUT4 i1_2_lut_adj_1321 (.I0(n33507), .I1(n8_adj_4374), .I2(GND_net), 
            .I3(GND_net), .O(n42213));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'hdddd;
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n28580));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_13_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n37256), .O(n2_adj_4257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n28579));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15381_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n28440));
    defparam i15381_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_13 (.CI(n37256), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n37257));
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n28578));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_12_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n37255), .O(n2_adj_4258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1322 (.I0(r_SM_Main_2__N_3516[0]), .I1(tx_active), 
            .I2(tx_transmit_N_3413), .I3(\FRAME_MATCHER.i_31__N_2523 ), 
            .O(n2_adj_4344));
    defparam i1_2_lut_3_lut_4_lut_adj_1322.LUT_INIT = 16'hfe00;
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n28577));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1323 (.I0(n3183), .I1(n2_adj_4344), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n23831), .O(n41663));
    defparam i1_2_lut_3_lut_4_lut_adj_1323.LUT_INIT = 16'he0ee;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n28576));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1324 (.I0(\data_out_frame[5] [0]), .I1(n42331), 
            .I2(\data_out_frame[4] [6]), .I3(\data_out_frame[7] [0]), .O(n27666));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_3_lut_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1325 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n42410), .I3(n26969), .O(n27414));
    defparam i1_2_lut_3_lut_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_CARRY add_43_12 (.CI(n37255), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n37256));
    SB_LUT4 i2_3_lut_4_lut_adj_1326 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(n42353), .I3(n42727), .O(Kp_23__N_836));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1545_i8_2_lut_3_lut_4_lut (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n42410), .I3(\data_in_frame[8] [7]), .O(n8_adj_4127));
    defparam equal_1545_i8_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15382_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n28441));
    defparam i15382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15383_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n28442));
    defparam i15383_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15384_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n28443));
    defparam i15384_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n28575));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n28574));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n28573));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n28572));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n28571));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n28570));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n28569));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n28568));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n28567));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n28566));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n28565));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n28564));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n28563));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n28562));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n28561));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n28560));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n28559));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n28558));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n28557));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n28556));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n28555));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n28554));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n28553));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n28552));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n28551));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n28550));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n28549));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n28548));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n28547));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n28546));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n28545));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n28544));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n28543));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n28542));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(CLK_c), 
           .D(n28541));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18]_c [1]), .C(CLK_c), 
           .D(n28540));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(CLK_c), 
           .D(n28539));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n28538));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n28537));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n28536));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18][6] ), .C(CLK_c), 
           .D(n28535));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n28534));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n28533));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n28532));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n28531));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n28530));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n28529));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n28528));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n28527));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n28526));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(CLK_c), 
           .D(n28525));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(CLK_c), 
           .D(n28524));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n28523));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n28522));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(CLK_c), 
           .D(n28521));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n28520));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n28519));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n28518));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n28517));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n28516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n28515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n28514));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n28513));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n28296));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15385_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n28444));
    defparam i15385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n28512));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n28511));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n28510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n28509));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n28508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n28507));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15386_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n28445));
    defparam i15386_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n28164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n28506));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n28505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n28504));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n28503));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n28502));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n28501));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n28500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n28499));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15387_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n28446));
    defparam i15387_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15388_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42213), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n28447));
    defparam i15388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n28498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n28497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n28496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n28495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n28494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n28493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n28492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n28491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n28490));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n28489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n28488));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n28487));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n28486));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n28485));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n28484));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n28483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n28482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n28481));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n28480));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n28479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n28478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n28477));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n28476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n28475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n28474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n28473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n28472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n28471));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n28470));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n28469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n28468));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n28467));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n28466));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n28465));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n28464));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n28463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n28462));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15373_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n28432));
    defparam i15373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15374_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n28433));
    defparam i15374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1327 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n42410), .I3(n42269), .O(Kp_23__N_1210));
    defparam i1_2_lut_3_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1328 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[5] [6]), .O(n27660));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1329 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(n42413), .I3(\data_in_frame[8] [4]), .O(n27381));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1330 (.I0(n26870), .I1(n42400), .I2(\data_in_frame[0] [0]), 
            .I3(Kp_23__N_990), .O(n42413));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i15375_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n28434));
    defparam i15375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n28461));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n28460));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15376_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n28435));
    defparam i15376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n28459));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n28458));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n28457));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n28456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n28455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n28454));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n28453));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1331 (.I0(n27066), .I1(\data_in_frame[5] [5]), 
            .I2(n27347), .I3(\data_in_frame[7] [7]), .O(n42265));
    defparam i1_2_lut_3_lut_4_lut_adj_1331.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n28452));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n28451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n28450));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15377_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n28436));
    defparam i15377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15378_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n28437));
    defparam i15378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15379_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n28438));
    defparam i15379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_2_lut_4_lut (.I0(\data_in_frame[10] [5]), .I1(n10_adj_4162), 
            .I2(\data_in_frame[17] [5]), .I3(n42696), .O(n17_adj_4280));
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15380_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42219), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n28439));
    defparam i15380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n28449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n28448));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1332 (.I0(\data_in_frame[10] [5]), .I1(n10_adj_4162), 
            .I2(\data_in_frame[17] [5]), .I3(n40662), .O(n40652));
    defparam i1_2_lut_4_lut_adj_1332.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n28447));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n28446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n28445));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n28444));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n28443));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n28442));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n28441));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n28440));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n28439));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33677_3_lut_4_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[4]), 
            .I2(n81), .I3(n359), .O(tx_transmit_N_3413));   // verilog/coms.v(214[11:56])
    defparam i33677_3_lut_4_lut.LUT_INIT = 16'h070f;
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n28438));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n28437));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n28436));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n28435));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n28434));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n28433));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1333 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[2] [1]), .O(n42400));
    defparam i2_3_lut_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n28432));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1334 (.I0(n27278), .I1(n26762), .I2(\data_out_frame[14] [4]), 
            .I3(GND_net), .O(n27321));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1334.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n28431));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n28430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n28429));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1335 (.I0(\FRAME_MATCHER.state [3]), .I1(n23831), 
            .I2(n3183), .I3(n1_adj_4309), .O(n41665));
    defparam i1_3_lut_4_lut_adj_1335.LUT_INIT = 16'haa80;
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n28428));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1336 (.I0(n33507), .I1(n8_adj_4373), .I2(GND_net), 
            .I3(GND_net), .O(n42222));
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'hdddd;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n28427));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n28426));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n28425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n28424));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n28423));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n28422));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n28421));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n28420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n28419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n28418));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n28417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n28416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n28415));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n28414));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n28413));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n28410));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n28409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n28408));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n28407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n28406));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n28405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n28403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n28402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n28401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n28400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n28399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n28398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n28397));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1337 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(n40128), .I3(n27026), .O(n42756));
    defparam i1_2_lut_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n28396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n28395));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(n27278), .I1(n26762), .I2(n26822), 
            .I3(GND_net), .O(n1794));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n28394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n28393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n28392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n28391));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n28390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n28389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n28388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n28387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n28386));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n28385));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n28384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n28383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n28382));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n28381));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n28380));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n28379));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15365_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n28424));
    defparam i15365_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n28378));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n28377));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n28376));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n28375));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n28374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n28373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n28372));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n28371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n28370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n28369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n28368));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n28367));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n28366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n28365));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n28364));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n28363));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1339 (.I0(\data_out_frame[19] [3]), .I1(n42528), 
            .I2(\data_out_frame[25] [6]), .I3(n40598), .O(n42834));
    defparam i2_3_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n28362));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15366_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n28425));
    defparam i15366_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n28361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n28360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n28359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n28358));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1340 (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[11] [7]), .I3(\data_out_frame[12] [0]), 
            .O(n42598));
    defparam i1_2_lut_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n28357));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15367_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n28426));
    defparam i15367_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n28356));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1341 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n42909));
    defparam i1_2_lut_3_lut_adj_1341.LUT_INIT = 16'h9696;
    SB_LUT4 i15368_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n28427));
    defparam i15368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n28355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n28354));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1342 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[6] [1]), .O(n6_adj_4362));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n28353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n28352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n28351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n28350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n28349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n28348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n28347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n28346));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n28345));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n28344));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n28343));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n28342));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n26725));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n28341));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15369_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n28428));
    defparam i15369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1344 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(n42810), .I3(\data_out_frame[5] [1]), .O(n27103));
    defparam i2_3_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n28340));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n28339));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_4_lut (.I0(n27324), .I1(\data_out_frame[17] [0]), .I2(\data_out_frame[16] [7]), 
            .I3(\data_out_frame[16] [6]), .O(n6_adj_4359));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n28338));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n28337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n28336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n28335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n28334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n28333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n28332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n28331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n28330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n28329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n28328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n28327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n28326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n28325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n28324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n28323));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n28322));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1345 (.I0(\data_in_frame[8] [7]), .I1(n27414), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1221));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n28321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n28320));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15370_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n28429));
    defparam i15370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n28319));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n28318));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n28317));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n28316));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n28315));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15371_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n28430));
    defparam i15371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n28314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n28313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n28312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n28311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n28310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n28309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n28308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n28307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n28306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n28305));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15372_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42216), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n28431));
    defparam i15372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1346 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(Kp_23__N_869), .I3(GND_net), .O(n43987));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_11_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n37254), .O(n2_adj_4259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i9_4_lut_adj_1347 (.I0(n43987), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[1] [1]), .O(n26_adj_4375));
    defparam i9_4_lut_adj_1347.LUT_INIT = 16'h4010;
    SB_LUT4 i13_4_lut_adj_1348 (.I0(n27340), .I1(n26_adj_4375), .I2(\data_in_frame[0] [6]), 
            .I3(n42416), .O(n30_adj_4376));
    defparam i13_4_lut_adj_1348.LUT_INIT = 16'h4004;
    SB_LUT4 i6_4_lut_adj_1349 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_869), 
            .I2(n42252), .I3(n42367), .O(n23_adj_4377));
    defparam i6_4_lut_adj_1349.LUT_INIT = 16'h1248;
    SB_LUT4 i1_2_lut_4_lut_adj_1350 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[4] [1]), .I3(n42862), .O(n6_adj_4357));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i31547_2_lut (.I0(n27360), .I1(n26838), .I2(GND_net), .I3(GND_net), 
            .O(n46425));
    defparam i31547_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1351 (.I0(n23_adj_4377), .I1(n30_adj_4376), .I2(n24130), 
            .I3(n26774), .O(n32));
    defparam i15_4_lut_adj_1351.LUT_INIT = 16'h0008;
    SB_LUT4 i4_4_lut_adj_1352 (.I0(n42696), .I1(Kp_23__N_1466), .I2(n40235), 
            .I3(n42865), .O(n10_adj_4369));
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1353 (.I0(n2_adj_4341), .I1(n4_adj_4342), 
            .I2(n23831), .I3(n3183), .O(n5_adj_4378));
    defparam i1_2_lut_3_lut_4_lut_adj_1353.LUT_INIT = 16'hfeee;
    SB_CARRY add_43_11 (.CI(n37254), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n37255));
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n42862));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n28304));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i10_4_lut_adj_1355 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[1] [2]), .O(n27_adj_4379));
    defparam i10_4_lut_adj_1355.LUT_INIT = 16'h8000;
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n28303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n28302));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16_4_lut_adj_1356 (.I0(n27_adj_4379), .I1(n32), .I2(n46425), 
            .I3(n22_adj_4380), .O(\FRAME_MATCHER.state_31__N_2624 [3]));
    defparam i16_4_lut_adj_1356.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[6] [0]), 
            .I2(n42909), .I3(GND_net), .O(n6_adj_4364));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1358 (.I0(\data_out_frame[12] [4]), .I1(n1516), 
            .I2(\data_out_frame[14] [6]), .I3(n42344), .O(n27324));
    defparam i2_3_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1359 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[6] [5]), .O(n42874));
    defparam i1_2_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[4]), 
            .I2(n26646), .I3(GND_net), .O(n59));   // verilog/coms.v(214[11:56])
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'hf8f8;
    SB_LUT4 equal_125_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4381));   // verilog/coms.v(154[7:23])
    defparam equal_125_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 add_43_10_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n37253), .O(n2_adj_4261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1361 (.I0(n33507), .I1(n8_adj_4381), .I2(GND_net), 
            .I3(GND_net), .O(n42225));
    defparam i1_2_lut_adj_1361.LUT_INIT = 16'hdddd;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[15] [5]), .I3(n42556), .O(n26_adj_4334));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1362 (.I0(\data_out_frame[12] [4]), .I1(n1516), 
            .I2(\data_out_frame[14] [5]), .I3(n26762), .O(n27223));
    defparam i2_3_lut_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1363 (.I0(\FRAME_MATCHER.state [2]), .I1(n7_adj_4343), 
            .I2(n36017), .I3(\FRAME_MATCHER.state_31__N_2624 [3]), .O(n41733));
    defparam i1_4_lut_adj_1363.LUT_INIT = 16'hcdcc;
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n28301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n28300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n28299));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1364 (.I0(\data_out_frame[5] [6]), .I1(n27287), 
            .I2(\data_out_frame[10] [0]), .I3(\data_out_frame[5] [2]), .O(n6_adj_4361));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1365 (.I0(Kp_23__N_1221), .I1(n42871), .I2(\data_in_frame[16] [0]), 
            .I3(n42693), .O(n12_adj_4382));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1366 (.I0(\data_in_frame[9] [1]), .I1(n12_adj_4382), 
            .I2(\data_in_frame[18] [2]), .I3(n42705), .O(n42825));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42295));
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h6666;
    SB_LUT4 i5_2_lut_4_lut_adj_1368 (.I0(\data_out_frame[5] [6]), .I1(n27287), 
            .I2(\data_out_frame[10] [0]), .I3(n42364), .O(n16_adj_4312));   // verilog/coms.v(74[16:27])
    defparam i5_2_lut_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1369 (.I0(\FRAME_MATCHER.state [4]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41669));
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1370 (.I0(\FRAME_MATCHER.state [5]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41805));
    defparam i1_2_lut_adj_1370.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1371 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [2]), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[11] [4]), 
            .O(n42853));
    defparam i2_3_lut_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1372 (.I0(\FRAME_MATCHER.state [6]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41737));
    defparam i1_2_lut_adj_1372.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1373 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[4] [2]), .O(n27705));
    defparam i1_2_lut_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n28298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n28297));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15357_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n28416));
    defparam i15357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15358_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n28417));
    defparam i15358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1374 (.I0(\FRAME_MATCHER.state [7]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41739));
    defparam i1_2_lut_adj_1374.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1375 (.I0(n42338), .I1(\data_out_frame[8] [7]), 
            .I2(n27666), .I3(\data_out_frame[11] [3]), .O(n42708));
    defparam i2_3_lut_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i15359_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n28418));
    defparam i15359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15360_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n28419));
    defparam i15360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_10 (.CI(n37253), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n37254));
    SB_LUT4 equal_126_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4160));   // verilog/coms.v(154[7:23])
    defparam equal_126_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15361_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n28420));
    defparam i15361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1376 (.I0(\FRAME_MATCHER.state [8]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41803));
    defparam i1_2_lut_adj_1376.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_9_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n37252), .O(n2_adj_4263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1377 (.I0(\FRAME_MATCHER.state [9]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41801));
    defparam i1_2_lut_adj_1377.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1378 (.I0(\data_out_frame[13] [4]), .I1(n40283), 
            .I2(n27554), .I3(n27679), .O(n40517));
    defparam i2_3_lut_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(n40652), .I1(n40578), .I2(\data_in_frame[19] [6]), 
            .I3(GND_net), .O(n39733));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_CARRY add_43_9 (.CI(n37252), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n37253));
    SB_LUT4 i15362_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n28421));
    defparam i15362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_8_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n37251), .O(n2_adj_4265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(\data_in_frame[1] [0]), .I1(n42407), 
            .I2(GND_net), .I3(GND_net), .O(n26903));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1381 (.I0(\FRAME_MATCHER.state [10]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41741));
    defparam i1_2_lut_adj_1381.LUT_INIT = 16'h8888;
    SB_CARRY add_43_8 (.CI(n37251), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n37252));
    SB_LUT4 add_43_7_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n37250), .O(n2_adj_4267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1382 (.I0(\FRAME_MATCHER.state [11]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41799));
    defparam i1_2_lut_adj_1382.LUT_INIT = 16'h8888;
    SB_LUT4 i15363_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n28422));
    defparam i15363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1383 (.I0(n42338), .I1(n42718), .I2(\data_out_frame[11] [3]), 
            .I3(\data_out_frame[11] [4]), .O(n10_adj_4319));
    defparam i2_2_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n26861));
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1385 (.I0(n40542), .I1(n40604), .I2(n42544), 
            .I3(GND_net), .O(n10_adj_4315));
    defparam i2_2_lut_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(\FRAME_MATCHER.state [12]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41797));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h8888;
    SB_LUT4 i15364_3_lut_4_lut (.I0(n10_adj_4370), .I1(n42203), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n28423));
    defparam i15364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_7 (.CI(n37250), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n37251));
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[12] [0]), .I3(GND_net), .O(n27498));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[10] [5]), .I3(\data_out_frame[8] [4]), .O(n9_adj_4323));   // verilog/coms.v(71[16:27])
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[15] [5]), .I3(GND_net), .O(n42780));
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1389 (.I0(n26870), .I1(n42400), .I2(\data_in_frame[0] [0]), 
            .I3(GND_net), .O(Kp_23__N_993));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1390 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[4] [7]), 
            .I2(n42671), .I3(\data_out_frame[13] [7]), .O(n42847));
    defparam i1_2_lut_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1391 (.I0(\FRAME_MATCHER.state [13]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41795));
    defparam i1_2_lut_adj_1391.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1392 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[14] [1]), .I3(GND_net), .O(n10_adj_4304));
    defparam i1_2_lut_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_6_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n37249), .O(n2_adj_4269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(\FRAME_MATCHER.state [14]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41743));
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [6]), 
            .I2(n43813), .I3(GND_net), .O(n39642));
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'h6969;
    SB_LUT4 i3_3_lut_4_lut (.I0(n27066), .I1(n42258), .I2(n42443), .I3(\data_in_frame[10] [2]), 
            .O(n11));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34337 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n49287));
    defparam byte_transmit_counter_0__bdd_4_lut_34337.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(\FRAME_MATCHER.state [15]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41793));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h8888;
    SB_CARRY add_43_6 (.CI(n37249), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n37250));
    SB_LUT4 add_43_5_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n37248), .O(n2_adj_4271)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1396 (.I0(n42563), .I1(n42810), .I2(\data_out_frame[5] [1]), 
            .I3(n42847), .O(n6_adj_4303));
    defparam i1_2_lut_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1397 (.I0(\FRAME_MATCHER.state [16]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41791));
    defparam i1_2_lut_adj_1397.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1398 (.I0(n40052), .I1(n42462), .I2(\data_out_frame[25] [1]), 
            .I3(n42886), .O(n6_adj_4299));
    defparam i1_2_lut_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1399 (.I0(n27041), .I1(n42538), .I2(n40578), 
            .I3(n40652), .O(n6_adj_4358));
    defparam i1_2_lut_3_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(n27041), .I1(n42538), .I2(\data_in_frame[19] [2]), 
            .I3(GND_net), .O(n42768));
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1401 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n42277));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1401.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(\FRAME_MATCHER.state [17]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41789));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h8888;
    SB_CARRY add_43_5 (.CI(n37248), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n37249));
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n27340));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1404 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [5]), 
            .I2(n26771), .I3(n1191), .O(n42680));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1405 (.I0(\FRAME_MATCHER.state [18]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41787));
    defparam i1_2_lut_adj_1405.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1406 (.I0(\data_in_frame[0] [4]), .I1(n42255), 
            .I2(\data_in_frame[2] [1]), .I3(Kp_23__N_869), .O(n22_adj_4380));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_4_lut_adj_1406.LUT_INIT = 16'h0990;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(\FRAME_MATCHER.state [19]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41785));
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1408 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26942));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1408.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1409 (.I0(\data_out_frame[25] [0]), .I1(\data_out_frame[20] [3]), 
            .I2(n39724), .I3(n42312), .O(n42840));
    defparam i1_2_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1410 (.I0(n26235), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[15] [4]), .I3(\data_out_frame[15] [5]), 
            .O(n4));
    defparam i1_2_lut_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1411 (.I0(\data_in_frame[13] [2]), .I1(n42900), 
            .I2(\data_in_frame[10] [6]), .I3(\data_in_frame[10] [7]), .O(n42619));
    defparam i3_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1412 (.I0(\data_in_frame[0] [4]), .I1(n42255), 
            .I2(n42750), .I3(n10_adj_4354), .O(n40128));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1413 (.I0(\data_in_frame[0] [4]), .I1(n42255), 
            .I2(\data_in_frame[5] [2]), .I3(n42744), .O(n27026));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1414 (.I0(n63_adj_4154), .I1(n63), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n92[1]));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_adj_1414.LUT_INIT = 16'h8080;
    SB_LUT4 add_43_4_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n37247), .O(n2_adj_4273)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(n63_adj_4154), .I1(n63), .I2(n63_adj_4159), 
            .I3(GND_net), .O(n23831));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'h8080;
    SB_LUT4 i15347_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n28406));
    defparam i15347_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_3_lut_adj_1416 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [7]), 
            .I2(n42662), .I3(GND_net), .O(n8_adj_4384));
    defparam i3_3_lut_adj_1416.LUT_INIT = 16'h9696;
    SB_LUT4 i15348_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n28407));
    defparam i15348_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15349_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n28408));
    defparam i15349_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n49287_bdd_4_lut (.I0(n49287), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n49290));
    defparam n49287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15350_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n28409));
    defparam i15350_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15351_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n28410));
    defparam i15351_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15354_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n28413));
    defparam i15354_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1417 (.I0(n40128), .I1(n27417), .I2(\data_in_frame[9] [4]), 
            .I3(GND_net), .O(n40629));
    defparam i1_2_lut_3_lut_adj_1417.LUT_INIT = 16'h9696;
    SB_LUT4 i15355_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n28414));
    defparam i15355_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15356_3_lut_4_lut (.I0(n10_adj_4370), .I1(n43891), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n28415));
    defparam i15356_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(n40128), .I1(n27417), .I2(n42434), 
            .I3(GND_net), .O(n8_adj_4195));
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1419 (.I0(\data_in_frame[15] [4]), .I1(n27381), 
            .I2(n8_adj_4384), .I3(n42619), .O(n40662));
    defparam i1_4_lut_adj_1419.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1420 (.I0(n40114), .I1(\data_out_frame[20] [1]), 
            .I2(n42645), .I3(\data_out_frame[20] [5]), .O(n42551));
    defparam i1_2_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1421 (.I0(\FRAME_MATCHER.state [20]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41783));
    defparam i1_2_lut_adj_1421.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1422 (.I0(\data_out_frame[5] [0]), .I1(n42331), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[4] [5]), .O(n27492));   // verilog/coms.v(71[16:62])
    defparam i1_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(n2122), .I1(n42588), .I2(\data_out_frame[25] [4]), 
            .I3(GND_net), .O(n42831));
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1424 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(n42801), .O(n6_adj_4281));
    defparam i1_2_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\FRAME_MATCHER.state [21]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41781));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1426 (.I0(n2122), .I1(n42588), .I2(n40073), 
            .I3(\data_out_frame[25] [5]), .O(n42610));
    defparam i2_3_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i20466_2_lut_3_lut (.I0(n2482), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n33507));
    defparam i20466_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_adj_1427 (.I0(\FRAME_MATCHER.state [22]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41779));
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1428 (.I0(n3183), .I1(n2_adj_4344), .I2(n42940), 
            .I3(n42231), .O(n39_adj_4385));
    defparam i1_3_lut_4_lut_adj_1428.LUT_INIT = 16'hef00;
    SB_LUT4 i1_2_lut_4_lut_adj_1429 (.I0(\data_out_frame[20] [3]), .I1(n39724), 
            .I2(n42312), .I3(n39761), .O(n39689));
    defparam i1_2_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1430 (.I0(\FRAME_MATCHER.state [23]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41777));
    defparam i1_2_lut_adj_1430.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1431 (.I0(n26482), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n85));
    defparam i1_2_lut_3_lut_adj_1431.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(\FRAME_MATCHER.state [24]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41725));
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1433 (.I0(n26238), .I1(n40114), .I2(n42645), 
            .I3(\data_out_frame[20] [5]), .O(n42616));
    defparam i2_3_lut_4_lut_adj_1433.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(\FRAME_MATCHER.state [25]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41729));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(n27210), .I1(n42465), .I2(n43940), 
            .I3(\data_out_frame[19] [5]), .O(n39632));
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(\FRAME_MATCHER.state [26]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41775));
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1437 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[16] [1]), .I3(\data_in_frame[14] [1]), .O(n30));
    defparam i1_2_lut_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1438 (.I0(\FRAME_MATCHER.state [27]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41773));
    defparam i1_2_lut_adj_1438.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1439 (.I0(n42367), .I1(n42724), .I2(\data_in_frame[4] [5]), 
            .I3(n27337), .O(n42410));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1440 (.I0(n26238), .I1(n42646), .I2(\data_out_frame[20] [5]), 
            .I3(\data_out_frame[25] [7]), .O(n10_adj_4220));
    defparam i2_2_lut_4_lut_adj_1440.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1441 (.I0(\FRAME_MATCHER.state [28]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41771));
    defparam i1_2_lut_adj_1441.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1442 (.I0(\data_in_frame[19] [1]), .I1(n26223), 
            .I2(n42768), .I3(\data_in_frame[21] [3]), .O(n43504));
    defparam i2_3_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1443 (.I0(\FRAME_MATCHER.state [29]), .I1(n4_adj_4342), 
            .I2(n2_adj_4341), .I3(n1_adj_4386), .O(n8_adj_4208));
    defparam i1_4_lut_adj_1443.LUT_INIT = 16'haaa8;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(n42367), .I1(n42724), .I2(\data_in_frame[6] [5]), 
            .I3(n42388), .O(Kp_23__N_1095));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_in_frame[11] [4]), .I1(n42385), .I2(\data_in_frame[16] [1]), 
            .I3(GND_net), .O(n16_adj_4199));
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15330_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n28389));
    defparam i15330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15331_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n28390));
    defparam i15331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15332_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n28391));
    defparam i15332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15333_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n28392));
    defparam i15333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1445 (.I0(n26969), .I1(n10), .I2(\data_in_frame[9] [2]), 
            .I3(n42693), .O(n6_adj_4192));
    defparam i1_2_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 i15334_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n28393));
    defparam i15334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15335_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n28394));
    defparam i15335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15336_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n28395));
    defparam i15336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15337_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42225), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n28396));
    defparam i15337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1446 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[9] [0]), .I3(GND_net), .O(n27547));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1446.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1447 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[6] [6]), .I3(\data_out_frame[9] [2]), .O(n42238));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1448 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[4] [7]), 
            .I2(n42671), .I3(GND_net), .O(n27121));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1448.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1449 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[4] [7]), 
            .I2(n10_adj_4325), .I3(n42338), .O(n42877));   // verilog/coms.v(73[16:34])
    defparam i5_3_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1450 (.I0(\data_out_frame[11] [4]), .I1(n27666), 
            .I2(n42238), .I3(n27492), .O(n12_adj_4306));
    defparam i3_3_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_out_frame[11] [4]), .I1(n27666), 
            .I2(n42238), .I3(GND_net), .O(n6_adj_4321));
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 i15322_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n28381));
    defparam i15322_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1452 (.I0(\data_in_frame[9] [3]), .I1(n10), 
            .I2(n27417), .I3(GND_net), .O(n27438));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i15323_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n28382));
    defparam i15323_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15324_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n28383));
    defparam i15324_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15325_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n28384));
    defparam i15325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1453 (.I0(n1475), .I1(tx_transmit_N_3413), 
            .I2(n23831), .I3(\FRAME_MATCHER.i_31__N_2523 ), .O(n1_adj_4308));
    defparam i1_3_lut_4_lut_adj_1453.LUT_INIT = 16'he000;
    SB_LUT4 i15326_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n28385));
    defparam i15326_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15327_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n28386));
    defparam i15327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15328_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n28387));
    defparam i15328_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15329_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42222), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n28388));
    defparam i15329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15314_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n28373));
    defparam i15314_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1454 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n33507), .O(n43891));
    defparam i2_3_lut_4_lut_adj_1454.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1455 (.I0(\FRAME_MATCHER.state [30]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41769));
    defparam i1_2_lut_adj_1455.LUT_INIT = 16'h8888;
    SB_LUT4 i15315_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n28374));
    defparam i15315_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15316_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n28375));
    defparam i15316_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1456 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n33507), .O(n42203));
    defparam i2_3_lut_4_lut_adj_1456.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n26622), .I3(GND_net), .O(n26617));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'hfefe;
    SB_LUT4 i15317_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n28376));
    defparam i15317_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_3_lut_4_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[5] [7]), .O(n42856));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15318_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n28377));
    defparam i15318_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15319_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n28378));
    defparam i15319_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15320_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n28379));
    defparam i15320_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15321_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42213), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n28380));
    defparam i15321_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2149_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4144));
    defparam i2149_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i15306_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n28365));
    defparam i15306_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1458 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [6]), 
            .I2(n42633), .I3(n39699), .O(n27041));
    defparam i2_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1459 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n6014));
    defparam i1_2_lut_3_lut_adj_1459.LUT_INIT = 16'h0202;
    SB_LUT4 i2_2_lut_3_lut_adj_1460 (.I0(\data_in_frame[12] [1]), .I1(n40128), 
            .I2(\data_in_frame[12] [2]), .I3(GND_net), .O(n10_adj_4185));
    defparam i2_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i15307_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n28366));
    defparam i15307_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15308_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n28367));
    defparam i15308_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1461 (.I0(n40257), .I1(n42538), .I2(\data_in_frame[19] [3]), 
            .I3(GND_net), .O(n42525));
    defparam i1_2_lut_3_lut_adj_1461.LUT_INIT = 16'h9696;
    SB_LUT4 i15309_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n28368));
    defparam i15309_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1462 (.I0(\data_in_frame[16] [6]), .I1(n42906), 
            .I2(n42844), .I3(n39699), .O(n43998));
    defparam i2_3_lut_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1463 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [3]), .O(n27347));
    defparam i2_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i17076_3_lut (.I0(\data_out_frame[18]_c [1]), .I1(\displacement[17] ), 
            .I2(n23943), .I3(GND_net), .O(n28540));
    defparam i17076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15310_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n28369));
    defparam i15310_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15311_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n28370));
    defparam i15311_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15312_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n28371));
    defparam i15312_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15313_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42219), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n28372));
    defparam i15313_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1464 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n87), .I3(n1), .O(n27762));   // verilog/coms.v(112[11:16])
    defparam i3_3_lut_4_lut_adj_1464.LUT_INIT = 16'h0004;
    SB_LUT4 i3_4_lut_3_lut (.I0(n42777), .I1(n39642), .I2(n2063), .I3(GND_net), 
            .O(n42601));
    defparam i3_4_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1465 (.I0(n44460), .I1(n42777), .I2(n42831), 
            .I3(\data_out_frame[23] [2]), .O(n42486));
    defparam i2_3_lut_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i15298_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n28357));
    defparam i15298_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15299_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n28358));
    defparam i15299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15300_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n28359));
    defparam i15300_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15301_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n28360));
    defparam i15301_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1466 (.I0(\data_in_frame[2] [3]), .I1(n42246), 
            .I2(n26838), .I3(\data_in_frame[4] [5]), .O(n42404));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i15302_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n28361));
    defparam i15302_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1467 (.I0(n31), .I1(n24130), .I2(n26617), 
            .I3(n78), .O(n27753));
    defparam i2_3_lut_4_lut_adj_1467.LUT_INIT = 16'h0100;
    SB_LUT4 i15303_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n28362));
    defparam i15303_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1468 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n26622), .O(n5_adj_4173));
    defparam i2_3_lut_4_lut_adj_1468.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1469 (.I0(\data_in_frame[10] [4]), .I1(n26999), 
            .I2(n27061), .I3(GND_net), .O(n42657));
    defparam i1_2_lut_3_lut_adj_1469.LUT_INIT = 16'h9696;
    SB_LUT4 i15304_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n28363));
    defparam i15304_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15305_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42216), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n28364));
    defparam i15305_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1362_2_lut_3_lut (.I0(n31), .I1(n24130), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n5785));
    defparam i1362_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i6_2_lut_3_lut (.I0(n6_adj_4300), .I1(n42673), .I2(\data_out_frame[15] [5]), 
            .I3(GND_net), .O(n20_adj_4296));
    defparam i6_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1470 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(n42407), .I3(\data_in_frame[3] [0]), .O(n27534));
    defparam i2_3_lut_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1471 (.I0(n6_adj_4300), .I1(n42673), .I2(n42494), 
            .I3(n40582), .O(n44460));
    defparam i2_3_lut_4_lut_adj_1471.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1472 (.I0(\data_in_frame[7] [6]), .I1(n42391), 
            .I2(n27026), .I3(GND_net), .O(n42434));
    defparam i1_2_lut_3_lut_adj_1472.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1473 (.I0(\data_in_frame[7] [6]), .I1(n42391), 
            .I2(n10_adj_4177), .I3(Kp_23__N_1233), .O(n27639));
    defparam i5_3_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1474 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n44_adj_4229));   // verilog/coms.v(231[5:23])
    defparam i16_4_lut_adj_1474.LUT_INIT = 16'hfffe;
    SB_LUT4 i15290_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n28349));
    defparam i15290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_3_lut_4_lut (.I0(\data_in_frame[7] [6]), .I1(n42391), .I2(n27026), 
            .I3(n23), .O(n28));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'hff9f;
    SB_LUT4 i1_2_lut_3_lut_adj_1475 (.I0(n27066), .I1(\data_in_frame[6] [1]), 
            .I2(Kp_23__N_836), .I3(GND_net), .O(n6_adj_4171));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1475.LUT_INIT = 16'h9696;
    SB_LUT4 i15291_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n28350));
    defparam i15291_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15292_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n28351));
    defparam i15292_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15293_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n28352));
    defparam i15293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1476 (.I0(n33507), .I1(n8_adj_4160), .I2(n10_adj_4387), 
            .I3(GND_net), .O(n42230));
    defparam i1_2_lut_3_lut_adj_1476.LUT_INIT = 16'hfdfd;
    SB_LUT4 i15294_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n28353));
    defparam i15294_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1477 (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4154), 
            .I2(n63), .I3(GND_net), .O(n29941));   // verilog/coms.v(112[11:16])
    defparam i1_3_lut_adj_1477.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_456_Select_2_i5_4_lut (.I0(n63_adj_4159), .I1(\FRAME_MATCHER.i_31__N_2524 ), 
            .I2(n3303), .I3(n29941), .O(n5_adj_4388));
    defparam select_456_Select_2_i5_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i15295_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n28354));
    defparam i15295_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15296_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n28355));
    defparam i15296_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1478 (.I0(n5_adj_4388), .I1(n63_adj_4159), .I2(n3183), 
            .I3(n29941), .O(n6_adj_4389));
    defparam i1_4_lut_adj_1478.LUT_INIT = 16'heaaa;
    SB_LUT4 i20543_3_lut (.I0(n63_adj_4159), .I1(n4452), .I2(n29941), 
            .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2720 [2]));   // verilog/coms.v(259[6] 261[9])
    defparam i20543_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_2_lut_3_lut_adj_1479 (.I0(n33507), .I1(n8_adj_4160), .I2(n10_adj_4370), 
            .I3(GND_net), .O(n42229));
    defparam i1_2_lut_3_lut_adj_1479.LUT_INIT = 16'hfdfd;
    SB_LUT4 i4_4_lut_adj_1480 (.I0(n7_adj_4371), .I1(\FRAME_MATCHER.state_31__N_2720 [2]), 
            .I2(n6_adj_4389), .I3(n52), .O(n49530));
    defparam i4_4_lut_adj_1480.LUT_INIT = 16'hfafe;
    SB_LUT4 i15297_3_lut_4_lut (.I0(n10_adj_4387), .I1(n42203), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n28356));
    defparam i15297_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_135_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4387));   // verilog/coms.v(154[7:23])
    defparam equal_135_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [4]), 
            .I2(\data_out_frame[20] [2]), .I3(n2206), .O(n42645));
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1482 (.I0(n40052), .I1(n42462), .I2(n42840), 
            .I3(n42627), .O(n42903));
    defparam i2_3_lut_4_lut_adj_1482.LUT_INIT = 16'h9669;
    SB_LUT4 i15282_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n28341));
    defparam i15282_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15283_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n28342));
    defparam i15283_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15284_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n28343));
    defparam i15284_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i33750_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n27998));
    defparam i33750_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 equal_143_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4370));   // verilog/coms.v(154[7:23])
    defparam equal_143_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1483 (.I0(n36013), .I1(\FRAME_MATCHER.i_31__N_2524 ), 
            .I2(n3303), .I3(n42231), .O(n5_adj_4390));
    defparam i1_4_lut_adj_1483.LUT_INIT = 16'heeea;
    SB_LUT4 i3_4_lut_adj_1484 (.I0(n5_adj_4390), .I1(n39_adj_4385), .I2(n85), 
            .I3(n27_adj_4348), .O(n49529));
    defparam i3_4_lut_adj_1484.LUT_INIT = 16'hefee;
    SB_LUT4 i15285_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n28344));
    defparam i15285_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15286_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n28345));
    defparam i15286_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15287_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n28346));
    defparam i15287_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15288_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n28347));
    defparam i15288_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15289_3_lut_4_lut (.I0(n10_adj_4387), .I1(n43891), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n28348));
    defparam i15289_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15238_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n28297));
    defparam i15238_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15239_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n28298));
    defparam i15239_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15240_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n28299));
    defparam i15240_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15241_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n28300));
    defparam i15241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15237_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n28296));
    defparam i15237_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15234_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n28293));
    defparam i15234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15235_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n28294));
    defparam i15235_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15236_3_lut_4_lut (.I0(n8_adj_4363), .I1(n42206), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n28295));
    defparam i15236_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1485 (.I0(\data_out_frame[20] [3]), .I1(n39724), 
            .I2(\data_out_frame[24] [0]), .I3(\data_out_frame[23] [5]), 
            .O(n42771));
    defparam i2_3_lut_4_lut_adj_1485.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1486 (.I0(n26235), .I1(\data_out_frame[17] [6]), 
            .I2(n42783), .I3(GND_net), .O(n6_adj_4292));
    defparam i1_2_lut_3_lut_adj_1486.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1487 (.I0(n26235), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n10_adj_4276));
    defparam i2_2_lut_3_lut_adj_1487.LUT_INIT = 16'h9696;
    SB_LUT4 i15274_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n28333));
    defparam i15274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15275_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n28334));
    defparam i15275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15276_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n28335));
    defparam i15276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15277_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n28336));
    defparam i15277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15278_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n28337));
    defparam i15278_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15279_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n28338));
    defparam i15279_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15280_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n28339));
    defparam i15280_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15281_3_lut_4_lut (.I0(n8_adj_4160), .I1(n42206), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n28340));
    defparam i15281_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_137_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4363));   // verilog/coms.v(154[7:23])
    defparam equal_137_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_138_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4372));   // verilog/coms.v(154[7:23])
    defparam equal_138_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_adj_1488 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[5] [7]), .I3(n42797), .O(n6_adj_4163));
    defparam i1_2_lut_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i15266_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n28325));
    defparam i15266_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15267_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n28326));
    defparam i15267_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15268_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n28327));
    defparam i15268_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15269_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n28328));
    defparam i15269_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1489 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n42449));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1489.LUT_INIT = 16'h9696;
    SB_LUT4 i15270_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n28329));
    defparam i15270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15271_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n28330));
    defparam i15271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15272_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n28331));
    defparam i15272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15273_3_lut_4_lut (.I0(n8_adj_4381), .I1(n42206), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n28332));
    defparam i15273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1490 (.I0(n27210), .I1(n42312), .I2(n27181), 
            .I3(n42649), .O(n43837));
    defparam i2_3_lut_4_lut_adj_1490.LUT_INIT = 16'h6996;
    SB_LUT4 i34290_4_lut (.I0(n43085), .I1(\FRAME_MATCHER.state [3]), .I2(n84), 
            .I3(n34511), .O(n43097));
    defparam i34290_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i2_3_lut_4_lut_adj_1491 (.I0(n27210), .I1(n42312), .I2(n44027), 
            .I3(\data_out_frame[24] [4]), .O(n43664));
    defparam i2_3_lut_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1492 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n26482), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2524 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1492.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_1493 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n26617), .I3(GND_net), .O(n49));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1493.LUT_INIT = 16'h0202;
    SB_LUT4 i23033_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n26482), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n5_adj_4173), .O(n33593));   // verilog/coms.v(127[12] 300[6])
    defparam i23033_3_lut_4_lut.LUT_INIT = 16'hdfd0;
    SB_LUT4 i1_2_lut_3_lut_adj_1494 (.I0(\FRAME_MATCHER.state [1]), .I1(n26482), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2523 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1494.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_adj_1495 (.I0(\FRAME_MATCHER.state [1]), .I1(n26482), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n52));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1495.LUT_INIT = 16'hfdfd;
    SB_LUT4 i6_4_lut_3_lut (.I0(n42465), .I1(n40658), .I2(n42771), .I3(GND_net), 
            .O(n14_adj_4219));
    defparam i6_4_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1496 (.I0(n42528), .I1(n42465), .I2(\data_out_frame[19] [3]), 
            .I3(GND_net), .O(n40634));
    defparam i1_2_lut_3_lut_adj_1496.LUT_INIT = 16'h9696;
    SB_LUT4 i15258_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n28317));
    defparam i15258_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15259_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n28318));
    defparam i15259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15260_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n28319));
    defparam i15260_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15261_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n28320));
    defparam i15261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15262_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n28321));
    defparam i15262_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15263_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n28322));
    defparam i15263_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32788_2_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n47620));
    defparam i32788_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i15264_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n28323));
    defparam i15264_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15265_3_lut_4_lut (.I0(n8_adj_4373), .I1(n42206), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n28324));
    defparam i15265_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1497 (.I0(n26774), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[5] [2]), .I3(GND_net), .O(n42426));
    defparam i1_2_lut_3_lut_adj_1497.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46730), .I3(n46728), .O(n7_adj_4235));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_3_lut_adj_1498 (.I0(n23831), .I1(\FRAME_MATCHER.i_31__N_2524 ), 
            .I2(n3303), .I3(GND_net), .O(n4_adj_4342));
    defparam i1_3_lut_adj_1498.LUT_INIT = 16'h0808;
    SB_LUT4 i1_3_lut_adj_1499 (.I0(n771), .I1(n85), .I2(n23831), .I3(GND_net), 
            .O(n2_adj_4341));
    defparam i1_3_lut_adj_1499.LUT_INIT = 16'h1010;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46721), .I3(n46719), .O(n7_adj_4234));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1500 (.I0(\FRAME_MATCHER.state [2]), .I1(r_SM_Main_2__N_3516[0]), 
            .I2(tx_active), .I3(GND_net), .O(n6_adj_4161));
    defparam i1_2_lut_3_lut_adj_1500.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46715), .I3(n46713), .O(n7_adj_4233));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46709), .I3(n46707), .O(n7_adj_4232));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46703), .I3(n46701), .O(n7_adj_4231));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46697), .I3(n46695), .O(n7_adj_4230));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46685), .I3(n46683), .O(n7_adj_4225));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46688), .I3(n46686), .O(n7_adj_4228));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i4_4_lut_adj_1501 (.I0(n42385), .I1(\data_in_frame[16] [0]), 
            .I2(n39630), .I3(n42741), .O(n10_adj_4391));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i15250_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n28309));
    defparam i15250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15251_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n28310));
    defparam i15251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1502 (.I0(n52), .I1(n4452), .I2(\FRAME_MATCHER.i_31__N_2524 ), 
            .I3(n3303), .O(n4_c));
    defparam i1_3_lut_4_lut_adj_1502.LUT_INIT = 16'h11f1;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34328 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n49281));
    defparam byte_transmit_counter_0__bdd_4_lut_34328.LUT_INIT = 16'he4aa;
    SB_LUT4 i15252_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n28311));
    defparam i15252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(n23831), .I1(n3183), .I2(GND_net), 
            .I3(GND_net), .O(n1_adj_4386));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h8888;
    SB_LUT4 n49281_bdd_4_lut (.I0(n49281), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n49284));
    defparam n49281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1504 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n26688), .I3(\FRAME_MATCHER.i [1]), .O(n5));
    defparam i1_3_lut_4_lut_adj_1504.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_3_lut_adj_1505 (.I0(n4452), .I1(n52), .I2(n23831), .I3(GND_net), 
            .O(n1_adj_4309));
    defparam i1_3_lut_adj_1505.LUT_INIT = 16'h1010;
    SB_LUT4 i2_2_lut_4_lut_adj_1506 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[11] [1]), 
            .I2(n26999), .I3(\data_in_frame[10] [4]), .O(n10_adj_4157));
    defparam i2_2_lut_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1507 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(n42422), .O(n6_adj_4178));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i15253_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n28312));
    defparam i15253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(\FRAME_MATCHER.state [31]), .I1(n5_adj_4378), 
            .I2(GND_net), .I3(GND_net), .O(n41721));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1509 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [7]), 
            .I2(n10_adj_4391), .I3(\data_in_frame[17] [7]), .O(n40235));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 i15254_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n28313));
    defparam i15254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34323 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n49275));
    defparam byte_transmit_counter_0__bdd_4_lut_34323.LUT_INIT = 16'he4aa;
    SB_LUT4 i15255_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n28314));
    defparam i15255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15256_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n28315));
    defparam i15256_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49275_bdd_4_lut (.I0(n49275), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n49278));
    defparam n49275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15257_3_lut_4_lut (.I0(n8_adj_4374), .I1(n42206), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n28316));
    defparam i15257_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15242_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n28301));
    defparam i15242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15243_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n28302));
    defparam i15243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34318 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n49269));
    defparam byte_transmit_counter_0__bdd_4_lut_34318.LUT_INIT = 16'he4aa;
    SB_LUT4 n49269_bdd_4_lut (.I0(n49269), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n49272));
    defparam n49269_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15244_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n28303));
    defparam i15244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[2] [3]), .I1(n42246), .I2(n42738), 
            .I3(\data_in_frame[5] [3]), .O(n20));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1510 (.I0(n27347), .I1(n42407), .I2(\data_in_frame[3] [1]), 
            .I3(\data_in_frame[0] [7]), .O(n42747));
    defparam i1_2_lut_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1511 (.I0(n27066), .I1(\data_in_frame[5] [5]), 
            .I2(n42566), .I3(GND_net), .O(n42391));
    defparam i1_2_lut_3_lut_adj_1511.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1512 (.I0(\data_in_frame[1] [0]), .I1(n42407), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [7]), .O(n27200));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34313 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n49263));
    defparam byte_transmit_counter_0__bdd_4_lut_34313.LUT_INIT = 16'he4aa;
    SB_LUT4 n49263_bdd_4_lut (.I0(n49263), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n49266));
    defparam n49263_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15245_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n28304));
    defparam i15245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_34421 (.I0(byte_transmit_counter[1]), 
            .I1(n47593), .I2(n47594), .I3(byte_transmit_counter[2]), .O(n49257));
    defparam byte_transmit_counter_1__bdd_4_lut_34421.LUT_INIT = 16'he4aa;
    SB_LUT4 i15246_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n28305));
    defparam i15246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15247_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n28306));
    defparam i15247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1513 (.I0(\FRAME_MATCHER.state_31__N_2624 [3]), 
            .I1(\FRAME_MATCHER.state [0]), .I2(n26622), .I3(\FRAME_MATCHER.state [1]), 
            .O(n8_adj_4112));   // verilog/coms.v(127[12] 300[6])
    defparam i3_3_lut_4_lut_adj_1513.LUT_INIT = 16'h0200;
    SB_LUT4 i15248_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n28307));
    defparam i15248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15249_3_lut_4_lut (.I0(n8_adj_4372), .I1(n42206), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n28308));
    defparam i15249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_428_Select_1_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4275));
    defparam select_428_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_2_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4274));
    defparam select_428_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 n49257_bdd_4_lut (.I0(n49257), .I1(n17_adj_4168), .I2(n16_adj_4167), 
            .I3(byte_transmit_counter[2]), .O(n49260));
    defparam n49257_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_428_Select_3_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4272));
    defparam select_428_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_4_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4270));
    defparam select_428_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_5_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4268));
    defparam select_428_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_6_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4266));
    defparam select_428_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_7_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4264));
    defparam select_428_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_8_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4262));
    defparam select_428_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 select_428_Select_9_i3_2_lut_4_lut (.I0(n2482), .I1(n26617), 
            .I2(n84), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4260));
    defparam select_428_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'h4500;
    uart_tx tx (.CLK_c(CLK_c), .\r_SM_Main_2__N_3513[1] (\r_SM_Main_2__N_3513[1] ), 
            .r_SM_Main({r_SM_Main}), .GND_net(GND_net), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .n42123(n42123), .n27820(n27820), .tx_o(tx_o), .tx_data({tx_data}), 
            .\r_SM_Main_2__N_3516[0] (r_SM_Main_2__N_3516[0]), .n19247(n19247), 
            .n49552(n49552), .n28192(n28192), .tx_active(tx_active), .n4(n4_adj_6), 
            .n28212(n28212), .VCC_net(VCC_net), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.n4(n4_adj_7), .GND_net(GND_net), .r_SM_Main({r_SM_Main_adj_14}), 
            .r_Rx_Data(r_Rx_Data), .\r_SM_Main_2__N_3442[2] (\r_SM_Main_2__N_3442[2] ), 
            .CLK_c(CLK_c), .n27824(n27824), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_11 ), 
            .n26628(n26628), .n33696(n33696), .RX_N_10(RX_N_10), .n42126(n42126), 
            .n41813(n41813), .rx_data_ready(rx_data_ready), .n28224(n28224), 
            .rx_data({rx_data}), .n28182(n28182), .n28181(n28181), .n28180(n28180), 
            .n27784(n27784), .n28179(n28179), .n28178(n28178), .n28177(n28177), 
            .n28176(n28176), .n42185(n42185), .n28215(n28215), .VCC_net(VCC_net), 
            .n26633(n26633), .n4_adj_4(n4_adj_12), .n4_adj_5(n4_adj_13)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (CLK_c, \r_SM_Main_2__N_3513[1] , r_SM_Main, GND_net, 
            \r_Bit_Index[0] , n42123, n27820, tx_o, tx_data, \r_SM_Main_2__N_3516[0] , 
            n19247, n49552, n28192, tx_active, n4, n28212, VCC_net, 
            tx_enable) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output \r_SM_Main_2__N_3513[1] ;
    output [2:0]r_SM_Main;
    input GND_net;
    output \r_Bit_Index[0] ;
    output n42123;
    output n27820;
    output tx_o;
    input [7:0]tx_data;
    input \r_SM_Main_2__N_3516[0] ;
    output n19247;
    input n49552;
    input n28192;
    output tx_active;
    output n4;
    input n28212;
    input VCC_net;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n28096, n19908, n19909;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]n307;
    
    wire n49410, n49356, o_Tx_Serial_N_3544, n3;
    wire [2:0]r_SM_Main_2__N_3510;
    
    wire n28027, n23932;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n3_adj_4108, n49407, n49353, n8, n7, n38612, n38611, 
        n38610, n38609, n38608, n38607, n38606, n38605;
    
    SB_DFFESR r_Clock_Count_1553__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n1), 
            .D(n41[6]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1553__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n1), 
            .D(n41[0]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i6931_3_lut (.I0(n19908), .I1(\r_SM_Main_2__N_3513[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n19909));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6931_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1694_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1694_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2177074_i1_3_lut (.I0(n49410), .I1(n49356), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3544));
    defparam i2177074_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3544), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n42123));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21337_2_lut (.I0(n42123), .I1(\r_SM_Main_2__N_3513[1] ), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3510[0]));
    defparam i21337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1687_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1687_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR r_Clock_Count_1553__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n1), 
            .D(n41[5]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1553__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n1), 
            .D(n41[4]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1553__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n1), 
            .D(n41[3]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n27820), 
            .D(n307[1]), .R(n28027));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n27820), 
            .D(n307[2]), .R(n28027));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n23932), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n19909), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1553__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n1), 
            .D(n41[2]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1553__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n1), 
            .D(n41[1]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4108), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n23932), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n23932), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n23932), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n23932), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n23932), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n23932), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n23932), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i6273_2_lut (.I0(\r_SM_Main_2__N_3516[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n19247));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6273_2_lut.LUT_INIT = 16'h2222;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n49552));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n28192));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n49407));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49407_bdd_4_lut (.I0(n49407), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n49410));
    defparam n49407_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_34426 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n49353));
    defparam r_Bit_Index_0__bdd_4_lut_34426.LUT_INIT = 16'he4aa;
    SB_LUT4 n49353_bdd_4_lut (.I0(n49353), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n49356));
    defparam n49353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[2]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[8]), .I2(n8), 
            .I3(r_Clock_Count[4]), .O(n7));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut (.I0(n7), .I1(r_Clock_Count[5]), .I2(r_Clock_Count[7]), 
            .I3(r_Clock_Count[6]), .O(\r_SM_Main_2__N_3513[1] ));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33570_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3513[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n28096));
    defparam i33570_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR r_Clock_Count_1553__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n1), 
            .D(n41[8]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1553__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n1), 
            .D(n41[7]), .R(n28096));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3513[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 r_Clock_Count_1553_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n38612), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1553_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n38611), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_9 (.CI(n38611), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n38612));
    SB_LUT4 r_Clock_Count_1553_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n38610), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_8 (.CI(n38610), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n38611));
    SB_LUT4 r_Clock_Count_1553_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n38609), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_7 (.CI(n38609), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n38610));
    SB_LUT4 r_Clock_Count_1553_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n38608), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_6 (.CI(n38608), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n38609));
    SB_LUT4 r_Clock_Count_1553_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n38607), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_5 (.CI(n38607), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n38608));
    SB_LUT4 r_Clock_Count_1553_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n38606), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_4 (.CI(n38606), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n38607));
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n28212));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_1553_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n38605), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_3 (.CI(n38605), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n38606));
    SB_LUT4 r_Clock_Count_1553_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1553_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1553_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n38605));
    SB_LUT4 i10676_2_lut_3_lut (.I0(\r_SM_Main_2__N_3513[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4108));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i10676_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3516[0] ), 
            .I3(r_SM_Main[1]), .O(n23932));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3510[0]), .O(n28027));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_850 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3513[1] ), .O(n27820));
    defparam i1_3_lut_4_lut_adj_850.LUT_INIT = 16'h1101;
    SB_LUT4 i6930_3_lut_4_lut (.I0(\r_SM_Main_2__N_3516[0] ), .I1(n42123), 
            .I2(\r_SM_Main_2__N_3513[1] ), .I3(r_SM_Main[1]), .O(n19908));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6930_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n4, GND_net, r_SM_Main, r_Rx_Data, \r_SM_Main_2__N_3442[2] , 
            CLK_c, n27824, \r_Bit_Index[0] , n26628, n33696, RX_N_10, 
            n42126, n41813, rx_data_ready, n28224, rx_data, n28182, 
            n28181, n28180, n27784, n28179, n28178, n28177, n28176, 
            n42185, n28215, VCC_net, n26633, n4_adj_4, n4_adj_5) /* synthesis syn_module_defined=1 */ ;
    output n4;
    input GND_net;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    output \r_SM_Main_2__N_3442[2] ;
    input CLK_c;
    output n27824;
    output \r_Bit_Index[0] ;
    output n26628;
    output n33696;
    input RX_N_10;
    output n42126;
    input n41813;
    output rx_data_ready;
    input n28224;
    output [7:0]rx_data;
    input n28182;
    input n28181;
    input n28180;
    output n27784;
    input n28179;
    input n28178;
    input n28177;
    input n28176;
    input n42185;
    input n28215;
    input VCC_net;
    output n26633;
    output n4_adj_4;
    output n4_adj_5;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_2__N_3448;
    
    wire n47583, n34441;
    wire [7:0]n37;
    
    wire n27894;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n28094;
    wire [2:0]n326;
    
    wire n28029, n26500, n1, n34315, n3, r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_3445;
    
    wire n26492, n10, n8, n43022, n6, n38604, n38603, n38602, 
        n38601, n38600, n38599, n38598;
    
    SB_LUT4 equal_153_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_153_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i32817_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3448[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n47583));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i32817_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n47583), .I1(\r_SM_Main_2__N_3442[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n34441));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_DFFESR r_Clock_Count_1551__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n27894), 
            .D(n37[0]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n27824), 
            .D(n326[1]), .R(n28029));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n27824), 
            .D(n326[2]), .R(n28029));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut (.I0(n26500), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n26628));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20654_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33696));
    defparam i20654_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3448[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n34315), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i1672_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1672_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n42126));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21339_2_lut (.I0(n42126), .I1(\r_SM_Main_2__N_3442[2] ), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3445[0]));
    defparam i21339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1665_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1665_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n34441), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut_adj_847 (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[5]), 
            .I2(r_Clock_Count[7]), .I3(GND_net), .O(n26492));   // verilog/uart_rx.v(68[17:52])
    defparam i2_3_lut_adj_847.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[4]), .I2(n26492), 
            .I3(r_Clock_Count[2]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[1]), .I1(n10), .I2(r_Clock_Count[3]), 
            .I3(GND_net), .O(r_SM_Main_2__N_3448[0]));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i3_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[2]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21245_4_lut (.I0(r_Clock_Count[0]), .I1(n26492), .I2(n8), 
            .I3(r_Clock_Count[4]), .O(\r_SM_Main_2__N_3442[2] ));
    defparam i21245_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i28150_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_3448[0]), 
            .I3(GND_net), .O(n43022));
    defparam i28150_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n43022), .I2(\r_SM_Main_2__N_3442[2] ), 
            .I3(r_SM_Main[1]), .O(n28094));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n41813));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n28224));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1551__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n27894), 
            .D(n37[7]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3448[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i33573_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n27894));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i33573_4_lut.LUT_INIT = 16'h4555;
    SB_DFFESR r_Clock_Count_1551__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n27894), 
            .D(n37[6]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1551__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n27894), 
            .D(n37[5]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1551__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n27894), 
            .D(n37[4]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1551__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n27894), 
            .D(n37[3]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1551__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n27894), 
            .D(n37[2]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1551__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n27894), 
            .D(n37[1]), .R(n28094));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3445[0]), .O(n28029));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_848 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3442[2] ), .O(n27824));
    defparam i1_3_lut_4_lut_adj_848.LUT_INIT = 16'h1101;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n28182));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n28181));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n28180));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i13_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(\r_SM_Main_2__N_3442[2] ), 
            .I3(r_SM_Main[0]), .O(n27784));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h2055;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n28179));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n28178));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n28177));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n28176));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n42185));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1551_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n38604), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1551_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n38603), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1551_add_4_8 (.CI(n38603), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n38604));
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n28215));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1551_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n38602), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1551_add_4_7 (.CI(n38602), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n38603));
    SB_LUT4 r_Clock_Count_1551_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n38601), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1551_add_4_6 (.CI(n38601), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n38602));
    SB_LUT4 r_Clock_Count_1551_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n38600), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1551_add_4_5 (.CI(n38600), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n38601));
    SB_LUT4 r_Clock_Count_1551_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n38599), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1551_add_4_4 (.CI(n38599), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n38600));
    SB_LUT4 r_Clock_Count_1551_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n38598), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1551_add_4_3 (.CI(n38598), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n38599));
    SB_LUT4 r_Clock_Count_1551_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1551_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1551_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n38598));
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3442[2] ), .O(n26500));
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_849 (.I0(n26500), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n26633));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_849.LUT_INIT = 16'heeee;
    SB_LUT4 equal_157_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_157_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_155_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5));   // verilog/uart_rx.v(97[17:39])
    defparam equal_155_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_3_lut (.I0(n42126), .I1(\r_SM_Main_2__N_3442[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n34315));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_3_lut.LUT_INIT = 16'hc7c7;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (CLK_c, \state[3] , n6, GND_net, read, \state[0] , 
            enable_slow_N_4090, n4226, \state[1] , \state[2] , n7, 
            n28191, rw, n41955, data_ready, n41845, n41841, n43002, 
            n43073, n34306, \state_7__N_3987[0] , \state_7__N_4003[3] , 
            \saved_addr[0] , \state[0]_adj_2 , n5538, n33499, sda_enable, 
            scl_enable, n10, n6014, n8, VCC_net, n28202, data, 
            sda_out, n28194, n47597, scl, n26652, n28174, n28170, 
            n28169, n28168, n28167, n28166, n28165, n33700, n4, 
            n4_adj_3, n26657) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    output \state[3] ;
    output n6;
    input GND_net;
    input read;
    output \state[0] ;
    output enable_slow_N_4090;
    output [0:0]n4226;
    output \state[1] ;
    output \state[2] ;
    output n7;
    input n28191;
    output rw;
    input n41955;
    output data_ready;
    input n41845;
    input n41841;
    input n43002;
    output n43073;
    output n34306;
    output \state_7__N_3987[0] ;
    input \state_7__N_4003[3] ;
    output \saved_addr[0] ;
    output \state[0]_adj_2 ;
    output n5538;
    output n33499;
    output sda_enable;
    output scl_enable;
    output n10;
    input n6014;
    input n8;
    input VCC_net;
    input n28202;
    output [7:0]data;
    output sda_out;
    input n28194;
    output n47597;
    output scl;
    output n26652;
    input n28174;
    input n28170;
    input n28169;
    input n28168;
    input n28167;
    input n28166;
    input n28165;
    output n33700;
    output n4;
    output n4_adj_3;
    output n26657;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3889;
    
    wire n27871;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n28048, n26509, n28, n26, n27, n25, enable;
    wire [15:0]n3652;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n37349, n37348, n37347, n37346, n37345, n37344, n37343, 
        n37342, n37341, n37340, n37339, n37338, n37337, n37336, 
        n37335;
    
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[1]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[2]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[3]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[4]), .S(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[5]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[6]), .S(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[7]), .S(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[8]), .S(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[9]), .S(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[10]), .S(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[11]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[12]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[13]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[14]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[15]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i2_2_lut (.I0(\state[3] ), .I1(n26509), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n26509));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_907_Mux_0_i1_4_lut (.I0(read), .I1(n26509), .I2(\state[0] ), 
            .I3(enable_slow_N_4090), .O(n4226[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_907_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n4226[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i33622_2_lut (.I0(n26509), .I1(enable_slow_N_4090), .I2(GND_net), 
            .I3(GND_net), .O(n3652[5]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i33622_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n27871), 
            .D(delay_counter_15__N_3889[0]), .R(n28048));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i15033_2_lut (.I0(n27871), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28048));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15033_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n27871));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i2_2_lut_adj_846 (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut_adj_846.LUT_INIT = 16'heeee;
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n28191));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n41955));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_715_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n3652[5]), 
            .I3(n37349), .O(delay_counter_15__N_3889[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_715_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n3652[5]), 
            .I3(n37348), .O(delay_counter_15__N_3889[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_16 (.CI(n37348), .I0(delay_counter[14]), .I1(n3652[5]), 
            .CO(n37349));
    SB_LUT4 add_715_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n3652[5]), 
            .I3(n37347), .O(delay_counter_15__N_3889[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_15 (.CI(n37347), .I0(delay_counter[13]), .I1(n3652[5]), 
            .CO(n37348));
    SB_LUT4 add_715_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n3652[5]), 
            .I3(n37346), .O(delay_counter_15__N_3889[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_14 (.CI(n37346), .I0(delay_counter[12]), .I1(n3652[5]), 
            .CO(n37347));
    SB_LUT4 add_715_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n3652[5]), 
            .I3(n37345), .O(delay_counter_15__N_3889[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_13 (.CI(n37345), .I0(delay_counter[11]), .I1(n3652[5]), 
            .CO(n37346));
    SB_LUT4 add_715_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n3652[5]), 
            .I3(n37344), .O(delay_counter_15__N_3889[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_12 (.CI(n37344), .I0(delay_counter[10]), .I1(n3652[5]), 
            .CO(n37345));
    SB_LUT4 add_715_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n3652[5]), 
            .I3(n37343), .O(delay_counter_15__N_3889[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_11 (.CI(n37343), .I0(delay_counter[9]), .I1(n3652[5]), 
            .CO(n37344));
    SB_LUT4 add_715_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n3652[5]), 
            .I3(n37342), .O(delay_counter_15__N_3889[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_10 (.CI(n37342), .I0(delay_counter[8]), .I1(n3652[5]), 
            .CO(n37343));
    SB_LUT4 add_715_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n3652[5]), 
            .I3(n37341), .O(delay_counter_15__N_3889[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_9 (.CI(n37341), .I0(delay_counter[7]), .I1(n3652[5]), 
            .CO(n37342));
    SB_LUT4 add_715_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n3652[5]), 
            .I3(n37340), .O(delay_counter_15__N_3889[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_8 (.CI(n37340), .I0(delay_counter[6]), .I1(n3652[5]), 
            .CO(n37341));
    SB_LUT4 add_715_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n3652[5]), 
            .I3(n37339), .O(delay_counter_15__N_3889[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_7 (.CI(n37339), .I0(delay_counter[5]), .I1(n3652[5]), 
            .CO(n37340));
    SB_LUT4 add_715_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n3652[5]), 
            .I3(n37338), .O(delay_counter_15__N_3889[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_6 (.CI(n37338), .I0(delay_counter[4]), .I1(n3652[5]), 
            .CO(n37339));
    SB_LUT4 add_715_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n3652[5]), 
            .I3(n37337), .O(delay_counter_15__N_3889[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_5 (.CI(n37337), .I0(delay_counter[3]), .I1(n3652[5]), 
            .CO(n37338));
    SB_LUT4 add_715_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n3652[5]), 
            .I3(n37336), .O(delay_counter_15__N_3889[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_4 (.CI(n37336), .I0(delay_counter[2]), .I1(n3652[5]), 
            .CO(n37337));
    SB_LUT4 add_715_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n3652[5]), 
            .I3(n37335), .O(delay_counter_15__N_3889[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_3 (.CI(n37335), .I0(delay_counter[1]), .I1(n3652[5]), 
            .CO(n37336));
    SB_LUT4 add_715_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n3652[5]), 
            .I3(GND_net), .O(delay_counter_15__N_3889[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n3652[5]), 
            .CO(n37335));
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n41845));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n41841));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i28198_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n43002), 
            .I3(enable_slow_N_4090), .O(n43073));   // verilog/eeprom.v(51[5:9])
    defparam i28198_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 i21263_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4090), 
            .I3(GND_net), .O(n34306));   // verilog/eeprom.v(51[5:9])
    defparam i21263_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    i2c_controller i2c (.\state_7__N_3987[0] (\state_7__N_3987[0] ), .enable_slow_N_4090(enable_slow_N_4090), 
            .GND_net(GND_net), .CLK_c(CLK_c), .\state_7__N_4003[3] (\state_7__N_4003[3] ), 
            .\saved_addr[0] (\saved_addr[0] ), .\state[1] (state[1]), .\state[2] (\state[2] ), 
            .\state[0] (\state[0]_adj_2 ), .\state[3] (\state[3] ), .n5538(n5538), 
            .n33499(n33499), .enable(enable), .sda_enable(sda_enable), 
            .scl_enable(scl_enable), .n10(n10), .n6014(n6014), .n8(n8), 
            .VCC_net(VCC_net), .n28202(n28202), .data({data}), .sda_out(sda_out), 
            .n28194(n28194), .n47597(n47597), .scl(scl), .n26652(n26652), 
            .n28174(n28174), .n28170(n28170), .n28169(n28169), .n28168(n28168), 
            .n28167(n28167), .n28166(n28166), .n28165(n28165), .n33700(n33700), 
            .n4(n4), .n4_adj_1(n4_adj_3), .n26657(n26657)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (\state_7__N_3987[0] , enable_slow_N_4090, GND_net, 
            CLK_c, \state_7__N_4003[3] , \saved_addr[0] , \state[1] , 
            \state[2] , \state[0] , \state[3] , n5538, n33499, enable, 
            sda_enable, scl_enable, n10, n6014, n8, VCC_net, n28202, 
            data, sda_out, n28194, n47597, scl, n26652, n28174, 
            n28170, n28169, n28168, n28167, n28166, n28165, n33700, 
            n4, n4_adj_1, n26657) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state_7__N_3987[0] ;
    output enable_slow_N_4090;
    input GND_net;
    input CLK_c;
    input \state_7__N_4003[3] ;
    output \saved_addr[0] ;
    output \state[1] ;
    output \state[2] ;
    output \state[0] ;
    output \state[3] ;
    output n5538;
    output n33499;
    input enable;
    output sda_enable;
    output scl_enable;
    output n10;
    input n6014;
    input n8;
    input VCC_net;
    input n28202;
    output [7:0]data;
    output sda_out;
    input n28194;
    output n47597;
    output scl;
    output n26652;
    input n28174;
    input n28170;
    input n28169;
    input n28168;
    input n28167;
    input n28166;
    input n28165;
    output n33700;
    output n4;
    output n4_adj_1;
    output n26657;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n119;
    
    wire n27937;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n28142, enable_slow_N_4089;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n28097, n11, n11_adj_4091, n5, n47587, n47527, n11_adj_4092, 
        n47646, n10_c, n15, n11_adj_4093, n34105, state_7__N_3986, 
        n5531, n11_adj_4094, n33885, i2c_clk_N_4076, n7, n33, n37, 
        n28025, n34, n39, n10_adj_4095, n47621, n42037, n19389, 
        n5909, scl_enable_N_4077, n41891, sda_out_adj_4096, n34355, 
        n27835, n10_adj_4097, n15_adj_4099, n43008, n12, n44815, 
        n38648, n38647, n38646, n38645, n38644, n37546, n37545, 
        n37544, n37543, n37542, n37541, n37540;
    
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27937), .D(n119[6]), 
            .R(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27937), .D(n119[5]), 
            .R(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i33620_2_lut (.I0(\state_7__N_3987[0] ), .I1(enable_slow_N_4090), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4089));   // verilog/i2c_controller.v(62[6:32])
    defparam i33620_2_lut.LUT_INIT = 16'h7777;
    SB_DFFSR counter2_1555_1556__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n28097));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27937), .D(n119[4]), 
            .R(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27937), .D(n119[3]), 
            .R(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27937), .D(n119[2]), 
            .S(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27937), .D(n119[1]), 
            .S(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_4_lut (.I0(n11), .I1(n11_adj_4091), .I2(\state_7__N_4003[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'h5755;
    SB_LUT4 i32670_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n47587));   // verilog/i2c_controller.v(198[28:35])
    defparam i32670_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i32725_4_lut (.I0(n47587), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n47527));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i32725_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 i32967_4_lut (.I0(n47527), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(n11_adj_4092), .O(n47646));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i32967_4_lut.LUT_INIT = 16'h0322;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_c));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i33922_3_lut (.I0(n5538), .I1(n15), .I2(n11_adj_4093), .I3(GND_net), 
            .O(n34105));
    defparam i33922_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i33579_4_lut (.I0(state_7__N_3986), .I1(n5531), .I2(n11_adj_4094), 
            .I3(n33499), .O(n5538));
    defparam i33579_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i33753_2_lut (.I0(\state_7__N_4003[3] ), .I1(n11_adj_4091), 
            .I2(GND_net), .I3(GND_net), .O(n33885));
    defparam i33753_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n28097), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4076));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_841 (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_841.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n28025));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_842 (.I0(n34), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i1_2_lut_adj_842.LUT_INIT = 16'heeee;
    SB_LUT4 i21429_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_3986));
    defparam i21429_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i32966_4_lut (.I0(n10_adj_4095), .I1(n10_c), .I2(\state_7__N_4003[3] ), 
            .I3(enable), .O(n47621));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i32966_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut_adj_843 (.I0(\state[1] ), .I1(n7), .I2(n47621), .I3(\state[0] ), 
            .O(n42037));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_843.LUT_INIT = 16'ha088;
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n5909), 
            .D(n19389), .S(n28025));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4093));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4076));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4077));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n5538), .D(n33885), 
            .S(n34105));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4096), .C(i2c_clk), .E(n41891), 
            .D(n47646));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n5538), .D(n5), 
            .S(n34355));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27937), .D(n119[0]), 
            .S(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE enable_slow_120 (.Q(\state_7__N_3987[0] ), .C(CLK_c), .E(n27835), 
            .D(enable_slow_N_4089));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4097));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4097), .I2(counter2[0]), 
            .I3(GND_net), .O(n28097));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_102_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4095));   // verilog/i2c_controller.v(44[32:47])
    defparam equal_102_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28136_2_lut (.I0(\state_7__N_4003[3] ), .I1(n15_adj_4099), 
            .I2(GND_net), .I3(GND_net), .O(n43008));
    defparam i28136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n5531));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n5531), .I1(n43008), .I2(n6014), .I3(n37), 
            .O(n27937));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n28202));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27937), .D(n119[7]), 
            .R(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1856_2_lut (.I0(sda_out_adj_4096), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i1856_2_lut.LUT_INIT = 16'h8888;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n28194));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n5538), .D(n42037), 
            .S(n44815));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i32696_3_lut_4_lut (.I0(n11_adj_4094), .I1(n11_adj_4093), .I2(enable_slow_N_4090), 
            .I3(\state_7__N_3987[0] ), .O(n47597));
    defparam i32696_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 counter2_1555_1556_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n38648), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1555_1556_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1555_1556_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n38647), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1555_1556_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1555_1556_add_4_6 (.CI(n38647), .I0(GND_net), .I1(counter2[4]), 
            .CO(n38648));
    SB_LUT4 counter2_1555_1556_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n38646), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1555_1556_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1555_1556_add_4_5 (.CI(n38646), .I0(GND_net), .I1(counter2[3]), 
            .CO(n38647));
    SB_LUT4 counter2_1555_1556_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n38645), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1555_1556_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1555_1556_add_4_4 (.CI(n38645), .I0(GND_net), .I1(counter2[2]), 
            .CO(n38646));
    SB_LUT4 counter2_1555_1556_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n38644), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1555_1556_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1555_1556_add_4_3 (.CI(n38644), .I0(GND_net), .I1(counter2[1]), 
            .CO(n38645));
    SB_LUT4 counter2_1555_1556_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1555_1556_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1555_1556_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n38644));
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n37546), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n37545), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n37545), .I0(counter[6]), .I1(VCC_net), 
            .CO(n37546));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n37544), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n37544), .I0(counter[5]), .I1(VCC_net), 
            .CO(n37545));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n37543), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n37543), .I0(counter[4]), .I1(VCC_net), 
            .CO(n37544));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n37542), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n37542), .I0(counter[3]), .I1(VCC_net), 
            .CO(n37543));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n37541), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n37541), .I0(counter[2]), .I1(VCC_net), 
            .CO(n37542));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n37540), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n37540), .I0(counter[1]), .I1(VCC_net), 
            .CO(n37541));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n37540));
    SB_LUT4 i33803_3_lut_4_lut (.I0(n11_adj_4094), .I1(n11_adj_4093), .I2(n15_adj_4099), 
            .I3(n5538), .O(n34355));
    defparam i33803_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i20559_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i20559_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4091));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 equal_102_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4090));
    defparam equal_102_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_844 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n26652));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_844.LUT_INIT = 16'heeee;
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n28174));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n28170));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n28169));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n28168));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n28167));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n28166));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n28165));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1555_1556__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n28097));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1555_1556__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n28097));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1555_1556__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n28097));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1555_1556__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n28097));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1555_1556__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n28097));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 state_7__I_0_138_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4094));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_138_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i20658_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33700));
    defparam i20658_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_161_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_161_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_163_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_163_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_845 (.I0(n15), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n26657));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_845.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28101_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n43008), .O(n28142));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i28101_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 state_7__I_0_143_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i33627_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n41891));
    defparam i33627_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i21412_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(n15_adj_4099), .O(scl_enable_N_4077));
    defparam i21412_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i22_3_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n11_adj_4092));
    defparam i22_3_lut_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 equal_104_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15_adj_4099));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_104_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i33925_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n5538), .O(n44815));
    defparam i33925_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 i21232_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33499));
    defparam i21232_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(\state_7__N_3987[0] ), .I2(enable_slow_N_4090), 
            .I3(GND_net), .O(n27835));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i33633_4_lut_4_lut (.I0(\state[2] ), .I1(n11_adj_4092), .I2(\state[1] ), 
            .I3(n39), .O(n5909));
    defparam i33633_4_lut_4_lut.LUT_INIT = 16'hef00;
    SB_LUT4 i33624_2_lut_3_lut (.I0(\state[2] ), .I1(n11_adj_4092), .I2(\state[0] ), 
            .I3(GND_net), .O(n19389));
    defparam i33624_2_lut_3_lut.LUT_INIT = 16'h0404;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n48297, VCC_net, INHA_c, clk32MHz, n26499, pwm_counter, 
            GND_net, n26497) /* synthesis syn_module_defined=1 */ ;
    input n48297;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n26499;
    output [31:0]pwm_counter;
    input GND_net;
    input n26497;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n43658, n18, n24, n22, n26, n21, pwm_counter_31__N_711;
    wire [31:0]n133;
    
    wire n38566, n38565, n38564, n38563, n38562, n38561, n38560, 
        n38559, n38558, n38557, n38556, n38555, n38554, n38553, 
        n38552, n38551, n38550, n38549, n38548, n38547, n38546, 
        n38545, n38544, n38543, n38542, n38541, n38540, n38539, 
        n38538, n38537, n38536;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n48297), 
            .R(n26499));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n43658));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n43658), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n18));
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[22]), .I2(pwm_counter[14]), 
            .I3(pwm_counter[18]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(pwm_counter[21]), .I1(n26497), .I2(pwm_counter[16]), 
            .I3(pwm_counter[12]), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(pwm_counter[15]), .I1(n24), .I2(n18), .I3(pwm_counter[19]), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_2_lut (.I0(pwm_counter[11]), .I1(pwm_counter[20]), .I2(GND_net), 
            .I3(GND_net), .O(n21));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20773_4_lut (.I0(n21), .I1(pwm_counter[31]), .I2(n26), .I3(n22), 
            .O(pwm_counter_31__N_711));   // verilog/pwm.v(18[8:40])
    defparam i20773_4_lut.LUT_INIT = 16'h3332;
    SB_DFFSR pwm_counter_1548__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n133[10]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n133[11]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n133[12]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n133[13]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n133[14]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n133[15]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n133[16]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n133[17]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n133[18]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n133[19]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n133[20]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n133[21]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n133[22]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1548__i31 (.Q(pwm_counter[31]), .C(clk32MHz), .D(n133[31]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_1548_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[31]), 
            .I3(n38566), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1548_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n38565), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_32 (.CI(n38565), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n38566));
    SB_LUT4 pwm_counter_1548_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n38564), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_31 (.CI(n38564), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n38565));
    SB_LUT4 pwm_counter_1548_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n38563), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_30 (.CI(n38563), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n38564));
    SB_LUT4 pwm_counter_1548_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n38562), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_29 (.CI(n38562), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n38563));
    SB_LUT4 pwm_counter_1548_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n38561), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_28 (.CI(n38561), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n38562));
    SB_LUT4 pwm_counter_1548_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n38560), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_27 (.CI(n38560), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n38561));
    SB_LUT4 pwm_counter_1548_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n38559), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_26 (.CI(n38559), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n38560));
    SB_LUT4 pwm_counter_1548_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n38558), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_25 (.CI(n38558), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n38559));
    SB_LUT4 pwm_counter_1548_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n38557), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_24 (.CI(n38557), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n38558));
    SB_LUT4 pwm_counter_1548_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n38556), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_23 (.CI(n38556), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n38557));
    SB_LUT4 pwm_counter_1548_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n38555), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_22 (.CI(n38555), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n38556));
    SB_LUT4 pwm_counter_1548_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n38554), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_21 (.CI(n38554), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n38555));
    SB_LUT4 pwm_counter_1548_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n38553), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_20 (.CI(n38553), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n38554));
    SB_LUT4 pwm_counter_1548_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n38552), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_19 (.CI(n38552), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n38553));
    SB_LUT4 pwm_counter_1548_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n38551), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_18 (.CI(n38551), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n38552));
    SB_LUT4 pwm_counter_1548_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n38550), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_17 (.CI(n38550), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n38551));
    SB_LUT4 pwm_counter_1548_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n38549), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_16 (.CI(n38549), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n38550));
    SB_LUT4 pwm_counter_1548_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n38548), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_15 (.CI(n38548), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n38549));
    SB_LUT4 pwm_counter_1548_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n38547), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_14 (.CI(n38547), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n38548));
    SB_LUT4 pwm_counter_1548_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n38546), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_13 (.CI(n38546), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n38547));
    SB_LUT4 pwm_counter_1548_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n38545), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_12 (.CI(n38545), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n38546));
    SB_LUT4 pwm_counter_1548_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n38544), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_11 (.CI(n38544), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n38545));
    SB_LUT4 pwm_counter_1548_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n38543), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_10 (.CI(n38543), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n38544));
    SB_LUT4 pwm_counter_1548_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n38542), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_9 (.CI(n38542), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n38543));
    SB_LUT4 pwm_counter_1548_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n38541), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_8 (.CI(n38541), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n38542));
    SB_LUT4 pwm_counter_1548_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n38540), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_7 (.CI(n38540), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n38541));
    SB_LUT4 pwm_counter_1548_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n38539), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_6 (.CI(n38539), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n38540));
    SB_LUT4 pwm_counter_1548_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n38538), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_5 (.CI(n38538), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n38539));
    SB_LUT4 pwm_counter_1548_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n38537), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_4 (.CI(n38537), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n38538));
    SB_LUT4 pwm_counter_1548_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n38536), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_3 (.CI(n38536), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n38537));
    SB_LUT4 pwm_counter_1548_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1548_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1548_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n38536));
    
endmodule
