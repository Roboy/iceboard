// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Sep  8 14:33:26 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    
    wire n37306, n37307;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    
    wire n59719, n59718;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n59285, n25890, data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(352[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(360[15:20])
    
    wire pwm_setpoint_23__N_207, n12454, n12458, n12460, n12464, n12466, 
        n12470, n12472, n12476, n12478, n12482, n12484, n59284, 
        n260, n12490, n294, n298, n299, n300, n301, n302, n303, 
        n304, n305, n306, n307, n308, n309, n625, n623, n622, 
        n621, n59283, n59282, n58901;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n71386, n28392;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, GLC_N_400, 
        dti_N_404, RX_N_2, n1744, n1742;
    wire [31:0]motor_state_23__N_91;
    wire [32:0]encoder0_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
        n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        read_N_409, n4, n1319, n59717, n59281, n44741, n59716, 
        n59715, n59714, n59713, n71380, n1784, n1786, n1788, n1790, 
        n1792, n1794, n1796;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n1822, n1824;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [10:0]t0;   // verilog/neopixel.v(10[12:14])
    wire [1:0]state;   // verilog/neopixel.v(19[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(20[11:18])
    wire [5:0]color_bit_N_502;
    
    wire n58900, n59712, n59280, n59279, n59711, n25, n24, n23, 
        n22, n21, n59278, n59710, n59709, n71728, n20, n19, 
        n19_adj_5707, n17, n16, n15, n13, n12, n11, n10, n9, 
        n18, n17_adj_5708, n2821, n16_adj_5709;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n15_adj_5710, n14, n13_adj_5711, n59277, n2, n32, n31, 
        n30, n29, n28, n27, n26, n14_adj_5712, n15_adj_5713, n16_adj_5714, 
        n17_adj_5715, n18_adj_5716, n19_adj_5717, n20_adj_5718, n21_adj_5719, 
        n22_adj_5720, n23_adj_5721, n24_adj_5722, n25_adj_5723, n25_adj_5724, 
        n24_adj_5725, n23_adj_5726, n22_adj_5727, n21_adj_5728, n20_adj_5729, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active, n19_adj_5730, n18_adj_5731, n17_adj_5732, n16_adj_5733, 
        n15_adj_5734, n14_adj_5735, n13_adj_5736, n12_adj_5737;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n71722, n4930, n4929, n4928, 
        n4908, n4907, n4909, n4910, n4911, n4912, n4913, n4914, 
        n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
        n4923, n4924, n4925, n4926, n4927, n4_adj_5738, n3476, 
        n2874, n11_adj_5739, n10_adj_5740, n9_adj_5741, n78546, n8, 
        n59708, n59707, n35782, n59706, n71716, n1, n59705, n59704, 
        n69651, n66705, n66703, n66704, n29359, n66702, n66701, 
        n66578, n66700, n66699, n66698, n66697, n66696, n66695, 
        n66694, n66693, n66692, n66691, n66690, n66689, n66688, 
        n66687, n66686, n66685, n66684, n66683, n66682, n66681, 
        n66680, n66679, n66678, n66677, n66676, n66675, n66674, 
        n66673, n66672, n66671, n66670, n66669, n66668, n66667, 
        n66666, n66665, n66664, n66663, n66662, n66661, n66660, 
        n66659, n66658, n66657, n66656, n66655, n66654, n66653, 
        n66652, n66651, n66650, n66649, n66648, n66647, n66646, 
        n66645, n66644, n66643, n66642, n66581, n66582, n66583, 
        n66584, n66585, n66586, n66587, n29288, n66589, n66590, 
        n66591, n66592, n66593, n66594, n66595, n66596, n66579, 
        n29278, n66597, n66598, n66599, n66600, n66601, n66602, 
        n29271, n66603, n66604, n66605, n66606, n66607, n66608, 
        n66577, n29263, n66609, n29261, n66610, n66611, n66612, 
        n66613, n66614, n66615, n66616, n29253, n66617, n29251, 
        n66618, n66619, n66620, n66621, n66622, n66623, n29244, 
        n29243, n66624, n66625, n66626, n66627, n66628, n66629, 
        n29236, n29235, n66588, n66630, n29232, n29231, n66631, 
        n66632, n66634, n66635, n66636, n29224, n66580, n66637, 
        n66638, n66639, n66640, n66641, n69831, n29178, n59703, 
        n59702, n59701, n6, n67194, n59053, n59052, n58899, n59051, 
        n59050, n58898, n58897, n4_adj_5742, n59700, n59699, n71332, 
        n71326, n59698, n59697, n71320, n79447, n59696, n59049, 
        n59695, n59694, n59048, n59693, n59259, n58884, n59047, 
        n59258, n59046, n71314, n59045, n59257, n59044, n59692, 
        n59691, n59256, n59043, n7, n6_adj_5743, n7_adj_5744, n6_adj_5745, 
        n5, n4_adj_5746, n59255, n59042, n3, n2_adj_5747, n8_adj_5748, 
        n71308, n6_adj_5749, n71302, n71298, n59041, n71294, n59254, 
        n59040, n58896, n15_adj_5750, n71292, n8_adj_5751, n71282, 
        n59039, n78848, n59253, n71276, n59038, Kp_23__N_1389, n16_adj_5752, 
        n71270, n71264, n77825, n59690, n59689, n59252, n68753, 
        n59688, n59687, n71258, n68558, \FRAME_MATCHER.i_31__N_2509 , 
        n71252, n30193, n30190, n71250, n30187, n30184, n30181, 
        n45282, n30178, n30175, n30172, n30169, n30166, n30163, 
        n30160, n30157, n30154, n30151, n30148, n30145, n30141, 
        n30138, n30135, n30132, n30129, n30126, n30123, n30119, 
        n30118, n30117, n30116, n30115, n30114, n30113, n30112, 
        n30111, n30110, n30109, n30108, n30107, n59686, n59251, 
        n30013, n30012, n30008, n30007, n30003, n30002, n30001, 
        n30000, n29999, n29998, n29997, n29996, n29995, n29994, 
        n29993, n29991, n29990, n29989, n29988, n29987, n29986, 
        n29984, n29983, n45466, n29979, n29976, n29975, n29974, 
        n29973, n29972, n29970, n29969, n29968, n29967, n29966, 
        n29965, n29961, n29960, n29959, n29958, n29956, n29947, 
        n29943, n29941, n29937, n29936, n29934, n45456, n45352, 
        n45450, n29915, n29914, n45448, n29910, n45446, n29906, 
        n45438, n45432, n45428, n45424, n29872, n65964, n65966, 
        n29863, n29845, n29842, n29839, n29836, n29833, n45436, 
        n45330, n29830, n29827, n45440, n29824, n45462, n29821, 
        n68436, n29818, n29815, n29812, n45526, n29809, n29806, 
        n45516, n29803, n45514, n29800, n7_adj_5753, n6_adj_5754, 
        n5_adj_5755, n4_adj_5756, n22_adj_5757, n77535, n19_adj_5758, 
        n17_adj_5759, n16_adj_5760, n15_adj_5761, n31093, n31088, 
        n71236, n13_adj_5762, n11_adj_5763, n9_adj_5764, n8_adj_5765, 
        n7_adj_5766, n6_adj_5767, n5_adj_5768, n4_adj_5769, n71232, 
        n67800, n30_adj_5770, n23_adj_5771, n22_adj_5772, n21_adj_5773, 
        n19_adj_5774, n17_adj_5775, n16_adj_5776, n15_adj_5777, n13_adj_5778, 
        n11_adj_5779, n10_adj_5780, n9_adj_5781, n8_adj_5782, n7_adj_5783, 
        n6_adj_5784, n4_adj_5785, n16_adj_5786, n65962, n69799, n69075, 
        n31046, n31039, n31038, n31034, n31031, n31023, n31022, 
        n71220, n4_adj_5787, n4_adj_5788, n11_adj_5789, n30883, n71214, 
        n30873, n59685, n59684, n59683, n59682, n71212, n59681, 
        n59680, n30786, n30785, n30781, n30779, n30767, n59679, 
        n59678, n77533, control_update, n30762, n59677, n59676, 
        n59675, n59674;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n59673, n30758, n30751, n59672, n59671, n30748, n45398, 
        n59670, n59669, n71206, n30740, n105, n12452, n30734, 
        n239, n247, n258, n284, n291, n299_adj_5790, n313, n322, 
        n336, n337, n339, n340, n342, n343, n344, n345, n346, 
        n347, n348, n349, n350, n351, n352, n353, n354, n355, 
        n356, n357, n358, n359, n460, n461, n462, n467, n475, 
        n486, n5220, n71200, n5217, n29797, n59250, n30727, n59668, 
        n59667, n29794, n77191, n59666, n59665, n3165, n59664, 
        n59663, n77183, n59662, n59661, n5_adj_5791, n30714, n30713, 
        n30712, n30711, n30710, n59660, n11_adj_5792, n30709, n30708, 
        n30707, n59659;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3833, n30697, n30696, n30695, 
        position_31__N_3836, n30694, n59658, n59657, n59656, n59655, 
        n59654, n59653, n30693, n30692, n30691, n30690, n71578, 
        n23188, n59652, n59651, n15_adj_5793, n59650, n59649, n59648, 
        n59647, n30678, n30677, n59646, n59645, n59644;
    wire [1:0]a_new_adj_6010;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_6011;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5796, b_prev_adj_5797, debounce_cnt_N_3833_adj_5798, 
        n30676, n30675, n30674, n30673, position_31__N_3836_adj_5799, 
        n72377, n30672, n30671, n12_adj_5800, n11_adj_5801, n10_adj_5802, 
        n4_adj_5803, n3_adj_5804, n2_adj_5805, n30670, n30669, n30668, 
        n30667;
    wire [7:0]data_adj_6024;   // verilog/eeprom.v(23[12:16])
    
    wire n30666;
    wire [7:0]state_7__N_3918;
    
    wire n67730, n291_adj_5806, n71188, n5_adj_5807, n6903, n69884, 
        n30632, n45504;
    wire [15:0]data_adj_6031;   // verilog/tli4970.v(27[14:18])
    
    wire n37117, n30619, n30616, n59612, n59611, n15_adj_5816, n30603, 
        n30593, n30589, n30588, n5_adj_5817, n30585, n30584, n59610, 
        n30583, n59609, n30582, n12488, n59608, n30581, n30580, 
        n30579, n59607, n30578, state_7__N_4319, n30577, n71182, 
        n29775, n45500, n9_adj_5818, n8_adj_5819, n7_adj_5820, n6_adj_5821, 
        n5_adj_5822, n30576, n30555, n71574, n59606, n59605, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n45464, n45283;
    wire [24:0]o_Rx_DV_N_3488;
    wire [2:0]r_SM_Main_adj_6047;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_6048;   // verilog/uart_tx.v(33[16:29])
    
    wire n30517, n30516, n71176, n30515, n30514, n23025, n59604, 
        n59603, n77531, n30513, n30512, n30511, n30510, n30509, 
        n30508, n30507, n59602, n30505, n30503, n30502, n30501, 
        n30500, n30499, n30498, n30497, n30496, n30495, n59601;
    wire [7:0]state_adj_6057;   // verilog/i2c_controller.v(33[12:17])
    
    wire n78034, n59600, enable_slow_N_4213, n8_adj_5834, n30490, 
        n30489, n59599, n45494, n71170, n30481, n8_adj_5835;
    wire [7:0]state_7__N_4110;
    
    wire n30479, n6707, n30469, n59598, n59597;
    wire [7:0]state_7__N_4126;
    
    wire n30458, n59596, n71164, n30432, n29763, n29759, n59595, 
        n59594, n42994, n59593, n59592, n59591, n731, n71158, 
        n36832, n7761, n7760, n7759, n7758, n7757, n7756, n76681, 
        n828, n829, n830, n831, n832, n833, n834, n861, n896, 
        n897, n898, n899, n900, n901, n927, n928, n929, n930, 
        n931, n932, n933, n934, n935, n936, n937, n938, n939, 
        n940, n941, n942, n943, n944, n945, n946, n947, n948, 
        n949, n950, n951, n952, n953, n954, n955, n956, n957, 
        n960, n71150, n995, n996, n997, n998, n999, n1000, n1001, 
        n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
        n1059, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
        n1100, n1101, n71144, n1125, n1126, n1127, n1128, n1129, 
        n1130, n1131, n1132, n1133, n78873, n1158, n1193, n1194, 
        n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1224_adj_5836, 
        n1225_adj_5837, n1226_adj_5838, n1227_adj_5839, n1228_adj_5840, 
        n1229_adj_5841, n1230_adj_5842, n1231_adj_5843, n1232_adj_5844, 
        n1233_adj_5845, n78888, n1257, n1292, n1293, n1294, n1295, 
        n1296, n1297, n1298, n1299, n1300, n1301, n1323, n1324, 
        n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
        n1333, n71136, n1356, n1391, n1392, n1393, n1394, n1395, 
        n1396, n1397, n1398, n1399, n1400, n1401, n1422, n1423, 
        n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
        n1432, n1433, n1455, n1489, n1490, n1491, n1492, n1493, 
        n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
        n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
        n1529, n1530, n1531, n1532, n1533, n1554, n1589, n1590, 
        n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
        n1599, n1600, n1601, n71130, n67637, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n67635, n1653, n59549, n67633, n59548, 
        n41637, n82, n89, n41654, n1688, n1689, n1690, n1691, 
        n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
        n1700, n1701, n67631, n41669, n1719, n1720, n1721, n1722, 
        n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
        n1731, n1732, n1733, n79, n67628, n59547, n1752, n59546, 
        n59545, n71126, n67625, n1787, n1788_adj_5846, n1789, n1790_adj_5847, 
        n1791, n1792_adj_5848, n1793, n1794_adj_5849, n1795, n1796_adj_5850, 
        n1797, n1798, n1799, n1800, n1801, n1818, n1819, n1820, 
        n1821, n1822_adj_5851, n1823, n1824_adj_5852, n1825, n1826, 
        n1827, n1828, n1829, n1830, n1831, n1832, n1833, n59249, 
        n1851, n59544, n59543, n59542, n59541, n59540, n59539, 
        n59538, n59537, n1885, n1886, n1887, n1888, n1889, n1890, 
        n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
        n1899, n1900, n1901, n1917, n1918, n1919, n1920, n1921, 
        n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
        n1930, n1931, n1932, n1933, n78377, n1950, n71118, n1985, 
        n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
        n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, 
        n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
        n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, 
        n2032, n2033, n44559, n2049, n12_adj_5853, n2084, n2085, 
        n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, 
        n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, 
        n59536, n59535, n59248, n2115, n2116, n2117, n2118, n2119, 
        n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
        n2128, n2129, n2130, n2131, n2132, n2133, n59247, n59037, 
        n59534, n2148, n59533, n59532, n59246, n71112, n59531, 
        n59530, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
        n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
        n2198, n2199, n2200, n2201, n59529, n59245, n59244, n2214, 
        n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
        n2231, n2232, n2233, n59036, n59035, n2247, n59243, n2281, 
        n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
        n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
        n2298, n2299, n2300, n2301, n2313, n2314, n2315, n2316, 
        n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
        n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
        n2333, n59242, n2346, n59241, n59240, n59034, n59033, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n59239, n2445, n59238, n2480, n2481, 
        n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, 
        n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, 
        n2498, n2499, n2500, n2501, n59509, n2511, n2512, n2513, 
        n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, 
        n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, 
        n2530, n2531, n2532, n2533, n2544, n59508, n59507, n59506, 
        n59505, n59237, n59504, n2579, n2580, n2581, n2582, n2583, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
        n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
        n2600, n2601, n59503, n2610, n2611, n2612, n2613, n2614, 
        n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
        n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
        n2631, n2632, n2633, n2643, n59502, n59501, n59500, n59499, 
        n59498, n59497, n59236, n59496, n59495, n2677, n2678, 
        n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
        n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
        n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2709, 
        n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
        n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, 
        n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
        n2742, n59494, n59235, n59493, n59032, n2776, n2777, n2778, 
        n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
        n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, 
        n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2808, 
        n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
        n2817, n2818, n2819, n2820, n2821_adj_5854, n2822, n2823, 
        n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
        n2832, n2833, n59234, n2841, n59492, n59491, n2875, n2876, 
        n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
        n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
        n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
        n2901, n59490, n59233, n2907, n2908, n2909, n2910, n2911, 
        n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, 
        n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, 
        n2928, n2929, n2930, n2931, n2932, n2933, n59031, n78616, 
        n2940, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
        n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
        n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
        n2998, n2999, n3000, n3001, n3006, n3007, n3008, n3009, 
        n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
        n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
        n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
        n78970, n3039, n59232, n3074, n3075, n3076, n3077, n3078, 
        n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
        n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
        n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3105, 
        n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
        n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
        n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
        n3130, n3131, n3132, n3133, n79004, n3138, n59231, n27_adj_5855, 
        n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, 
        n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
        n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
        n3197, n3198, n3199, n3200, n3201, n3204, n3205, n3206, 
        n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
        n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
        n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
        n3231, n3232, n3233, n3237, n59230, n71102, n3272, n3273, 
        n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
        n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
        n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3298, 
        n3301, n71100, n71094, n59229, n59228, n71088, n59227, 
        n59226, n24_adj_5856, n62, n71082, n59225, n59463, n59462, 
        n59461, n59224, n59460, n59459, n59458, n59457, n59456, 
        n59223, n59455, n59454, n71076, n59222, n59453, n59452, 
        n59451, n71070, n23094, n59450, n59221, n59449, n59448, 
        n59447, n59220, n25921, n59446, n59445, n9_adj_5857, n15_adj_5858, 
        n25_adj_5859, n32_adj_5860, n34, n39, n41, n79636, n59219, 
        n58895, n59218, n28274, n28272, n77205, n71066, n28240, 
        n59217, n59216, n28194, n58883, n59215, n45468, n28174, 
        n59214, n59213, n59212, n30398, n30395, n28130, n71058, 
        n59211, n28117, n4_adj_5861, n30392, n28099, n9_adj_5862, 
        n16_adj_5863, n20_adj_5864, n22_adj_5865, n25_adj_5866, n79624, 
        n33, n35, n37, n41_adj_5867, n79618, n79612, n21_adj_5868, 
        n79606, n37_adj_5869, n78778, n8_adj_5870, n10_adj_5871, n25_adj_5872, 
        n79600, n34_adj_5873, n36, n38, n79594, n38_adj_5874, n40, 
        n24_adj_5875, n79588, n79582, n28076, n2_adj_5876, n3_adj_5877, 
        n4_adj_5878, n5_adj_5879, n6_adj_5880, n7_adj_5881, n8_adj_5882, 
        n9_adj_5883, n10_adj_5884, n11_adj_5885, n12_adj_5886, n13_adj_5887, 
        n14_adj_5888, n15_adj_5889, n16_adj_5890, n17_adj_5891, n18_adj_5892, 
        n19_adj_5893, n20_adj_5894, n21_adj_5895, n22_adj_5896, n23_adj_5897, 
        n24_adj_5898, n25_adj_5899, n26_adj_5900, n27_adj_5901, n28_adj_5902, 
        n29_adj_5903, n30_adj_5904, n31_adj_5905, n32_adj_5906, n30388, 
        n59210, n59427, n59209, n59208, n59426, n59425, n59207, 
        n59424, n59206, n59423, n59422, n59421, n59205, n59204, 
        n59203, n71048, n58882, n44711, n77576, n44639, n71044, 
        n59420, n59419, n45370, n28051, n30382, n59418, n59417, 
        n71038, n78351, n60154, n60153, n59416, n59415, n60152, 
        n60151, n60150, n60149, n59414, n59413, n8_adj_5907, n59202, 
        n59412, n60148, n7_adj_5908, n59411, n59410, n67203, n25869, 
        n59201, n28027, n347_adj_5909, n59200, n59199, n59198, n59197, 
        n59196, n59195, n59194, n71026, n59193, n71020, n79576, 
        n27_adj_5910, n59192, n59191, n59190, n59189, n59188, n10_adj_5911, 
        n30_adj_5912, n59187, n59186, n25895, n59185, n78517, n71010, 
        n71004, n59184, n68474, n71002, n71000, n59183, n59182, 
        n59181, n58894, n59180, n58893, n59179, n58892, n58881, 
        n77575, n70984, n58999, n58998, n58997, n72383, n58996, 
        n58995, n58994, n58993, n79570, n68536, n137, n44574, 
        n70978, n51, n70976, n110, n70972, n79564, n78262, n70962, 
        n56, n38_adj_5913, n58992, n70954, n58991, n58990, n78215, 
        n70950, n75815, n6_adj_5914, n58989, n58988, n27243, n66576, 
        n70946, n58987, n58986, n27203, n27184, n58985, n70940, 
        n44675, n79243, n5_adj_5915, n67584, n79558, n67085, n27089, 
        n62972, n58984, n58983, n70934, n69738, n70932, n26999, 
        n78102, n79240, n79237, n78754, n70926, n70924, n70922, 
        n26760, n58982, n72380, n58981, n58980, n79234, n24_adj_5916, 
        n26619, n67135, n79552, n53108, n26875, n78020, n70906, 
        n70904, n12_adj_5917, n75797, n4_adj_5918, n6_adj_5919, n8_adj_5920, 
        n9_adj_5921, n11_adj_5922, n13_adj_5923, n14_adj_5924, n15_adj_5925, 
        n4_adj_5926, n6_adj_5927, n8_adj_5928, n9_adj_5929, n58979, 
        n25590, n70896, n38_adj_5930, n39_adj_5931, n40_adj_5932, 
        n41_adj_5933, n42, n43, n44, n45, n29756, n29755, n29752, 
        n79546, n26311, n79540, n6_adj_5934, n58978, n58977, n58891, 
        n58890, n67235, n62302, n78490, n77865, n29438, n70888, 
        n69558, n67238, n62277, n70882, n70878, n69065, n66744, 
        n66743, n66742, n66741, n66740, n66739, n66738, n66737, 
        n66736, n66735, n66734, n66733, n66732, n66731, n66730, 
        n66729, n66728, n66727, n66726, n66725, n29387, n66724, 
        n66723, n66722, n66721, n66720, n66719, n66718, n66717, 
        n66716, n66715, n66714, n66713, n29374, n70868, n66712, 
        n66711, n66710, n66867, n72039, n66872, n66866, n28730, 
        n66862, n28717, n28715, n28713, n66853, n28703, n28672, 
        n29155, n28664, n28662, n28656, n77694, n77693, n70860, 
        n58880, n77685, n44782, n10_adj_5935, n59386, n59385, n59384, 
        n8_adj_5936, n59383, n20468, n11851, n11849, n62510, n70854, 
        n6_adj_5937, n78095, n66709, n65800, n72378, n70848, n70846, 
        n20421, n59135, n59134, n30375, n30372, n30368, n30365, 
        n30362, n30355, n68441, n30349, n59133, n77684, n59132, 
        n58889, n70840, n59131, n29749, n45484, n79150, n79126, 
        n79120, n79114, n59382, n29746, n59130, n75727, n59129, 
        n59128, n68518, n25773, n29740, n25776, n59381, n78728, 
        n70830, n75719, n59127, n59126, n29734, n70824, n29731, 
        n68507, n59125, n77147, n25932, n59124, n59380, n70818, 
        n45520, n30267, n45496, n30264, n29727, n30261, n70812, 
        n30258, n30255, n30252, n30249, n70810, n59379, n70808, 
        n59378, n59377, n5_adj_5938, n70806, n36361, n25419, n59123, 
        n59376, n78463, n25421, n59375, n58879, n59374, n59373, 
        n59372, n59371, n59370, n59910, n59909, n59908, n59907, 
        n59906, n59905, n59904, n59903, n70784, n59902, n59901, 
        n59900, n59899, n59354, n59898, n59897, n59353, n59896, 
        n59895, n59894, n59893, n59892, n59891, n59890, n59889, 
        n59352, n59888, n59887, n59886, n59885, n59351, n59884, 
        n59350, n59883, n59882, n59881, n59880, n59879, n59349, 
        n59878, n70774, n59348, n59877, n70770, n59876, n59875, 
        n59874, n59873, n59872, n59871, n59870, n59869, n59868, 
        n59347, n70766, n59346, n59867, n59345, n59866, n59865, 
        n59344, n70760, n10_adj_5939, n59343, n59864, n14_adj_5940, 
        n59863, n59862, n59861, n59860, n59859, n13_adj_5941, n59858, 
        n59857, n59342, n59856, n59341, n59855, n59854, n59853, 
        n59852, n59851, n59850, n70754, n59849, n59848, n59847, 
        n59340, n59846, n59339, n59845, n59844, n59843, n59842, 
        n59841, n59840, n59839, n59838, n59837, n59836, n59835, 
        n76526, n59834, n59833, n70746, n59832, n59831, n79880, 
        n59830, n59829, n76520, n59828, n59827, n70740, n59826, 
        n59825, n59824, n59823, n59822, n58888, n59821, n59820, 
        n70734, n70732, n59819, n62281, n59818, n59817, n59816, 
        n59815, n59814, n59813, n79417, n59812, n59811, n59810, 
        n59809, n59808, n59318, n59317, n58887, n70718, n59807, 
        n59806, n59805, n59316, n59804, n59315, n59314, n70716, 
        n79414, n59803, n59802, n59801, n59800, n59313, n59799, 
        n59798, n59797, n59796, n59795, n59794, n59312, n59793, 
        n70714, n59792, n59311, n59310, n59309, n59791, n59790, 
        n59789, n59308, n59307, n59788, n58886, n59787, n59786, 
        n59785, n59784, n59783, n59782, n59306, n59781, n70712, 
        n59780, n59305, n59304, n58878, n59779, n70710, n13_adj_5942, 
        n15_adj_5943, n17_adj_5944, n25_adj_5945, n29_adj_5946, n31_adj_5947, 
        n35_adj_5948, n59778, n39_adj_5949, n49, n59777, n59776, 
        n59, n61, n59775, n59774, n59773, n59772, n59771, n59770, 
        n59769, n59768, n70704, n59767, n59766, n70702, n59765, 
        n59764, n59763, n8_adj_5950, n59762, n59761, n59760, n59759, 
        n59758, n70692, n78688, n59757, n59756, n12456, n70690, 
        n59755, n12450, n70688, n36147, n12462, n59754, n59753, 
        n58907, n66633, n12468, n72458, n58906, n59752, n12474, 
        n70686, n59751, n58586, n12480, n70684, n12486, n5_adj_5951, 
        n11_adj_5952, n58905, n70682, n12492, n70680, n77215, n59750, 
        n29369, n59749, n20467, n58877, n66708, n29367, n21158, 
        n29366, n58885, n21154, n59748, n59747, n66707, n66945, 
        n58904, n59746, n59745, n11914, n59744, n58903, n59743, 
        n59742, n59741, n58902, n10_adj_5953, n76403, n34689, n66706, 
        n59290, n59740, n70662, n59289, n25406, n59739, n59738, 
        n25771, n17_adj_5954, n61457, n59288, n20422, n61795, n76395, 
        n59737, n59736, n61432, n59287, n59286, n59735, n59734, 
        n26475, n75570, n59733, n59732, n61406, n59731, n77749, 
        n59730, n6_adj_5955, n61396, n78647, n77334, n59729, n68527, 
        n59728, n59727, n59726, n24045, n25912, n25885, n78151, 
        n59725, n75568, n59724, n59723, n59722, n59721, n59720, 
        n77333, n76359, n76324, n78612, n76303, n5_adj_5956, n69858, 
        n75564, n17_adj_5957, n25_adj_5958, n72168, n64972, n75562, 
        n24_adj_5959, n69393, n65060, n78096, n67629, n10_adj_5960, 
        n75317, n75301, n67243, n78930, n66790, n75275, n75272, 
        n75269, n67500, n67274, n67213, n34_adj_5961, n67361, n69463, 
        n75251, n75250, n70388, n75247, n75246, n69575, n69567, 
        n69502, n67425, n78917, n67578, n72460, n72459, n70372, 
        n66979, n69485, n67596, n67599, n70356, n4_adj_5962, n14_adj_5963, 
        n10_adj_5964, n78152, n70340, n66852, n70324, n6_adj_5965, 
        n75544, n4_adj_5966, n70308, n70292, n8_adj_5967, n7_adj_5968, 
        n68492, n70276, n75535, n68490, n65842, n66869, n69981, 
        n65866, n65870, n78580, n65874, n65878, n68571, n65884, 
        n65888, n65892, n65896, n65900, n78022, n65960, n68498, 
        n72094, n8_adj_5969, n65990, n65994, n65998, n75437, n75123, 
        n67259, n68433, n68431, n66142, n78373, n68582, n78265, 
        n75098, n75097, n78869, n78937, n75094, n75093, n68452, 
        n77519, n7_adj_5970;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n59771), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n28027), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i61349_4_lut (.I0(n15_adj_5777), .I1(n13_adj_5778), .I2(n11_adj_5779), 
            .I3(n76681), .O(n77205));
    defparam i61349_4_lut.LUT_INIT = 16'hfeff;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i61335_4_lut (.I0(n21_adj_5773), .I1(n19_adj_5774), .I2(n17_adj_5775), 
            .I3(n77205), .O(n77191));
    defparam i61335_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61969_4_lut (.I0(current[15]), .I1(n23_adj_5771), .I2(duty[12]), 
            .I3(n77191), .O(n77825));
    defparam i61969_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i60503_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n77825), .O(n76359));
    defparam i60503_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5785));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i61291_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5777), .O(n77147));
    defparam i61291_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5770));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i61893_3_lut (.I0(n4_adj_5785), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n77749));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61893_3_lut.LUT_INIT = 16'h8e8e;
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4126[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i60447_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n76324), .O(n76303));
    defparam i60447_4_lut.LUT_INIT = 16'h5adb;
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 LessThan_11_i35_rep_239_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n79880));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_239_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62164_3_lut (.I0(n30_adj_5770), .I1(n10_adj_5780), .I2(n77147), 
            .I3(GND_net), .O(n78020));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i62164_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .bit_ctr({Open_0, 
            Open_1, Open_2, bit_ctr[1:0]}), .\color_bit_N_502[1] (color_bit_N_502[1]), 
            .GND_net(GND_net), .neopxl_color({neopxl_color}), .timer({timer}), 
            .state({state}), .n29968(n29968), .t0({t0}), .n28194(n28194), 
            .\bit_ctr[3] (bit_ctr[3]), .\bit_ctr[4] (bit_ctr[4]), .VCC_net(VCC_net), 
            .n30584(n30584), .n30583(n30583), .n30582(n30582), .n30581(n30581), 
            .n30580(n30580), .n30579(n30579), .n30578(n30578), .n30577(n30577), 
            .n30576(n30576), .n30555(n30555), .n30479(n30479), .n65800(n65800), 
            .NEOPXL_c(NEOPXL_c), .n61457(n61457), .n61432(n61432), .\color_bit_N_502[2] (color_bit_N_502[2]), 
            .n44741(n44741), .n25406(n25406), .LED_c(LED_c), .n3165(n3165)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 i60547_4_lut (.I0(n77749), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n76403));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i60547_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i61837_3_lut (.I0(n6_adj_5784), .I1(duty[10]), .I2(n21_adj_5773), 
            .I3(GND_net), .O(n77693));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61837_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2039_5 (.CI(n59771), .I0(n3031), 
            .I1(VCC_net), .CO(n59772));
    SB_LUT4 i61838_3_lut (.I0(n77693), .I1(duty[11]), .I2(n23_adj_5771), 
            .I3(GND_net), .O(n77694));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61327_4_lut (.I0(current[15]), .I1(n23_adj_5771), .I2(duty[12]), 
            .I3(n75437), .O(n77183));
    defparam i61327_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5782), .I1(duty[9]), .I2(n19_adj_5774), 
            .I3(GND_net), .O(n16_adj_5776));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61684_3_lut (.I0(n77694), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n22_adj_5772));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61684_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61663_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n76359), .O(n77519));
    defparam i61663_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 encoder0_position_30__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n59770), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62359_4_lut (.I0(n76403), .I1(n78020), .I2(n79880), .I3(n76303), 
            .O(n78215));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i62359_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_30__I_0_add_2039_4 (.CI(n59770), .I0(n3032), 
            .I1(GND_net), .CO(n59771));
    SB_LUT4 encoder0_position_30__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n59769), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61679_3_lut (.I0(n22_adj_5772), .I1(n16_adj_5776), .I2(n77183), 
            .I3(GND_net), .O(n77535));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61679_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62409_4_lut (.I0(n77535), .I1(n78215), .I2(n79880), .I3(n77519), 
            .O(n78265));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i62409_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_30__I_0_add_2039_3 (.CI(n59769), .I0(n3033), 
            .I1(VCC_net), .CO(n59770));
    SB_LUT4 encoder0_position_30__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n59769));
    SB_LUT4 i62406_4_lut (.I0(n78265), .I1(duty[19]), .I2(current[15]), 
            .I3(duty[18]), .O(n78262));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i62406_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 encoder0_position_30__I_0_add_1972_29_lut (.I0(n78612), .I1(n2907), 
            .I2(VCC_net), .I3(n59768), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n59767), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_28 (.CI(n59767), .I0(n2908), 
            .I1(VCC_net), .CO(n59768));
    SB_LUT4 encoder0_position_30__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n59766), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(n78262), .I1(current[15]), .I2(duty[21]), .I3(duty[20]), 
            .O(n5_adj_5938));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n5_adj_5938), .I1(duty[23]), .I2(n51), .I3(duty[22]), 
            .O(n11851));
    defparam i7_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i15601_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n66852), .I3(GND_net), .O(n29815));   // verilog/coms.v(130[12] 305[6])
    defparam i15601_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15598_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n66852), .I3(GND_net), .O(n29812));   // verilog/coms.v(130[12] 305[6])
    defparam i15598_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16362_3_lut (.I0(t0[9]), .I1(timer[9]), .I2(n3165), .I3(GND_net), 
            .O(n30576));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16363_3_lut (.I0(t0[8]), .I1(timer[8]), .I2(n3165), .I3(GND_net), 
            .O(n30577));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16364_3_lut (.I0(t0[7]), .I1(timer[7]), .I2(n3165), .I3(GND_net), 
            .O(n30578));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16365_3_lut (.I0(t0[6]), .I1(timer[6]), .I2(n3165), .I3(GND_net), 
            .O(n30579));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16366_3_lut (.I0(t0[5]), .I1(timer[5]), .I2(n3165), .I3(GND_net), 
            .O(n30580));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16367_3_lut (.I0(t0[4]), .I1(timer[4]), .I2(n3165), .I3(GND_net), 
            .O(n30581));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16368_3_lut (.I0(t0[3]), .I1(timer[3]), .I2(n3165), .I3(GND_net), 
            .O(n30582));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16369_3_lut (.I0(t0[2]), .I1(timer[2]), .I2(n3165), .I3(GND_net), 
            .O(n30583));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16370_3_lut (.I0(t0[1]), .I1(timer[1]), .I2(n3165), .I3(GND_net), 
            .O(n30584));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16371_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n23025), .I3(GND_net), .O(n30585));   // verilog/coms.v(130[12] 305[6])
    defparam i16371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62760_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78616));
    defparam i62760_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5708));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_91[4]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15595_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n66852), .I3(GND_net), .O(n29809));   // verilog/coms.v(130[12] 305[6])
    defparam i15595_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16374_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n23025), .I3(GND_net), .O(n30588));   // verilog/coms.v(130[12] 305[6])
    defparam i16374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16375_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n23025), .I3(GND_net), .O(n30589));   // verilog/coms.v(130[12] 305[6])
    defparam i16375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15592_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n66852), .I3(GND_net), .O(n29806));   // verilog/coms.v(130[12] 305[6])
    defparam i15592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5709));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i59845_2_lut (.I0(n79), .I1(n8_adj_5834), .I2(GND_net), .I3(GND_net), 
            .O(n75247));   // verilog/coms.v(94[13:20])
    defparam i59845_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i27536_4_lut (.I0(n75247), .I1(n75246), .I2(rx_data[5]), .I3(\data_in_frame[17] [5]), 
            .O(n41669));   // verilog/coms.v(94[13:20])
    defparam i27536_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i27537_3_lut (.I0(n41669), .I1(\data_in_frame[17] [5]), .I2(reset), 
            .I3(GND_net), .O(n30593));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30473_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i30473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30598_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i30598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15789_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n23025), .I3(GND_net), .O(n30003));   // verilog/coms.v(130[12] 305[6])
    defparam i15789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15589_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n66852), .I3(GND_net), .O(n29803));   // verilog/coms.v(130[12] 305[6])
    defparam i15589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15794_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n30008));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15586_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n66852), .I3(GND_net), .O(n29800));   // verilog/coms.v(130[12] 305[6])
    defparam i15586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i63032_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78888));
    defparam i63032_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16389_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n23025), .I3(GND_net), .O(n30603));   // verilog/coms.v(130[12] 305[6])
    defparam i16389_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1972_27 (.CI(n59766), .I0(n2909), 
            .I1(VCC_net), .CO(n59767));
    SB_LUT4 i589_2_lut (.I0(n1319), .I1(n44574), .I2(GND_net), .I3(GND_net), 
            .O(n2821));   // verilog/TinyFPGA_B.v(384[18] 386[12])
    defparam i589_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16053_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n28730), 
            .I3(GND_net), .O(n30267));   // verilog/coms.v(130[12] 305[6])
    defparam i16053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n59765), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15583_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n66852), .I3(GND_net), .O(n29797));   // verilog/coms.v(130[12] 305[6])
    defparam i15583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16817_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n31031));   // verilog/coms.v(130[12] 305[6])
    defparam i16817_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i63002_2_lut (.I0(n23188), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i63002_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i15580_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n66852), .I3(GND_net), .O(n29794));   // verilog/coms.v(130[12] 305[6])
    defparam i15580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i56321_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n72168));
    defparam i56321_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i63205_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6903), .I2(n72168), 
            .I3(n25_adj_5958), .O(n17_adj_5957));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i63205_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i15799_3_lut (.I0(a_prev_adj_5796), .I1(a_new_adj_6010[1]), 
            .I2(debounce_cnt_N_3833_adj_5798), .I3(GND_net), .O(n30013));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15799_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16874_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n31088));   // verilog/coms.v(130[12] 305[6])
    defparam i16874_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1972_26 (.CI(n59765), .I0(n2910), 
            .I1(VCC_net), .CO(n59766));
    SB_LUT4 i16402_3_lut (.I0(\data_in_frame[17] [6]), .I1(rx_data[6]), 
            .I2(n28715), .I3(GND_net), .O(n30616));   // verilog/coms.v(130[12] 305[6])
    defparam i16402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16405_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n23025), .I3(GND_net), .O(n30619));   // verilog/coms.v(130[12] 305[6])
    defparam i16405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16050_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n28730), 
            .I3(GND_net), .O(n30264));   // verilog/coms.v(130[12] 305[6])
    defparam i16050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n59764), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15893_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[1]), .I2(n5_adj_5791), 
            .I3(n25895), .O(n30107));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15893_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16047_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n28730), 
            .I3(GND_net), .O(n30261));   // verilog/coms.v(130[12] 305[6])
    defparam i16047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16044_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n28730), 
            .I3(GND_net), .O(n30258));   // verilog/coms.v(130[12] 305[6])
    defparam i16044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15549_3_lut (.I0(\data_in_frame[19] [7]), .I1(rx_data[7]), 
            .I2(n69075), .I3(GND_net), .O(n29763));   // verilog/coms.v(130[12] 305[6])
    defparam i15549_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16041_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n28730), 
            .I3(GND_net), .O(n30255));   // verilog/coms.v(130[12] 305[6])
    defparam i16041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15894_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[2]), .I2(n5_adj_5817), 
            .I3(n25895), .O(n30108));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15894_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16038_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n28730), 
            .I3(GND_net), .O(n30252));   // verilog/coms.v(130[12] 305[6])
    defparam i16038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15545_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n69075), .I3(GND_net), .O(n29759));   // verilog/coms.v(130[12] 305[6])
    defparam i15545_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [2]), 
            .I2(\data_out_frame[20] [1]), .I3(GND_net), .O(n67085));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY encoder0_position_30__I_0_add_1972_25 (.CI(n59764), .I0(n2911), 
            .I1(VCC_net), .CO(n59765));
    SB_LUT4 i16035_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n28730), 
            .I3(GND_net), .O(n30249));   // verilog/coms.v(130[12] 305[6])
    defparam i16035_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n59763), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16418_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n23025), .I3(GND_net), .O(n30632));   // verilog/coms.v(130[12] 305[6])
    defparam i16418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1972_24 (.CI(n59763), .I0(n2912), 
            .I1(VCC_net), .CO(n59764));
    SB_LUT4 i15895_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[3]), .I2(n44711), 
            .I3(n25895), .O(n30109));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15895_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5710));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15896_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[4]), .I2(n5_adj_5807), 
            .I3(n25885), .O(n30110));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15896_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15897_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[5]), .I2(n5_adj_5791), 
            .I3(n25885), .O(n30111));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15897_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15898_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[6]), .I2(n5_adj_5817), 
            .I3(n25885), .O(n30112));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15898_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n59762), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15899_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[7]), .I2(n44711), 
            .I3(n25885), .O(n30113));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15899_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15900_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[8]), .I2(n5_adj_5807), 
            .I3(n25869), .O(n30114));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15900_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_30__I_0_add_1972_23 (.CI(n59762), .I0(n2913), 
            .I1(VCC_net), .CO(n59763));
    SB_LUT4 i15901_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[9]), .I2(n5_adj_5791), 
            .I3(n25869), .O(n30115));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15901_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_3812_i6_3_lut (.I0(encoder0_position[5]), .I1(n27), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15902_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[10]), .I2(n5_adj_5817), 
            .I3(n25869), .O(n30116));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15902_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15903_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[11]), .I2(n44711), 
            .I3(n25869), .O(n30117));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15903_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n59761), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_22 (.CI(n59761), .I0(n2914), 
            .I1(VCC_net), .CO(n59762));
    SB_LUT4 i20486_3_lut (.I0(n28730), .I1(rx_data[0]), .I2(\data_in_frame[9] [0]), 
            .I3(GND_net), .O(n30666));   // verilog/coms.v(94[13:20])
    defparam i20486_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i16453_3_lut (.I0(current[11]), .I1(data_adj_6031[11]), .I2(n28099), 
            .I3(GND_net), .O(n30667));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15904_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[12]), .I2(n5_adj_5807), 
            .I3(n25912), .O(n30118));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15904_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16454_3_lut (.I0(current[10]), .I1(data_adj_6031[10]), .I2(n28099), 
            .I3(GND_net), .O(n30668));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16455_3_lut (.I0(current[9]), .I1(data_adj_6031[9]), .I2(n28099), 
            .I3(GND_net), .O(n30669));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16456_3_lut (.I0(current[8]), .I1(data_adj_6031[8]), .I2(n28099), 
            .I3(GND_net), .O(n30670));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16457_3_lut (.I0(current[7]), .I1(data_adj_6031[7]), .I2(n28099), 
            .I3(GND_net), .O(n30671));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16458_3_lut (.I0(current[6]), .I1(data_adj_6031[6]), .I2(n28099), 
            .I3(GND_net), .O(n30672));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16459_3_lut (.I0(current[5]), .I1(data_adj_6031[5]), .I2(n28099), 
            .I3(GND_net), .O(n30673));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63586 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[17] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[0]), .O(n79414));
    defparam byte_transmit_counter_1__bdd_4_lut_63586.LUT_INIT = 16'he4aa;
    SB_LUT4 i16460_3_lut (.I0(current[4]), .I1(data_adj_6031[4]), .I2(n28099), 
            .I3(GND_net), .O(n30674));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16461_3_lut (.I0(current[3]), .I1(data_adj_6031[3]), .I2(n28099), 
            .I3(GND_net), .O(n30675));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16462_3_lut (.I0(current[2]), .I1(data_adj_6031[2]), .I2(n28099), 
            .I3(GND_net), .O(n30676));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16463_3_lut (.I0(current[1]), .I1(data_adj_6031[1]), .I2(n28099), 
            .I3(GND_net), .O(n30677));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n59760), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16464_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n23025), .I3(GND_net), .O(n30678));   // verilog/coms.v(130[12] 305[6])
    defparam i16464_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1972_21 (.CI(n59760), .I0(n2915), 
            .I1(VCC_net), .CO(n59761));
    SB_LUT4 encoder0_position_30__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n59759), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_20 (.CI(n59759), .I0(n2916), 
            .I1(VCC_net), .CO(n59760));
    SB_LUT4 encoder0_position_30__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n59758), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_19 (.CI(n59758), .I0(n2917), 
            .I1(VCC_net), .CO(n59759));
    SB_LUT4 encoder0_position_30__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n59757), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_18 (.CI(n59757), .I0(n2918), 
            .I1(VCC_net), .CO(n59758));
    SB_LUT4 encoder0_position_30__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n59756), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_17 (.CI(n59756), .I0(n2919), 
            .I1(VCC_net), .CO(n59757));
    SB_LUT4 encoder0_position_30__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n59755), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_16 (.CI(n59755), .I0(n2920), 
            .I1(VCC_net), .CO(n59756));
    SB_LUT4 i15542_3_lut (.I0(\data_in_frame[19] [5]), .I1(rx_data[5]), 
            .I2(n69075), .I3(GND_net), .O(n29756));   // verilog/coms.v(130[12] 305[6])
    defparam i15542_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15905_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[15]), .I2(n44711), 
            .I3(n25912), .O(n30119));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15905_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n59754), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_15 (.CI(n59754), .I0(n2921), 
            .I1(VCC_net), .CO(n59755));
    SB_LUT4 encoder0_position_30__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n59753), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_14 (.CI(n59753), .I0(n2922), 
            .I1(VCC_net), .CO(n59754));
    SB_LUT4 encoder0_position_30__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n59752), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_30__I_0_add_1972_13 (.CI(n59752), .I0(n2923), 
            .I1(VCC_net), .CO(n59753));
    SB_LUT4 encoder0_position_30__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n59751), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_12 (.CI(n59751), .I0(n2924), 
            .I1(VCC_net), .CO(n59752));
    SB_LUT4 n79414_bdd_4_lut (.I0(n79414), .I1(\data_out_frame[18] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[0]), 
            .O(n79417));
    defparam n79414_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n59750), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15909_3_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), .I2(n66867), 
            .I3(GND_net), .O(n30123));   // verilog/coms.v(130[12] 305[6])
    defparam i15909_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1972_11 (.CI(n59750), .I0(n2925), 
            .I1(VCC_net), .CO(n59751));
    SB_LUT4 encoder0_position_30__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15912_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n66867), 
            .I3(GND_net), .O(n30126));   // verilog/coms.v(130[12] 305[6])
    defparam i15912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n59749), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_10 (.CI(n59749), .I0(n2926), 
            .I1(VCC_net), .CO(n59750));
    SB_LUT4 encoder0_position_30__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n59748), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i15915_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n66867), 
            .I3(GND_net), .O(n30129));   // verilog/coms.v(130[12] 305[6])
    defparam i15915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1773_3_lut (.I0(n2610), .I1(n2677), 
            .I2(n2643), .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51829_3_lut (.I0(n3), .I1(n7757), .I2(n67628), .I3(GND_net), 
            .O(n67629));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51829_3_lut.LUT_INIT = 16'hcaca;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_30__I_0_add_1972_9 (.CI(n59748), .I0(n2927), 
            .I1(VCC_net), .CO(n59749));
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i16476_3_lut (.I0(baudrate[23]), .I1(data_adj_6024[7]), .I2(n28272), 
            .I3(GND_net), .O(n30690));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16477_3_lut (.I0(baudrate[22]), .I1(data_adj_6024[6]), .I2(n28272), 
            .I3(GND_net), .O(n30691));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n59747), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16478_3_lut (.I0(baudrate[21]), .I1(data_adj_6024[5]), .I2(n28272), 
            .I3(GND_net), .O(n30692));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16478_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1972_8 (.CI(n59747), .I0(n2928), 
            .I1(VCC_net), .CO(n59748));
    SB_LUT4 i16479_3_lut (.I0(baudrate[20]), .I1(data_adj_6024[4]), .I2(n28272), 
            .I3(GND_net), .O(n30693));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n59746), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_7 (.CI(n59746), .I0(n2929), 
            .I1(GND_net), .CO(n59747));
    SB_LUT4 encoder0_position_30__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n59745), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_6 (.CI(n59745), .I0(n2930), 
            .I1(GND_net), .CO(n59746));
    SB_LUT4 encoder0_position_30__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n59744), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_5 (.CI(n59744), .I0(n2931), 
            .I1(VCC_net), .CO(n59745));
    SB_LUT4 i16480_3_lut (.I0(baudrate[19]), .I1(data_adj_6024[3]), .I2(n28272), 
            .I3(GND_net), .O(n30694));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16481_3_lut (.I0(baudrate[18]), .I1(data_adj_6024[2]), .I2(n28272), 
            .I3(GND_net), .O(n30695));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16482_3_lut (.I0(baudrate[17]), .I1(data_adj_6024[1]), .I2(n28272), 
            .I3(GND_net), .O(n30696));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16482_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i16483_3_lut (.I0(baudrate[16]), .I1(data_adj_6024[0]), .I2(n28272), 
            .I3(GND_net), .O(n30697));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16483_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n59743), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_4 (.CI(n59743), .I0(n2932), 
            .I1(GND_net), .CO(n59744));
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n59742), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1972_3 (.CI(n59742), .I0(n2933), 
            .I1(VCC_net), .CO(n59743));
    SB_LUT4 encoder0_position_30__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n59742));
    SB_LUT4 encoder0_position_30__I_0_add_1905_28_lut (.I0(GND_net), .I1(n2808), 
            .I2(VCC_net), .I3(n59741), .O(n2875)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n59740), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_27 (.CI(n59740), .I0(n2809), 
            .I1(VCC_net), .CO(n59741));
    SB_LUT4 encoder0_position_30__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n59739), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_26 (.CI(n59739), .I0(n2810), 
            .I1(VCC_net), .CO(n59740));
    SB_LUT4 i15918_3_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), .I2(n66867), 
            .I3(GND_net), .O(n30132));   // verilog/coms.v(130[12] 305[6])
    defparam i15918_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n59738), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_25 (.CI(n59738), .I0(n2811), 
            .I1(VCC_net), .CO(n59739));
    SB_LUT4 encoder0_position_30__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n59737), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_24 (.CI(n59737), .I0(n2812), 
            .I1(VCC_net), .CO(n59738));
    SB_LUT4 i51830_3_lut (.I0(encoder0_position[29]), .I1(n67629), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n59736), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1905_23 (.CI(n59736), .I0(n2813), 
            .I1(VCC_net), .CO(n59737));
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n59735), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i56603_3_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n72459));
    defparam i56603_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1905_22 (.CI(n59735), .I0(n2814), 
            .I1(VCC_net), .CO(n59736));
    SB_LUT4 encoder0_position_30__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n59734), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_21 (.CI(n59734), .I0(n2815), 
            .I1(VCC_net), .CO(n59735));
    SB_LUT4 encoder0_position_30__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n59733), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i56602_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[6] [7]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n72458));
    defparam i56602_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1905_20 (.CI(n59733), .I0(n2816), 
            .I1(VCC_net), .CO(n59734));
    SB_LUT4 i56604_4_lut (.I0(n72459), .I1(n28392), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n72460));
    defparam i56604_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 encoder0_position_30__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n59732), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_19 (.CI(n59732), .I0(n2817), 
            .I1(VCC_net), .CO(n59733));
    SB_LUT4 encoder0_position_30__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n59731), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_18 (.CI(n59731), .I0(n2818), 
            .I1(VCC_net), .CO(n59732));
    SB_CARRY add_151_14 (.CI(n58888), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n58889));
    SB_LUT4 encoder0_position_30__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n59730), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_17 (.CI(n59730), .I0(n2819), 
            .I1(VCC_net), .CO(n59731));
    SB_LUT4 encoder0_position_30__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n59729), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_16 (.CI(n59729), .I0(n2820), 
            .I1(VCC_net), .CO(n59730));
    SB_LUT4 encoder0_position_30__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821_adj_5854), 
            .I2(VCC_net), .I3(n59728), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_15 (.CI(n59728), .I0(n2821_adj_5854), 
            .I1(VCC_net), .CO(n59729));
    SB_LUT4 encoder0_position_30__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n59727), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_14 (.CI(n59727), .I0(n2822), 
            .I1(VCC_net), .CO(n59728));
    SB_LUT4 i16493_3_lut (.I0(baudrate[7]), .I1(data_adj_6024[7]), .I2(n28274), 
            .I3(GND_net), .O(n30707));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n59726), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16494_3_lut (.I0(baudrate[6]), .I1(data_adj_6024[6]), .I2(n28274), 
            .I3(GND_net), .O(n30708));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16495_3_lut (.I0(baudrate[5]), .I1(data_adj_6024[5]), .I2(n28274), 
            .I3(GND_net), .O(n30709));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16496_3_lut (.I0(baudrate[4]), .I1(data_adj_6024[4]), .I2(n28274), 
            .I3(GND_net), .O(n30710));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16496_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1905_13 (.CI(n59726), .I0(n2823), 
            .I1(VCC_net), .CO(n59727));
    SB_LUT4 encoder0_position_30__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n59725), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_12 (.CI(n59725), .I0(n2824), 
            .I1(VCC_net), .CO(n59726));
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n59724), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i16497_3_lut (.I0(baudrate[3]), .I1(data_adj_6024[3]), .I2(n28274), 
            .I3(GND_net), .O(n30711));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16497_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1905_11 (.CI(n59724), .I0(n2825), 
            .I1(VCC_net), .CO(n59725));
    SB_LUT4 i16498_3_lut (.I0(baudrate[2]), .I1(data_adj_6024[2]), .I2(n28274), 
            .I3(GND_net), .O(n30712));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16499_3_lut (.I0(baudrate[1]), .I1(data_adj_6024[1]), .I2(n28274), 
            .I3(GND_net), .O(n30713));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n59723), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_10 (.CI(n59723), .I0(n2826), 
            .I1(VCC_net), .CO(n59724));
    SB_LUT4 encoder0_position_30__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n59722), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_9 (.CI(n59722), .I0(n2827), 
            .I1(VCC_net), .CO(n59723));
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28130), 
            .D(n1238), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_1034_15_lut (.I0(n78848), .I1(n1521), 
            .I2(VCC_net), .I3(n59259), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15921_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n66867), 
            .I3(GND_net), .O(n30135));   // verilog/coms.v(130[12] 305[6])
    defparam i15921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15924_3_lut (.I0(\data_in_frame[4] [5]), .I1(rx_data[5]), .I2(n66867), 
            .I3(GND_net), .O(n30138));   // verilog/coms.v(130[12] 305[6])
    defparam i15924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15927_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n66867), 
            .I3(GND_net), .O(n30141));   // verilog/coms.v(130[12] 305[6])
    defparam i15927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n59721), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_8 (.CI(n59721), .I0(n2828), 
            .I1(VCC_net), .CO(n59722));
    SB_LUT4 encoder0_position_30__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n59720), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_7 (.CI(n59720), .I0(n2829), 
            .I1(GND_net), .CO(n59721));
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n58879), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n59719), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5805), .I3(n59053), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(n62281), .I1(n61406), .I2(n26619), .I3(n6_adj_5743), 
            .O(n25419));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_30__I_0_add_1905_6 (.CI(n59719), .I0(n2830), 
            .I1(GND_net), .CO(n59720));
    SB_LUT4 i16500_3_lut (.I0(baudrate[0]), .I1(data_adj_6024[0]), .I2(n28274), 
            .I3(GND_net), .O(n30714));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15931_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n66867), 
            .I3(GND_net), .O(n30145));   // verilog/coms.v(130[12] 305[6])
    defparam i15931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n59718), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_5 (.CI(n59718), .I0(n2831), 
            .I1(VCC_net), .CO(n59719));
    SB_LUT4 encoder0_position_30__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5711));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n59258), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n58887), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_14 (.CI(n59258), .I0(n1522), 
            .I1(VCC_net), .CO(n59259));
    SB_LUT4 encoder0_position_30__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n59257), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5804), .I3(n59052), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5800));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n59052), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5804), .CO(n59053));
    SB_CARRY encoder0_position_30__I_0_add_1034_13 (.CI(n59257), .I0(n1523), 
            .I1(VCC_net), .CO(n59258));
    SB_LUT4 encoder0_position_30__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n59717), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_91[5]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1905_4 (.CI(n59717), .I0(n2832), 
            .I1(GND_net), .CO(n59718));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5803), .I3(n59051), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_13 (.CI(n58887), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n58888));
    SB_LUT4 mux_243_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_91[6]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n59716), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n59256), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_3 (.CI(n59716), .I0(n2833), 
            .I1(VCC_net), .CO(n59717));
    SB_LUT4 encoder0_position_30__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5801));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5802));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n59051), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5803), .CO(n59052));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5818));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_12 (.CI(n59256), .I0(n1524), 
            .I1(VCC_net), .CO(n59257));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5819));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5822), .I3(n59050), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n59716));
    SB_LUT4 encoder0_position_30__I_0_add_1838_27_lut (.I0(GND_net), .I1(n2709), 
            .I2(VCC_net), .I3(n59715), .O(n2776)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n59714), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15934_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n66866), 
            .I3(GND_net), .O(n30148));   // verilog/coms.v(130[12] 305[6])
    defparam i15934_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_26 (.CI(n59714), .I0(n2710), 
            .I1(VCC_net), .CO(n59715));
    SB_LUT4 encoder0_position_30__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n59713), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n59255), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_11 (.CI(n59255), .I0(n1525), 
            .I1(VCC_net), .CO(n59256));
    SB_CARRY encoder0_position_30__I_0_add_1838_25 (.CI(n59713), .I0(n2711), 
            .I1(VCC_net), .CO(n59714));
    SB_LUT4 encoder0_position_30__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n59712), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n59050), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5822), .CO(n59051));
    SB_CARRY encoder0_position_30__I_0_add_1838_24 (.CI(n59712), .I0(n2712), 
            .I1(VCC_net), .CO(n59713));
    SB_LUT4 encoder0_position_30__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n59711), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5821), .I3(n59049), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_23 (.CI(n59711), .I0(n2713), 
            .I1(VCC_net), .CO(n59712));
    SB_LUT4 encoder0_position_30__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n59254), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_10 (.CI(n59254), .I0(n1526), 
            .I1(VCC_net), .CO(n59255));
    SB_LUT4 encoder0_position_30__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n59710), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_22 (.CI(n59710), .I0(n2714), 
            .I1(VCC_net), .CO(n59711));
    SB_LUT4 encoder0_position_30__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n59709), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_21 (.CI(n59709), .I0(n2715), 
            .I1(VCC_net), .CO(n59710));
    SB_LUT4 encoder0_position_30__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n59708), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n59253), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15538_3_lut (.I0(\data_in_frame[19] [4]), .I1(rx_data[4]), 
            .I2(n69075), .I3(GND_net), .O(n29752));   // verilog/coms.v(130[12] 305[6])
    defparam i15538_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1034_9 (.CI(n59253), .I0(n1527), 
            .I1(VCC_net), .CO(n59254));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n59049), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5821), .CO(n59050));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5820), .I3(n59048), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_20 (.CI(n59708), .I0(n2716), 
            .I1(VCC_net), .CO(n59709));
    SB_LUT4 encoder0_position_30__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n59707), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n59048), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5820), .CO(n59049));
    SB_CARRY encoder0_position_30__I_0_add_1838_19 (.CI(n59707), .I0(n2717), 
            .I1(VCC_net), .CO(n59708));
    SB_LUT4 encoder0_position_30__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n59706), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_18 (.CI(n59706), .I0(n2718), 
            .I1(VCC_net), .CO(n59707));
    SB_LUT4 encoder0_position_30__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225_adj_5837));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15535_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n69075), .I3(GND_net), .O(n29749));   // verilog/coms.v(130[12] 305[6])
    defparam i15535_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28130), 
            .D(n1237), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i15937_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n66866), 
            .I3(GND_net), .O(n30151));   // verilog/coms.v(130[12] 305[6])
    defparam i15937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15940_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n66866), 
            .I3(GND_net), .O(n30154));   // verilog/coms.v(130[12] 305[6])
    defparam i15940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n59705), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i836_3_lut (.I0(n1225_adj_5837), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_17 (.CI(n59705), .I0(n2719), 
            .I1(VCC_net), .CO(n59706));
    SB_LUT4 encoder0_position_30__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n59704), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_16 (.CI(n59704), .I0(n2720), 
            .I1(VCC_net), .CO(n59705));
    SB_LUT4 i15943_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n66866), 
            .I3(GND_net), .O(n30157));   // verilog/coms.v(130[12] 305[6])
    defparam i15943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15946_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n66866), 
            .I3(GND_net), .O(n30160));   // verilog/coms.v(130[12] 305[6])
    defparam i15946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n59703), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_15 (.CI(n59703), .I0(n2721), 
            .I1(VCC_net), .CO(n59704));
    SB_LUT4 encoder0_position_30__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n59702), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_14 (.CI(n59702), .I0(n2722), 
            .I1(VCC_net), .CO(n59703));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5819), .I3(n59047), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n59701), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_13 (.CI(n59701), .I0(n2723), 
            .I1(VCC_net), .CO(n59702));
    SB_LUT4 encoder0_position_30__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n59252), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n59700), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5820));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1034_8 (.CI(n59252), .I0(n1528), 
            .I1(VCC_net), .CO(n59253));
    SB_CARRY encoder0_position_30__I_0_add_1838_12 (.CI(n59700), .I0(n2724), 
            .I1(VCC_net), .CO(n59701));
    SB_LUT4 encoder0_position_30__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n59699), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n59047), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5819), .CO(n59048));
    SB_CARRY encoder0_position_30__I_0_add_1838_11 (.CI(n59699), .I0(n2725), 
            .I1(VCC_net), .CO(n59700));
    SB_LUT4 encoder0_position_30__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n59698), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_10 (.CI(n59698), .I0(n2726), 
            .I1(VCC_net), .CO(n59699));
    SB_LUT4 encoder0_position_30__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n59697), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_9 (.CI(n59697), .I0(n2727), 
            .I1(VCC_net), .CO(n59698));
    SB_LUT4 encoder0_position_30__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n59251), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n59696), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_8 (.CI(n59696), .I0(n2728), 
            .I1(VCC_net), .CO(n59697));
    SB_CARRY encoder0_position_30__I_0_add_1034_7 (.CI(n59251), .I0(n1529), 
            .I1(GND_net), .CO(n59252));
    SB_LUT4 encoder0_position_30__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n59695), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n59250), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_7 (.CI(n59695), .I0(n2729), 
            .I1(GND_net), .CO(n59696));
    SB_CARRY encoder0_position_30__I_0_add_1034_6 (.CI(n59250), .I0(n1530), 
            .I1(GND_net), .CO(n59251));
    SB_LUT4 encoder0_position_30__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n59249), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n59694), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5818), .I3(n59046), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n59046), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5818), .CO(n59047));
    SB_CARRY encoder0_position_30__I_0_add_1838_6 (.CI(n59694), .I0(n2730), 
            .I1(GND_net), .CO(n59695));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5802), .I3(n59045), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n59693), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16513_3_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(n28715), .I3(GND_net), .O(n30727));   // verilog/coms.v(130[12] 305[6])
    defparam i16513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15532_3_lut (.I0(\data_in_frame[19] [2]), .I1(rx_data[2]), 
            .I2(n69075), .I3(GND_net), .O(n29746));   // verilog/coms.v(130[12] 305[6])
    defparam i15532_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5821));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1838_5 (.CI(n59693), .I0(n2731), 
            .I1(VCC_net), .CO(n59694));
    SB_LUT4 encoder0_position_30__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n59692), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_4 (.CI(n59692), .I0(n2732), 
            .I1(GND_net), .CO(n59693));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n59045), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5802), .CO(n59046));
    SB_LUT4 encoder0_position_30__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n59691), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5801), .I3(n59044), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_3 (.CI(n59691), .I0(n2733), 
            .I1(VCC_net), .CO(n59692));
    SB_LUT4 i15949_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n66866), 
            .I3(GND_net), .O(n30163));   // verilog/coms.v(130[12] 305[6])
    defparam i15949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n59691));
    SB_LUT4 i16520_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n23025), .I3(GND_net), .O(n30734));   // verilog/coms.v(130[12] 305[6])
    defparam i16520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n58886), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_26_lut (.I0(GND_net), .I1(n2610), 
            .I2(VCC_net), .I3(n59690), .O(n2677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n59044), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5801), .CO(n59045));
    SB_LUT4 encoder0_position_30__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n59689), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5800), .I3(n59043), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_25 (.CI(n59689), .I0(n2611), 
            .I1(VCC_net), .CO(n59690));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5822));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15526_3_lut (.I0(\data_in_frame[19] [0]), .I1(rx_data[0]), 
            .I2(n69075), .I3(GND_net), .O(n29740));   // verilog/coms.v(130[12] 305[6])
    defparam i15526_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n59688), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_24 (.CI(n59688), .I0(n2612), 
            .I1(VCC_net), .CO(n59689));
    SB_LUT4 encoder0_position_30__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n59687), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[18] [7]), .I1(n28656), .I2(n28713), 
            .I3(rx_data[7]), .O(n65884));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i16526_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n28713), .I3(GND_net), .O(n30740));   // verilog/coms.v(130[12] 305[6])
    defparam i16526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15520_3_lut (.I0(\data_in_frame[18] [6]), .I1(rx_data[6]), 
            .I2(n28713), .I3(GND_net), .O(n29734));   // verilog/coms.v(130[12] 305[6])
    defparam i15520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_2_lut (.I0(n291), .I1(n239), .I2(GND_net), .I3(GND_net), 
            .O(n37_adj_5869));
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1771_23 (.CI(n59687), .I0(n2613), 
            .I1(VCC_net), .CO(n59688));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n59043), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5800), .CO(n59044));
    SB_LUT4 i15517_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n28713), .I3(GND_net), .O(n29731));   // verilog/coms.v(130[12] 305[6])
    defparam i15517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1819 (.I0(\data_in_frame[18] [4]), .I1(n28656), 
            .I2(n28713), .I3(rx_data[4]), .O(n65888));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1819.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n59686), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_22 (.CI(n59686), .I0(n2614), 
            .I1(VCC_net), .CO(n59687));
    SB_LUT4 encoder0_position_30__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n59685), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_5 (.CI(n59249), .I0(n1531), 
            .I1(VCC_net), .CO(n59250));
    SB_CARRY encoder0_position_30__I_0_add_1771_21 (.CI(n59685), .I0(n2615), 
            .I1(VCC_net), .CO(n59686));
    SB_LUT4 encoder0_position_30__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n59248), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_4 (.CI(n59248), .I0(n1532), 
            .I1(GND_net), .CO(n59249));
    SB_LUT4 i16534_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n21154), .I3(n4_adj_5962), .O(n30748));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i16534_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 encoder0_position_30__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n59684), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5711), .I3(n59042), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59810_3_lut (.I0(state_7__N_4110[0]), .I1(n11_adj_5789), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n75317));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i59810_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i16_4_lut (.I0(state_adj_6057[0]), .I1(n75317), .I2(n6707), 
            .I3(n44639), .O(n8_adj_5969));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 i16537_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[0]), 
            .I2(n10_adj_5953), .I3(n25890), .O(n30751));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16537_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1771_20 (.CI(n59684), .I0(n2616), 
            .I1(VCC_net), .CO(n59685));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n59042), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5711), .CO(n59043));
    SB_LUT4 i12_4_lut_adj_1820 (.I0(\data_in_frame[18] [3]), .I1(n28656), 
            .I2(n28713), .I3(rx_data[3]), .O(n65892));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1820.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5803));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n59683), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16544_3_lut (.I0(n67800), .I1(r_Bit_Index[0]), .I2(n28240), 
            .I3(GND_net), .O(n30758));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16544_3_lut.LUT_INIT = 16'h1414;
    SB_CARRY encoder0_position_30__I_0_add_1771_19 (.CI(n59683), .I0(n2617), 
            .I1(VCC_net), .CO(n59684));
    SB_LUT4 i16548_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n70292), 
            .I3(n27_adj_5855), .O(n30762));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16548_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n59682), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n59247), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_3 (.CI(n59247), .I0(n1533), 
            .I1(VCC_net), .CO(n59248));
    SB_CARRY encoder0_position_30__I_0_add_1771_18 (.CI(n59682), .I0(n2618), 
            .I1(VCC_net), .CO(n59683));
    SB_LUT4 encoder0_position_30__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n59681), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14), .I3(n59041), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_17 (.CI(n59681), .I0(n2619), 
            .I1(VCC_net), .CO(n59682));
    SB_LUT4 encoder0_position_30__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n59680), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_16 (.CI(n59680), .I0(n2620), 
            .I1(VCC_net), .CO(n59681));
    SB_LUT4 encoder0_position_30__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n59679), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_15 (.CI(n59679), .I0(n2621), 
            .I1(VCC_net), .CO(n59680));
    SB_LUT4 encoder0_position_30__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16553_4_lut (.I0(CS_MISO_c), .I1(data_adj_6031[0]), .I2(n11_adj_5792), 
            .I3(state_7__N_4319), .O(n30767));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16553_4_lut.LUT_INIT = 16'hccca;
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n59678), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_14 (.CI(n59678), .I0(n2622), 
            .I1(VCC_net), .CO(n59679));
    SB_LUT4 encoder0_position_30__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n59677), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1821 (.I0(\data_in_frame[18] [2]), .I1(n28656), 
            .I2(n28713), .I3(rx_data[2]), .O(n65896));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1821.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_30__I_0_add_1771_13 (.CI(n59677), .I0(n2623), 
            .I1(VCC_net), .CO(n59678));
    SB_LUT4 encoder0_position_30__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n59676), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28130), 
            .D(n1236), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28130), 
            .D(n1235), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28130), 
            .D(n1234), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_CARRY encoder0_position_30__I_0_add_1771_12 (.CI(n59676), .I0(n2624), 
            .I1(VCC_net), .CO(n59677));
    SB_LUT4 encoder0_position_30__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n59675), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28130), 
            .D(n1233), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i7_2_lut (.I0(PWMLimit[20]), .I1(setpoint[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5867));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_2_lut (.I0(PWMLimit[18]), .I1(setpoint[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13_2_lut (.I0(PWMLimit[4]), .I1(setpoint[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5862));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(n8_adj_5835), .I1(n41637), .I2(GND_net), .I3(GND_net), 
            .O(n28656));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28130), 
            .D(n1232), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28130), 
            .D(n1231), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28130), 
            .D(n1230), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1822 (.I0(\data_in_frame[18] [1]), .I1(n28656), 
            .I2(n28713), .I3(rx_data[1]), .O(n65900));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1822.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_30__I_0_add_1771_11 (.CI(n59675), .I0(n2625), 
            .I1(VCC_net), .CO(n59676));
    SB_LUT4 i16565_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n23094), .I3(GND_net), .O(n30779));   // verilog/coms.v(130[12] 305[6])
    defparam i16565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16567_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n23094), .I3(GND_net), .O(n30781));   // verilog/coms.v(130[12] 305[6])
    defparam i16567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59651_4_lut (.I0(data_ready), .I1(n6903), .I2(n24_adj_5959), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n75269));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i59651_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i60243_2_lut (.I0(n24_adj_5959), .I1(n6903), .I2(GND_net), 
            .I3(GND_net), .O(n75272));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i60243_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n75272), .I1(n75269), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5965), .O(n64972));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i16571_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n23094), .I3(GND_net), .O(n30785));   // verilog/coms.v(130[12] 305[6])
    defparam i16571_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n59247));
    SB_LUT4 encoder0_position_30__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n59674), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_14_lut (.I0(GND_net), .I1(n1422), 
            .I2(VCC_net), .I3(n59246), .O(n1489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_10 (.CI(n59674), .I0(n2626), 
            .I1(VCC_net), .CO(n59675));
    SB_LUT4 encoder0_position_30__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n59673), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n59041), .I0(encoder0_position_scaled[11]), 
            .I1(n14), .CO(n59042));
    SB_LUT4 encoder0_position_30__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n59245), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_13 (.CI(n59245), .I0(n1423), 
            .I1(VCC_net), .CO(n59246));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5710), .I3(n59040), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5957));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_CARRY encoder0_position_30__I_0_add_1771_9 (.CI(n59673), .I0(n2627), 
            .I1(VCC_net), .CO(n59674));
    SB_LUT4 encoder0_position_30__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n59672), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_8 (.CI(n59672), .I0(n2628), 
            .I1(VCC_net), .CO(n59673));
    SB_LUT4 encoder0_position_30__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n59671), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n59244), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_12 (.CI(n59244), .I0(n1424), 
            .I1(VCC_net), .CO(n59245));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n59040), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5710), .CO(n59041));
    SB_CARRY encoder0_position_30__I_0_add_1771_7 (.CI(n59671), .I0(n2629), 
            .I1(GND_net), .CO(n59672));
    SB_LUT4 encoder0_position_30__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n59670), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_6 (.CI(n59670), .I0(n2630), 
            .I1(GND_net), .CO(n59671));
    SB_LUT4 i20492_3_lut (.I0(n16_adj_5863), .I1(PWMLimit[8]), .I2(setpoint[8]), 
            .I3(GND_net), .O(n34689));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i20492_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5709), .I3(n59039), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_2_lut_adj_1823 (.I0(PWMLimit[16]), .I1(setpoint[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i7_2_lut_adj_1823.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n59039), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5709), .CO(n59040));
    SB_LUT4 i63017_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78873));
    defparam i63017_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_2_lut_adj_1824 (.I0(PWMLimit[12]), .I1(setpoint[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5866));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i9_2_lut_adj_1824.LUT_INIT = 16'h6666;
    SB_LUT4 i23696_3_lut (.I0(n20_adj_5864), .I1(PWMLimit[10]), .I2(setpoint[10]), 
            .I3(GND_net), .O(n22_adj_5865));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i23696_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i12_2_lut (.I0(PWMLimit[4]), .I1(n475), .I2(GND_net), .I3(GND_net), 
            .O(n35782));
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21973_3_lut (.I0(n24_adj_5875), .I1(PWMLimit[12]), .I2(n467), 
            .I3(GND_net), .O(n36147));
    defparam i21973_3_lut.LUT_INIT = 16'hb2b2;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n59669), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_5 (.CI(n59669), .I0(n2631), 
            .I1(VCC_net), .CO(n59670));
    SB_LUT4 encoder0_position_30__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n59668), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_4 (.CI(n59668), .I0(n2632), 
            .I1(GND_net), .CO(n59669));
    SB_LUT4 encoder0_position_30__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n59667), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n59243), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_3 (.CI(n59667), .I0(n2633), 
            .I1(VCC_net), .CO(n59668));
    SB_LUT4 encoder0_position_30__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n59667));
    SB_CARRY encoder0_position_30__I_0_add_967_11 (.CI(n59243), .I0(n1425), 
            .I1(VCC_net), .CO(n59244));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5708), .I3(n59038), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_25_lut (.I0(n78616), .I1(n2511), 
            .I2(VCC_net), .I3(n59666), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n59665), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_24 (.CI(n59665), .I0(n2512), 
            .I1(VCC_net), .CO(n59666));
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n59664), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n59242), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_23 (.CI(n59664), .I0(n2513), 
            .I1(VCC_net), .CO(n59665));
    SB_LUT4 encoder0_position_30__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n59663), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_22 (.CI(n59663), .I0(n2514), 
            .I1(VCC_net), .CO(n59664));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n59038), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5708), .CO(n59039));
    SB_LUT4 encoder0_position_30__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n59662), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_21 (.CI(n59662), .I0(n2515), 
            .I1(VCC_net), .CO(n59663));
    SB_CARRY encoder0_position_30__I_0_add_967_10 (.CI(n59242), .I0(n1426), 
            .I1(VCC_net), .CO(n59243));
    SB_LUT4 encoder0_position_30__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n59661), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n59241), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_20 (.CI(n59661), .I0(n2516), 
            .I1(VCC_net), .CO(n59662));
    SB_LUT4 encoder0_position_30__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n59660), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18), .I3(n59037), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_19 (.CI(n59660), .I0(n2517), 
            .I1(VCC_net), .CO(n59661));
    SB_LUT4 encoder0_position_30__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n59659), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_18 (.CI(n59659), .I0(n2518), 
            .I1(VCC_net), .CO(n59660));
    SB_LUT4 encoder0_position_30__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n59658), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_17 (.CI(n59658), .I0(n2519), 
            .I1(VCC_net), .CO(n59659));
    SB_LUT4 encoder0_position_30__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n59657), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_9 (.CI(n59241), .I0(n1427), 
            .I1(VCC_net), .CO(n59242));
    SB_CARRY encoder0_position_30__I_0_add_1704_16 (.CI(n59657), .I0(n2520), 
            .I1(VCC_net), .CO(n59658));
    SB_LUT4 encoder0_position_30__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n59656), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_15 (.CI(n59656), .I0(n2521), 
            .I1(VCC_net), .CO(n59657));
    SB_LUT4 encoder0_position_30__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n59655), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_14 (.CI(n59655), .I0(n2522), 
            .I1(VCC_net), .CO(n59656));
    SB_LUT4 encoder0_position_30__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n59654), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n59240), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_2_lut (.I0(n299_adj_5790), .I1(n247), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_5868));
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1704_13 (.CI(n59654), .I0(n2523), 
            .I1(VCC_net), .CO(n59655));
    SB_LUT4 encoder0_position_30__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n59653), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_12 (.CI(n59653), .I0(n2524), 
            .I1(VCC_net), .CO(n59654));
    SB_LUT4 encoder0_position_30__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n59652), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31409_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n45504));
    defparam i31409_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_30__I_0_add_1704_11 (.CI(n59652), .I0(n2525), 
            .I1(VCC_net), .CO(n59653));
    SB_CARRY encoder0_position_30__I_0_add_967_8 (.CI(n59240), .I0(n1428), 
            .I1(VCC_net), .CO(n59241));
    SB_LUT4 encoder0_position_30__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n59239), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n59651), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_10 (.CI(n59651), .I0(n2526), 
            .I1(VCC_net), .CO(n59652));
    SB_LUT4 encoder0_position_30__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n59650), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_9 (.CI(n59650), .I0(n2527), 
            .I1(VCC_net), .CO(n59651));
    SB_LUT4 encoder0_position_30__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n59649), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_8 (.CI(n59649), .I0(n2528), 
            .I1(VCC_net), .CO(n59650));
    SB_LUT4 encoder0_position_30__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n59648), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1825 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[11] [6]), 
            .I2(n66979), .I3(n6_adj_5934), .O(n27089));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1825.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_30__I_0_add_1704_7 (.CI(n59648), .I0(n2529), 
            .I1(GND_net), .CO(n59649));
    SB_LUT4 encoder0_position_30__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n59647), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_7 (.CI(n59239), .I0(n1429), 
            .I1(GND_net), .CO(n59240));
    SB_CARRY encoder0_position_30__I_0_add_1704_6 (.CI(n59647), .I0(n2530), 
            .I1(GND_net), .CO(n59648));
    SB_LUT4 encoder0_position_30__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n59646), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_5 (.CI(n59646), .I0(n2531), 
            .I1(VCC_net), .CO(n59647));
    SB_LUT4 encoder0_position_30__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n59238), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n59645), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_6 (.CI(n59238), .I0(n1430), 
            .I1(GND_net), .CO(n59239));
    SB_CARRY encoder0_position_30__I_0_add_1704_4 (.CI(n59645), .I0(n2532), 
            .I1(GND_net), .CO(n59646));
    SB_LUT4 encoder0_position_30__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n59644), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n59237), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_3 (.CI(n59644), .I0(n2533), 
            .I1(VCC_net), .CO(n59645));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n59037), .I0(encoder0_position_scaled[7]), 
            .I1(n18), .CO(n59038));
    SB_CARRY encoder0_position_30__I_0_add_967_5 (.CI(n59237), .I0(n1431), 
            .I1(VCC_net), .CO(n59238));
    SB_LUT4 encoder0_position_30__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23148_3_lut (.I0(n239), .I1(n291), .I2(n284), .I3(GND_net), 
            .O(n37306));
    defparam i23148_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n59644));
    SB_LUT4 i23149_3_lut (.I0(n37306), .I1(IntegralLimit[18]), .I2(n258), 
            .I3(GND_net), .O(n37307));
    defparam i23149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1826 (.I0(n37307), .I1(Ki[4]), .I2(GND_net), 
            .I3(GND_net), .O(n347_adj_5909));
    defparam i1_2_lut_adj_1826.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n59236), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28879_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n5_adj_5951));   // verilog/coms.v(105[12:33])
    defparam i28879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n1));   // verilog/coms.v(105[12:33])
    defparam i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_967_4 (.CI(n59236), .I0(n1432), 
            .I1(GND_net), .CO(n59237));
    SB_LUT4 i30474_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i30474_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n59235), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19), .I3(n59036), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62791_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78647));
    defparam i62791_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_967_3 (.CI(n59235), .I0(n1433), 
            .I1(VCC_net), .CO(n59236));
    SB_CARRY add_151_12 (.CI(n58886), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n58887));
    SB_LUT4 encoder0_position_30__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n59036), .I0(encoder0_position_scaled[6]), 
            .I1(n19), .CO(n59037));
    SB_LUT4 i8_2_lut (.I0(deadband[12]), .I1(n467), .I2(GND_net), .I3(GND_net), 
            .O(n25_adj_5872));
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n70868));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n59035), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i63081_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78937));
    defparam i63081_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62521_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78377));
    defparam i62521_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5782));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_30__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n59235));
    SB_LUT4 encoder0_position_30__I_0_add_900_13_lut (.I0(n78888), .I1(n1323), 
            .I2(VCC_net), .I3(n59234), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n59233), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_12 (.CI(n59233), .I0(n1324), 
            .I1(VCC_net), .CO(n59234));
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5964));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1827 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n70954));
    defparam i1_2_lut_adj_1827.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n59035), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n59036));
    SB_LUT4 encoder0_position_30__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i63016_4_lut (.I0(n70954), .I1(n1125), .I2(n70868), .I3(n45504), 
            .O(n1158));
    defparam i63016_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 mux_3812_i22_3_lut (.I0(encoder0_position[21]), .I1(n11_adj_5739), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n936));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31333_3_lut (.I0(n937), .I1(n1232_adj_5844), .I2(n1233_adj_5845), 
            .I3(GND_net), .O(n45428));
    defparam i31333_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i6_4_lut (.I0(dti_counter[7]), .I1(dti_counter[4]), .I2(dti_counter[5]), 
            .I3(dti_counter[6]), .O(n14_adj_5963));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1828 (.I0(dti_counter[0]), .I1(n14_adj_5963), .I2(n10_adj_5964), 
            .I3(dti_counter[3]), .O(n23188));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n59232), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_5 (.CI(n58879), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n58880));
    SB_CARRY encoder0_position_30__I_0_add_900_11 (.CI(n59232), .I0(n1325), 
            .I1(VCC_net), .CO(n59233));
    SB_LUT4 mux_1677_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), 
            .I3(GND_net), .O(n11914));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n12492));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 n11851_bdd_4_lut (.I0(n11851), .I1(current[15]), .I2(duty[18]), 
            .I3(n11849), .O(n79636));
    defparam n11851_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n59034), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21595_3_lut (.I0(n8_adj_5870), .I1(deadband[4]), .I2(n475), 
            .I3(GND_net), .O(n10_adj_5871));
    defparam i21595_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i1_3_lut_adj_1829 (.I0(n1226_adj_5838), .I1(n1227_adj_5839), 
            .I2(n1228_adj_5840), .I3(GND_net), .O(n70962));
    defparam i1_3_lut_adj_1829.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_1677_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n12490));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n28130), 
            .D(n1229), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n28130), 
            .D(n1228), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 mux_1677_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n12488));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n12486));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i63114_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78970));
    defparam i63114_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1677_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n12484));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i59712_2_lut_4_lut (.I0(duty[6]), .I1(n304), .I2(duty[5]), 
            .I3(n305), .O(n75568));
    defparam i59712_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1830 (.I0(n1229_adj_5841), .I1(n45428), .I2(n1230_adj_5842), 
            .I3(n1231_adj_5843), .O(n68433));
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'ha080;
    SB_LUT4 i63031_4_lut (.I0(n1225_adj_5837), .I1(n1224_adj_5836), .I2(n68433), 
            .I3(n70962), .O(n1257));
    defparam i63031_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_1677_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n12482));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233_adj_5845));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31329_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n45424));
    defparam i31329_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n70784));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'hfffe;
    SB_LUT4 i16809_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n31023));   // verilog/coms.v(130[12] 305[6])
    defparam i16809_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1677_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n12480));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n12478));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n1329), .I1(n45424), .I2(n1330), .I3(n1331), 
            .O(n68431));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'ha080;
    SB_LUT4 mux_1677_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n12476));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n12474));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n12472));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i63047_4_lut (.I0(n68431), .I1(n1323), .I2(n1324), .I3(n70784), 
            .O(n1356));
    defparam i63047_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i844_3_lut (.I0(n1233_adj_5845), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31401_4_lut (.I0(n939), .I1(n1431), .I2(n1432), .I3(n1433), 
            .O(n45496));
    defparam i31401_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1833 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n70976));
    defparam i1_2_lut_adj_1833.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1834 (.I0(n1429), .I1(n70976), .I2(n45496), .I3(n1430), 
            .O(n70978));
    defparam i1_4_lut_adj_1834.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_adj_1835 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(GND_net), 
            .O(n70984));
    defparam i1_3_lut_adj_1835.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_1677_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n12470));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i63064_4_lut (.I0(n1423), .I1(n70984), .I2(n70978), .I3(n1422), 
            .O(n1455));
    defparam i63064_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31238_3_lut (.I0(n940), .I1(n1532), .I2(n1533), .I3(GND_net), 
            .O(n45330));
    defparam i31238_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_1677_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n12468));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1836 (.I0(n1529), .I1(n45330), .I2(n1530), .I3(n1531), 
            .O(n68441));
    defparam i1_4_lut_adj_1836.LUT_INIT = 16'ha080;
    SB_LUT4 i1_3_lut_adj_1837 (.I0(n1522), .I1(n1524), .I2(n1526), .I3(GND_net), 
            .O(n70896));
    defparam i1_3_lut_adj_1837.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1838 (.I0(n1523), .I1(n1525), .I2(n1528), .I3(n1527), 
            .O(n70972));
    defparam i1_4_lut_adj_1838.LUT_INIT = 16'hfffe;
    SB_LUT4 i62995_4_lut (.I0(n70972), .I1(n1521), .I2(n70896), .I3(n68441), 
            .O(n1554));
    defparam i62995_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1840_3_lut (.I0(n2709), .I1(n2776), 
            .I2(n2742), .I3(GND_net), .O(n2808));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n12466));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31341_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n45436));
    defparam i31341_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_1677_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n12464));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n12462));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n12460));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i18_3_lut.LUT_INIT = 16'h3535;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i63148_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n79004));
    defparam i63148_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n28130), 
            .D(n1227), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i62495_1_lut (.I0(n45484), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78351));
    defparam i62495_1_lut.LUT_INIT = 16'h5555;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5942));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2189_3_lut (.I0(n3218), .I1(n3285), 
            .I2(n3237), .I3(GND_net), .O(n35_adj_5948));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_adj_1839 (.I0(n3231), .I1(n75097), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5915));
    defparam i16_4_lut_adj_1839.LUT_INIT = 16'hac0c;
    SB_LUT4 i1_4_lut_adj_1840 (.I0(n1625), .I1(n1626), .I2(n1627), .I3(n1628), 
            .O(n71020));
    defparam i1_4_lut_adj_1840.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1841 (.I0(n1629), .I1(n45436), .I2(n1630), .I3(n1631), 
            .O(n68452));
    defparam i1_4_lut_adj_1841.LUT_INIT = 16'ha080;
    SB_LUT4 i16669_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n30883));   // verilog/coms.v(130[12] 305[6])
    defparam i16669_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i59562_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n75093));
    defparam i59562_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 n79636_bdd_4_lut (.I0(n79636), .I1(duty[15]), .I2(n4915), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[15]));
    defparam n79636_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i2191_3_lut (.I0(n3220), .I1(n3287), 
            .I2(n3237), .I3(GND_net), .O(n31_adj_5947));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5943));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5944));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1842 (.I0(n1623), .I1(n1624), .I2(n68452), .I3(n71020), 
            .O(n71026));
    defparam i1_4_lut_adj_1842.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i62809_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n71026), 
            .O(n1653));
    defparam i62809_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1843 (.I0(n1724), .I1(n1723), .I2(n1728), .I3(n1726), 
            .O(n69575));
    defparam i1_4_lut_adj_1843.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i31343_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n45438));
    defparam i31343_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1844 (.I0(n69575), .I1(n1722), .I2(n1725), .I3(n1727), 
            .O(n70904));
    defparam i1_4_lut_adj_1844.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1845 (.I0(n1729), .I1(n70904), .I2(n45438), .I3(n1730), 
            .O(n70906));
    defparam i1_4_lut_adj_1845.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_30__I_0_i2194_3_lut (.I0(n3223), .I1(n3290), 
            .I2(n3237), .I3(GND_net), .O(n25_adj_5945));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1846 (.I0(n3226), .I1(n25_adj_5945), .I2(n3293), 
            .I3(n3237), .O(n70682));
    defparam i1_4_lut_adj_1846.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1847 (.I0(n3222), .I1(n15_adj_5943), .I2(n3289), 
            .I3(n3237), .O(n70680));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i1907_3_lut (.I0(n2808), .I1(n2875), 
            .I2(n2841), .I3(GND_net), .O(n2907));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1848 (.I0(n3219), .I1(n31_adj_5947), .I2(n3286), 
            .I3(n3237), .O(n70686));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(n3215), .I1(n17_adj_5944), .I2(n3282), 
            .I3(n3237), .O(n70688));
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2192_3_lut (.I0(n3221), .I1(n3288), 
            .I2(n3237), .I3(GND_net), .O(n29_adj_5946));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59706_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n75562));
    defparam i59706_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_30__I_0_i2187_3_lut (.I0(n3216), .I1(n3283), 
            .I2(n3237), .I3(GND_net), .O(n39_adj_5949));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1850 (.I0(n3217), .I1(n39_adj_5949), .I2(n3284), 
            .I3(n3237), .O(n71292));
    defparam i1_4_lut_adj_1850.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1851 (.I0(n3213), .I1(n71292), .I2(n3280), .I3(n3237), 
            .O(n71294));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1852 (.I0(n3225), .I1(n13_adj_5942), .I2(n3292), 
            .I3(n3237), .O(n70690));
    defparam i1_4_lut_adj_1852.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1853 (.I0(n3214), .I1(n35_adj_5948), .I2(n3281), 
            .I3(n3237), .O(n70692));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1854 (.I0(n75093), .I1(n5_adj_5915), .I2(n75094), 
            .I3(n3237), .O(n62972));
    defparam i1_4_lut_adj_1854.LUT_INIT = 16'h88c0;
    SB_LUT4 i1_4_lut_adj_1855 (.I0(n3224), .I1(n29_adj_5946), .I2(n3291), 
            .I3(n3237), .O(n70684));
    defparam i1_4_lut_adj_1855.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1856 (.I0(n70688), .I1(n70686), .I2(n70680), 
            .I3(n70682), .O(n70702));
    defparam i1_4_lut_adj_1856.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1857 (.I0(n70684), .I1(n62972), .I2(n70692), 
            .I3(n70690), .O(n70704));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2182_3_lut (.I0(n3211), .I1(n3278), 
            .I2(n3237), .I3(GND_net), .O(n49));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1858 (.I0(n71294), .I1(n3212), .I2(n3279), .I3(n3237), 
            .O(n69393));
    defparam i1_4_lut_adj_1858.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_30__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1859 (.I0(n69393), .I1(n49), .I2(n70704), .I3(n70702), 
            .O(n70710));
    defparam i1_4_lut_adj_1859.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1860 (.I0(n3210), .I1(n70710), .I2(n3277), .I3(n3237), 
            .O(n70712));
    defparam i1_4_lut_adj_1860.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1861 (.I0(n3209), .I1(n70712), .I2(n3276), .I3(n3237), 
            .O(n70714));
    defparam i1_4_lut_adj_1861.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1862 (.I0(n3208), .I1(n70714), .I2(n3275), .I3(n3237), 
            .O(n70716));
    defparam i1_4_lut_adj_1862.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1863 (.I0(n3207), .I1(n70716), .I2(n3274), .I3(n3237), 
            .O(n70718));
    defparam i1_4_lut_adj_1863.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62498_4_lut (.I0(n61), .I1(n72039), .I2(n59), .I3(n70718), 
            .O(n45484));
    defparam i62498_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_DFF read_197 (.Q(state_7__N_3918[0]), .C(clk16MHz), .D(n69981));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n67625));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n59231), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_10 (.CI(n59231), .I0(n1326), 
            .I1(VCC_net), .CO(n59232));
    SB_LUT4 encoder0_position_30__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i24_3_lut (.I0(encoder0_position[23]), .I1(n9_adj_5741), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n934));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11851_bdd_4_lut_63686 (.I0(n11851), .I1(current[15]), .I2(duty[17]), 
            .I3(n11849), .O(n79624));
    defparam n11851_bdd_4_lut_63686.LUT_INIT = 16'he4aa;
    SB_LUT4 n79624_bdd_4_lut (.I0(n79624), .I1(duty[14]), .I2(n4916), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[14]));
    defparam n79624_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i1_3_lut (.I0(encoder0_position[0]), .I1(n32), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1864 (.I0(n3226), .I1(n3227), .I2(GND_net), .I3(GND_net), 
            .O(n71298));
    defparam i1_2_lut_adj_1864.LUT_INIT = 16'heeee;
    SB_LUT4 i31278_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n45370));
    defparam i31278_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1865 (.I0(n3225), .I1(n71298), .I2(n3228), .I3(n3224), 
            .O(n71302));
    defparam i1_4_lut_adj_1865.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1866 (.I0(n3229), .I1(n45370), .I2(n3230), .I3(n3231), 
            .O(n68582));
    defparam i1_4_lut_adj_1866.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1867 (.I0(n3219), .I1(n3220), .I2(n3221), .I3(n71302), 
            .O(n71308));
    defparam i1_4_lut_adj_1867.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1868 (.I0(n3217), .I1(n3218), .I2(n71308), .I3(n68582), 
            .O(n71314));
    defparam i1_4_lut_adj_1868.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1869 (.I0(n3214), .I1(n3215), .I2(n3216), .I3(n71314), 
            .O(n71320));
    defparam i1_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1870 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n71320), 
            .O(n71326));
    defparam i1_4_lut_adj_1870.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1871 (.I0(n3213), .I1(n3209), .I2(n3222), .I3(n3223), 
            .O(n68753));
    defparam i1_4_lut_adj_1871.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1872 (.I0(n3207), .I1(n68753), .I2(n3208), .I3(n71326), 
            .O(n71332));
    defparam i1_4_lut_adj_1872.LUT_INIT = 16'hfffe;
    SB_LUT4 i63179_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n71332), 
            .O(n3237));
    defparam i63179_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i62540_4_lut (.I0(n1720), .I1(n1719), .I2(n70906), .I3(n1721), 
            .O(n1752));
    defparam i62540_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i31345_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n45440));
    defparam i31345_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1873 (.I0(n1825), .I1(n1827), .I2(n1826), .I3(n1828), 
            .O(n71038));
    defparam i1_4_lut_adj_1873.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1874 (.I0(n1829), .I1(n45440), .I2(n1830), .I3(n1831), 
            .O(n68490));
    defparam i1_4_lut_adj_1874.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_3_lut_adj_1875 (.I0(n1820), .I1(n1821), .I2(n1822_adj_5851), 
            .I3(GND_net), .O(n71048));
    defparam i1_3_lut_adj_1875.LUT_INIT = 16'hfefe;
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1876 (.I0(n1823), .I1(n68490), .I2(n1824_adj_5852), 
            .I3(n71038), .O(n71044));
    defparam i1_4_lut_adj_1876.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i62637_4_lut (.I0(n1818), .I1(n71044), .I2(n71048), .I3(n1819), 
            .O(n1851));
    defparam i62637_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1877 (.I0(n1928), .I1(n1926), .I2(n1924), .I3(n1927), 
            .O(n70878));
    defparam i1_4_lut_adj_1877.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i31260_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n45352));
    defparam i31260_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1878 (.I0(n1922), .I1(n70878), .I2(n1923), .I3(n1925), 
            .O(n70882));
    defparam i1_4_lut_adj_1878.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n28130), 
            .D(n1226), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n28130), 
            .D(n1225), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n28130), 
            .D(n1224), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n28130), 
            .D(n1223), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n28130), 
            .D(n1222), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n28130), 
            .D(n1221), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n28130), 
            .D(n1220), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n28130), 
            .D(n1219), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i1_4_lut_adj_1879 (.I0(n1929), .I1(n45352), .I2(n1930), .I3(n1931), 
            .O(n68474));
    defparam i1_4_lut_adj_1879.LUT_INIT = 16'ha080;
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n28130), 
            .D(n1218), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n28130), 
            .D(n1217), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n28130), 
            .D(n1216), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n28130), 
            .D(n1215), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n28130), 
            .D(n1214), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n28130), 
            .D(n1213), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n28130), 
            .D(n1212), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n28130), 
            .D(n1211), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n28130), 
            .D(n1210), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n28130), 
            .D(n1209), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n28130), 
            .D(n1208), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR dti_counter_2038__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n28174), 
            .D(n44), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n28174), 
            .D(n43), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n28174), 
            .D(n42), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n28174), 
            .D(n41_adj_5933), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n28174), 
            .D(n40_adj_5932), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n28174), 
            .D(n39_adj_5931), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n28174), 
            .D(n38_adj_5930), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n59034), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n59035));
    SB_LUT4 encoder0_position_30__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11851_bdd_4_lut_63676 (.I0(n11851), .I1(current[15]), .I2(duty[16]), 
            .I3(n11849), .O(n79618));
    defparam n11851_bdd_4_lut_63676.LUT_INIT = 16'he4aa;
    SB_LUT4 n79618_bdd_4_lut (.I0(n79618), .I1(duty[13]), .I2(n4917), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[13]));
    defparam n79618_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i2_3_lut (.I0(encoder0_position[1]), .I1(n31), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1880 (.I0(n3116), .I1(n3124), .I2(n3125), .I3(n3122), 
            .O(n70808));
    defparam i1_4_lut_adj_1880.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11851_bdd_4_lut_63671 (.I0(n11851), .I1(current[15]), .I2(duty[15]), 
            .I3(n11849), .O(n79612));
    defparam n11851_bdd_4_lut_63671.LUT_INIT = 16'he4aa;
    SB_LUT4 n79612_bdd_4_lut (.I0(n79612), .I1(duty[12]), .I2(n4918), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[12]));
    defparam n79612_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1881 (.I0(n3120), .I1(n3121), .I2(n3127), .I3(n3123), 
            .O(n70810));
    defparam i1_4_lut_adj_1881.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1882 (.I0(n3117), .I1(n3115), .I2(n3126), .I3(n3128), 
            .O(n70806));
    defparam i1_4_lut_adj_1882.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1883 (.I0(n70808), .I1(n3119), .I2(n3114), .I3(n3118), 
            .O(n70812));
    defparam i1_4_lut_adj_1883.LUT_INIT = 16'hfffe;
    SB_LUT4 dti_counter_2038_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n60154), .O(n38_adj_5930)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2038_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n60153), .O(n39_adj_5931)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31373_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n45468));
    defparam i31373_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1884 (.I0(n70812), .I1(n3113), .I2(n70806), .I3(n70810), 
            .O(n70818));
    defparam i1_4_lut_adj_1884.LUT_INIT = 16'hfffe;
    SB_CARRY dti_counter_2038_add_4_8 (.CI(n60153), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n60154));
    SB_LUT4 encoder0_position_30__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231_adj_5843));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2038_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n60152), .O(n40_adj_5932)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11851_bdd_4_lut_63666 (.I0(n11851), .I1(current[11]), .I2(duty[14]), 
            .I3(n11849), .O(n79606));
    defparam n11851_bdd_4_lut_63666.LUT_INIT = 16'he4aa;
    SB_LUT4 n79606_bdd_4_lut (.I0(n79606), .I1(duty[11]), .I2(n4919), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[11]));
    defparam n79606_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i842_3_lut (.I0(n1231_adj_5843), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1885 (.I0(n1920), .I1(n68474), .I2(n1921), .I3(n70882), 
            .O(n70888));
    defparam i1_4_lut_adj_1885.LUT_INIT = 16'hfffe;
    SB_CARRY dti_counter_2038_add_4_7 (.CI(n60152), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n60153));
    SB_LUT4 i1_4_lut_adj_1886 (.I0(n3129), .I1(n45468), .I2(n3130), .I3(n3131), 
            .O(n68536));
    defparam i1_4_lut_adj_1886.LUT_INIT = 16'ha080;
    SB_LUT4 i62520_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n70888), 
            .O(n1950));
    defparam i62520_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1887 (.I0(n3111), .I1(n68536), .I2(n3112), .I3(n70818), 
            .O(n70824));
    defparam i1_4_lut_adj_1887.LUT_INIT = 16'hfffe;
    SB_LUT4 i31431_4_lut (.I0(n945), .I1(n2031), .I2(n2032), .I3(n2033), 
            .O(n45526));
    defparam i31431_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 dti_counter_2038_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n60151), .O(n41_adj_5933)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1888 (.I0(n2024), .I1(n2025), .I2(n2027), .I3(GND_net), 
            .O(n71100));
    defparam i1_3_lut_adj_1888.LUT_INIT = 16'hfefe;
    SB_CARRY dti_counter_2038_add_4_6 (.CI(n60151), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n60152));
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n70824), 
            .O(n70830));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'hfffe;
    SB_LUT4 i63147_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n70830), 
            .O(n3138));
    defparam i63147_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 dti_counter_2038_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n60150), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11851_bdd_4_lut_63661 (.I0(n11851), .I1(current[10]), .I2(duty[13]), 
            .I3(n11849), .O(n79600));
    defparam n11851_bdd_4_lut_63661.LUT_INIT = 16'he4aa;
    SB_LUT4 n79600_bdd_4_lut (.I0(n79600), .I1(duty[10]), .I2(n4920), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[10]));
    defparam n79600_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1890 (.I0(n2028), .I1(n2026), .I2(GND_net), .I3(GND_net), 
            .O(n71214));
    defparam i1_2_lut_adj_1890.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1891 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n71214), 
            .O(n71220));
    defparam i1_4_lut_adj_1891.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1892 (.I0(n2029), .I1(n71100), .I2(n45526), .I3(n2030), 
            .O(n71102));
    defparam i1_4_lut_adj_1892.LUT_INIT = 16'heccc;
    SB_CARRY dti_counter_2038_add_4_5 (.CI(n60150), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n60151));
    SB_LUT4 i1_4_lut_adj_1893 (.I0(n2019), .I1(n2018), .I2(n2020), .I3(n71220), 
            .O(n69738));
    defparam i1_4_lut_adj_1893.LUT_INIT = 16'hfffe;
    SB_LUT4 i62901_4_lut (.I0(n2017), .I1(n2016), .I2(n69738), .I3(n71102), 
            .O(n2049));
    defparam i62901_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1894 (.I0(n2125), .I1(n2122), .I2(n2124), .I3(GND_net), 
            .O(n70732));
    defparam i1_3_lut_adj_1894.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR dti_counter_2038__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n28174), 
            .D(n45), .R(n29438));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1895 (.I0(n2127), .I1(n2128), .I2(n2126), .I3(n2123), 
            .O(n70734));
    defparam i1_4_lut_adj_1895.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11851_bdd_4_lut_63656 (.I0(n11851), .I1(current[9]), .I2(duty[12]), 
            .I3(n11849), .O(n79594));
    defparam n11851_bdd_4_lut_63656.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31361_3_lut (.I0(n946), .I1(n2132), .I2(n2133), .I3(GND_net), 
            .O(n45456));
    defparam i31361_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1896 (.I0(n2120), .I1(n2121), .I2(n70734), .I3(n70732), 
            .O(n70740));
    defparam i1_4_lut_adj_1896.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1897 (.I0(n2129), .I1(n45456), .I2(n2130), .I3(n2131), 
            .O(n68492));
    defparam i1_4_lut_adj_1897.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1898 (.I0(n2118), .I1(n68492), .I2(n2119), .I3(n70740), 
            .O(n70746));
    defparam i1_4_lut_adj_1898.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62925_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n70746), 
            .O(n2148));
    defparam i62925_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2038_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n60149), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n79594_bdd_4_lut (.I0(n79594), .I1(duty[9]), .I2(n4921), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n79594_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31355_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n45450));
    defparam i31355_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1899 (.I0(n2229), .I1(n45450), .I2(n2230), .I3(n2231), 
            .O(n68518));
    defparam i1_4_lut_adj_1899.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1900 (.I0(n2221), .I1(n2223), .I2(n2227), .I3(n2228), 
            .O(n71112));
    defparam i1_4_lut_adj_1900.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1901 (.I0(n2222), .I1(n2226), .I2(n2224), .I3(n2225), 
            .O(n71158));
    defparam i1_4_lut_adj_1901.LUT_INIT = 16'hfffe;
    SB_CARRY dti_counter_2038_add_4_4 (.CI(n60149), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n60150));
    SB_LUT4 encoder0_position_30__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n59230), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2038_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n60148), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_9 (.CI(n59230), .I0(n1327), 
            .I1(VCC_net), .CO(n59231));
    SB_LUT4 encoder0_position_30__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5767));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1902 (.I0(n2219), .I1(n2220), .I2(n71112), .I3(n68518), 
            .O(n71118));
    defparam i1_4_lut_adj_1902.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1903 (.I0(n2216), .I1(n2217), .I2(n2218), .I3(n71158), 
            .O(n71164));
    defparam i1_4_lut_adj_1903.LUT_INIT = 16'hfffe;
    SB_LUT4 i62875_4_lut (.I0(n2215), .I1(n71164), .I2(n71118), .I3(n2214), 
            .O(n2247));
    defparam i62875_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 n11851_bdd_4_lut_63651 (.I0(n11851), .I1(current[8]), .I2(duty[11]), 
            .I3(n11849), .O(n79588));
    defparam n11851_bdd_4_lut_63651.LUT_INIT = 16'he4aa;
    SB_LUT4 n79588_bdd_4_lut (.I0(n79588), .I1(duty[8]), .I2(n4922), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n79588_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i59863_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n75719));
    defparam i59863_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_30__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1904 (.I0(n2328), .I1(n2325), .I2(GND_net), .I3(GND_net), 
            .O(n70840));
    defparam i1_2_lut_adj_1904.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5765));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1905 (.I0(n2322), .I1(n2323), .I2(n2324), .I3(n2326), 
            .O(n70846));
    defparam i1_4_lut_adj_1905.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_2038_add_4_3 (.CI(n60148), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n60149));
    SB_LUT4 encoder0_position_30__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n59229), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_8 (.CI(n59229), .I0(n1328), 
            .I1(VCC_net), .CO(n59230));
    SB_LUT4 encoder0_position_30__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1906 (.I0(n2321), .I1(n70840), .I2(n2320), .I3(n2327), 
            .O(n70848));
    defparam i1_4_lut_adj_1906.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2038_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n59228), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_900_7 (.CI(n59228), .I0(n1329), 
            .I1(GND_net), .CO(n59229));
    SB_LUT4 i31371_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n45466));
    defparam i31371_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1907 (.I0(n3025), .I1(n3027), .I2(n3028), .I3(n3026), 
            .O(n71250));
    defparam i1_4_lut_adj_1907.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1908 (.I0(n71250), .I1(n3023), .I2(n3024), .I3(GND_net), 
            .O(n71252));
    defparam i1_3_lut_adj_1908.LUT_INIT = 16'hfefe;
    SB_CARRY dti_counter_2038_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n60148));
    SB_LUT4 i1_4_lut_adj_1909 (.I0(n3029), .I1(n45466), .I2(n3030), .I3(n3031), 
            .O(n68571));
    defparam i1_4_lut_adj_1909.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1910 (.I0(n3020), .I1(n3021), .I2(n3022), .I3(n71252), 
            .O(n71258));
    defparam i1_4_lut_adj_1910.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1911 (.I0(n3018), .I1(n3019), .I2(n71258), .I3(n68571), 
            .O(n71264));
    defparam i1_4_lut_adj_1911.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1912 (.I0(n3015), .I1(n3016), .I2(n3017), .I3(n71264), 
            .O(n71270));
    defparam i1_4_lut_adj_1912.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1913 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n71270), 
            .O(n71276));
    defparam i1_4_lut_adj_1913.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1914 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n71276), 
            .O(n71282));
    defparam i1_4_lut_adj_1914.LUT_INIT = 16'hfffe;
    SB_LUT4 i63113_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n71282), 
            .O(n3039));
    defparam i63113_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n59227), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n12458));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i19_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_30__I_0_add_900_6 (.CI(n59227), .I0(n1330), 
            .I1(GND_net), .CO(n59228));
    SB_LUT4 i62756_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78612));
    defparam i62756_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1677_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n12456));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n59226), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_900_5 (.CI(n59226), .I0(n1331), 
            .I1(VCC_net), .CO(n59227));
    SB_LUT4 encoder0_position_30__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n59225), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_4 (.CI(n59225), .I0(n1332), 
            .I1(GND_net), .CO(n59226));
    SB_LUT4 encoder0_position_30__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n59224), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62724_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78580));
    defparam i62724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n12454));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i62607_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78463));
    defparam i62607_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1677_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n12452));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i62690_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78546));
    defparam i62690_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_900_3 (.CI(n59224), .I0(n1333), 
            .I1(VCC_net), .CO(n59225));
    SB_LUT4 mux_1677_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n12450));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n59224));
    SB_LUT4 encoder0_position_30__I_0_add_833_12_lut (.I0(n78873), .I1(n1224_adj_5836), 
            .I2(VCC_net), .I3(n59223), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n11851_bdd_4_lut_63646 (.I0(n11851), .I1(current[7]), .I2(duty[10]), 
            .I3(n11849), .O(n79582));
    defparam n11851_bdd_4_lut_63646.LUT_INIT = 16'he4aa;
    SB_LUT4 i62661_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78517));
    defparam i62661_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62832_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78688));
    defparam i62832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62872_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78728));
    defparam i62872_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62922_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78778));
    defparam i62922_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62898_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78754));
    defparam i62898_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62517_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78373));
    defparam i62517_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_91[10]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i62634_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78490));
    defparam i62634_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n64972));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225_adj_5837), 
            .I2(VCC_net), .I3(n59222), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_11 (.CI(n59222), .I0(n1225_adj_5837), 
            .I1(VCC_net), .CO(n59223));
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30748));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226_adj_5838), 
            .I2(VCC_net), .I3(n59221), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_243_i14_3_lut (.I0(encoder0_position_scaled[13]), .I1(motor_state_23__N_91[13]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i14_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_30__I_0_add_833_10 (.CI(n59221), .I0(n1226_adj_5838), 
            .I1(VCC_net), .CO(n59222));
    SB_LUT4 mux_245_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5966), 
            .I2(commutation_state_prev[0]), .I3(dti_N_404), .O(n28027));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 encoder0_position_30__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227_adj_5839), 
            .I2(VCC_net), .I3(n59220), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_9 (.CI(n59220), .I0(n1227_adj_5839), 
            .I1(VCC_net), .CO(n59221));
    SB_LUT4 encoder0_position_30__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228_adj_5840), 
            .I2(VCC_net), .I3(n59219), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_8 (.CI(n59219), .I0(n1228_adj_5840), 
            .I1(VCC_net), .CO(n59220));
    SB_LUT4 encoder0_position_30__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229_adj_5841), 
            .I2(GND_net), .I3(n59218), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_7 (.CI(n59218), .I0(n1229_adj_5841), 
            .I1(GND_net), .CO(n59219));
    SB_LUT4 mux_243_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_91[14]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230_adj_5842), 
            .I2(GND_net), .I3(n59217), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_6 (.CI(n59217), .I0(n1230_adj_5842), 
            .I1(GND_net), .CO(n59218));
    SB_LUT4 encoder0_position_30__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231_adj_5843), 
            .I2(VCC_net), .I3(n59216), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_5 (.CI(n59216), .I0(n1231_adj_5843), 
            .I1(VCC_net), .CO(n59217));
    SB_LUT4 encoder0_position_30__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232_adj_5844), 
            .I2(GND_net), .I3(n59215), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_4 (.CI(n59215), .I0(n1232_adj_5844), 
            .I1(GND_net), .CO(n59216));
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_91[15]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[16]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_91[16]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i62992_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78848));
    defparam i62992_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233_adj_5845), 
            .I2(VCC_net), .I3(n59214), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_3 (.CI(n59214), .I0(n1233_adj_5845), 
            .I1(VCC_net), .CO(n59215));
    SB_LUT4 encoder0_position_30__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n59214));
    SB_LUT4 encoder0_position_30__I_0_add_1637_24_lut (.I0(n78517), .I1(n2412), 
            .I2(VCC_net), .I3(n59612), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n59611), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_11_lut (.I0(n78869), .I1(n1125), 
            .I2(VCC_net), .I3(n59213), .O(n1224_adj_5836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1637_23 (.CI(n59611), .I0(n2413), 
            .I1(VCC_net), .CO(n59612));
    SB_LUT4 encoder0_position_30__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n59212), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_10 (.CI(n59212), .I0(n1126), 
            .I1(VCC_net), .CO(n59213));
    SB_LUT4 encoder0_position_30__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n59610), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n59211), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_9 (.CI(n59211), .I0(n1127), 
            .I1(VCC_net), .CO(n59212));
    SB_CARRY encoder0_position_30__I_0_add_1637_22 (.CI(n59610), .I0(n2414), 
            .I1(VCC_net), .CO(n59611));
    SB_LUT4 i63061_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78917));
    defparam i63061_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n59210), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_8 (.CI(n59210), .I0(n1128), 
            .I1(VCC_net), .CO(n59211));
    SB_LUT4 encoder0_position_30__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n59609), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n59209), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_7 (.CI(n59209), .I0(n1129), 
            .I1(GND_net), .CO(n59210));
    SB_LUT4 i63013_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78869));
    defparam i63013_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_21 (.CI(n59609), .I0(n2415), 
            .I1(VCC_net), .CO(n59610));
    SB_LUT4 encoder0_position_30__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n59208), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i63074_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78930));
    defparam i63074_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_766_6 (.CI(n59208), .I0(n1130), 
            .I1(GND_net), .CO(n59209));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5906));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n59608), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n59207), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_5 (.CI(n59207), .I0(n1131), 
            .I1(VCC_net), .CO(n59208));
    SB_LUT4 i1_2_lut_4_lut_adj_1915 (.I0(commutation_state[0]), .I1(n4_adj_5966), 
            .I2(commutation_state_prev[0]), .I3(n44559), .O(n28174));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_1915.LUT_INIT = 16'hffde;
    SB_LUT4 i31353_3_lut (.I0(n948), .I1(n2332), .I2(n2333), .I3(GND_net), 
            .O(n45448));
    defparam i31353_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_30__I_0_add_1637_20 (.CI(n59608), .I0(n2416), 
            .I1(VCC_net), .CO(n59609));
    SB_LUT4 encoder0_position_30__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n59206), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_4 (.CI(n59206), .I0(n1132), 
            .I1(GND_net), .CO(n59207));
    SB_LUT4 encoder0_position_30__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n59607), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n59205), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_3 (.CI(n59205), .I0(n1133), 
            .I1(VCC_net), .CO(n59206));
    SB_CARRY encoder0_position_30__I_0_add_1637_19 (.CI(n59607), .I0(n2417), 
            .I1(VCC_net), .CO(n59608));
    SB_LUT4 encoder0_position_30__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n59205));
    SB_LUT4 encoder0_position_30__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n59606), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n59204), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n59203), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_18 (.CI(n59606), .I0(n2418), 
            .I1(VCC_net), .CO(n59607));
    SB_CARRY encoder0_position_30__I_0_add_699_9 (.CI(n59203), .I0(n1027), 
            .I1(VCC_net), .CO(n59204));
    SB_LUT4 encoder0_position_30__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n59202), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n59605), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_8 (.CI(n59202), .I0(n1028), 
            .I1(VCC_net), .CO(n59203));
    SB_LUT4 encoder0_position_30__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n59201), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1916 (.I0(n66979), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[10] [0]), .I3(n67361), .O(n10_adj_5960));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1916.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_30__I_0_add_1637_17 (.CI(n59605), .I0(n2419), 
            .I1(VCC_net), .CO(n59606));
    SB_CARRY encoder0_position_30__I_0_add_699_7 (.CI(n59201), .I0(n1029), 
            .I1(GND_net), .CO(n59202));
    SB_LUT4 encoder0_position_30__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n59200), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n59604), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5905));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5904));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut_adj_1917 (.I0(n30_adj_5912), .I1(n10_adj_5960), .I2(\data_out_frame[11] [7]), 
            .I3(GND_net), .O(n25421));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_adj_1917.LUT_INIT = 16'h9696;
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n58885), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n79582_bdd_4_lut (.I0(n79582), .I1(duty[7]), .I2(n4923), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n79582_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_699_6 (.CI(n59200), .I0(n1030), 
            .I1(GND_net), .CO(n59201));
    SB_LUT4 encoder0_position_30__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n59199), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_5 (.CI(n59199), .I0(n1031), 
            .I1(VCC_net), .CO(n59200));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5903));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5902));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5901));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5900));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_16 (.CI(n59604), .I0(n2420), 
            .I1(VCC_net), .CO(n59605));
    SB_LUT4 encoder0_position_30__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n59603), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_15 (.CI(n59603), .I0(n2421), 
            .I1(VCC_net), .CO(n59604));
    SB_LUT4 encoder0_position_30__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n59602), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_14 (.CI(n59602), .I0(n2422), 
            .I1(VCC_net), .CO(n59603));
    SB_LUT4 encoder0_position_30__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n59601), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_13 (.CI(n59601), .I0(n2423), 
            .I1(VCC_net), .CO(n59602));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5899));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n59600), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n59198), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_4 (.CI(n59198), .I0(n1032), 
            .I1(GND_net), .CO(n59199));
    SB_LUT4 encoder0_position_30__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n59197), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_12 (.CI(n59600), .I0(n2424), 
            .I1(VCC_net), .CO(n59601));
    SB_LUT4 encoder0_position_30__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n59599), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_11 (.CI(n59599), .I0(n2425), 
            .I1(VCC_net), .CO(n59600));
    SB_LUT4 encoder0_position_30__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n59598), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_10 (.CI(n59598), .I0(n2426), 
            .I1(VCC_net), .CO(n59599));
    SB_LUT4 encoder0_position_30__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n59597), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_9 (.CI(n59597), .I0(n2427), 
            .I1(VCC_net), .CO(n59598));
    SB_CARRY encoder0_position_30__I_0_add_699_3 (.CI(n59197), .I0(n1033), 
            .I1(VCC_net), .CO(n59198));
    SB_LUT4 encoder0_position_30__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n59197));
    SB_LUT4 encoder0_position_30__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n59596), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15229_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5966), 
            .I2(commutation_state_prev[0]), .I3(n44559), .O(n29438));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i15229_2_lut_4_lut.LUT_INIT = 16'h00de;
    SB_CARRY encoder0_position_30__I_0_add_1637_8 (.CI(n59596), .I0(n2428), 
            .I1(VCC_net), .CO(n59597));
    SB_LUT4 encoder0_position_30__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n59595), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n59196), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n59195), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_7 (.CI(n59595), .I0(n2429), 
            .I1(GND_net), .CO(n59596));
    SB_LUT4 encoder0_position_30__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n59594), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_8 (.CI(n59195), .I0(n928), 
            .I1(VCC_net), .CO(n59196));
    SB_LUT4 encoder0_position_30__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n59194), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_6 (.CI(n59594), .I0(n2430), 
            .I1(GND_net), .CO(n59595));
    SB_LUT4 encoder0_position_30__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n59593), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_7 (.CI(n59194), .I0(n929), 
            .I1(GND_net), .CO(n59195));
    SB_LUT4 encoder0_position_30__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n59193), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_5 (.CI(n59593), .I0(n2431), 
            .I1(VCC_net), .CO(n59594));
    SB_LUT4 encoder0_position_30__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n59592), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_4 (.CI(n59592), .I0(n2432), 
            .I1(GND_net), .CO(n59593));
    SB_LUT4 encoder0_position_30__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n59591), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_3 (.CI(n59591), .I0(n2433), 
            .I1(VCC_net), .CO(n59592));
    SB_LUT4 encoder0_position_30__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_6 (.CI(n59193), .I0(n930), 
            .I1(GND_net), .CO(n59194));
    SB_LUT4 encoder0_position_30__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n59192), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n59591));
    SB_CARRY encoder0_position_30__I_0_add_632_5 (.CI(n59192), .I0(n931), 
            .I1(VCC_net), .CO(n59193));
    SB_LUT4 encoder0_position_30__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n59191), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [5]), 
            .I2(n26475), .I3(\data_out_frame[16] [1]), .O(n26311));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_30__I_0_add_632_4 (.CI(n59191), .I0(n932), 
            .I1(GND_net), .CO(n59192));
    SB_LUT4 encoder0_position_30__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n59190), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11851_bdd_4_lut_63641 (.I0(n11851), .I1(current[6]), .I2(duty[9]), 
            .I3(n11849), .O(n79576));
    defparam n11851_bdd_4_lut_63641.LUT_INIT = 16'he4aa;
    SB_LUT4 n79576_bdd_4_lut (.I0(n79576), .I1(duty[6]), .I2(n4924), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n79576_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_632_3 (.CI(n59190), .I0(n933), 
            .I1(VCC_net), .CO(n59191));
    SB_LUT4 encoder0_position_30__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11851_bdd_4_lut_63636 (.I0(n11851), .I1(current[5]), .I2(duty[8]), 
            .I3(n11849), .O(n79570));
    defparam n11851_bdd_4_lut_63636.LUT_INIT = 16'he4aa;
    SB_LUT4 n79570_bdd_4_lut (.I0(n79570), .I1(duty[5]), .I2(n4925), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n79570_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n59190));
    SB_LUT4 encoder0_position_30__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n59189), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n59188), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_7 (.CI(n59188), .I0(n829), 
            .I1(GND_net), .CO(n59189));
    SB_LUT4 encoder0_position_30__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n59187), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_6 (.CI(n59187), .I0(n830), 
            .I1(GND_net), .CO(n59188));
    SB_LUT4 encoder0_position_30__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n59186), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_5 (.CI(n59186), .I0(n831), 
            .I1(VCC_net), .CO(n59187));
    SB_LUT4 i1_4_lut_adj_1918 (.I0(n2318), .I1(n2319), .I2(n70848), .I3(n70846), 
            .O(n70854));
    defparam i1_4_lut_adj_1918.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n59185), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_4 (.CI(n59185), .I0(n832), 
            .I1(GND_net), .CO(n59186));
    SB_LUT4 encoder0_position_30__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n59184), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_3 (.CI(n59184), .I0(n833), 
            .I1(VCC_net), .CO(n59185));
    SB_LUT4 n11851_bdd_4_lut_63631 (.I0(n11851), .I1(current[4]), .I2(duty[7]), 
            .I3(n11849), .O(n79564));
    defparam n11851_bdd_4_lut_63631.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n59184));
    SB_LUT4 n79564_bdd_4_lut (.I0(n79564), .I1(duty[4]), .I2(n4926), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n79564_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_2584_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n59183), 
            .O(n7756)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2584_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n59182), 
            .O(n7757)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n65060));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5898));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2584_6 (.CI(n59182), .I0(n622), .I1(GND_net), .CO(n59183));
    SB_LUT4 add_2584_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n59181), 
            .O(n7758)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2584_5 (.CI(n59181), .I0(n623), .I1(VCC_net), .CO(n59182));
    SB_LUT4 add_2584_4_lut (.I0(GND_net), .I1(n291_adj_5806), .I2(GND_net), 
            .I3(n59180), .O(n7759)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11851_bdd_4_lut_63626 (.I0(n11851), .I1(current[3]), .I2(duty[6]), 
            .I3(n11849), .O(n79558));
    defparam n11851_bdd_4_lut_63626.LUT_INIT = 16'he4aa;
    SB_CARRY add_2584_4 (.CI(n59180), .I0(n291_adj_5806), .I1(GND_net), 
            .CO(n59181));
    SB_LUT4 add_2584_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n59179), 
            .O(n7760)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2584_3 (.CI(n59179), .I0(n625), .I1(VCC_net), .CO(n59180));
    SB_LUT4 add_2584_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7761)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2584_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n59179));
    SB_LUT4 i15744_3_lut_4_lut (.I0(n1784), .I1(b_prev_adj_5797), .I2(a_new_adj_6010[1]), 
            .I3(position_31__N_3836_adj_5799), .O(n29958));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15744_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5804));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5805));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1919 (.I0(n2329), .I1(n45448), .I2(n2330), .I3(n2331), 
            .O(n68498));
    defparam i1_4_lut_adj_1919.LUT_INIT = 16'ha080;
    SB_LUT4 i15952_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n66866), 
            .I3(GND_net), .O(n30166));   // verilog/coms.v(130[12] 305[6])
    defparam i15952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5897));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28888_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[7]));
    defparam i28888_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5896));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1920 (.I0(n347), .I1(Ki[1]), .I2(GND_net), .I3(GND_net), 
            .O(n110));
    defparam i1_2_lut_adj_1920.LUT_INIT = 16'h8888;
    SB_LUT4 mux_243_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_91[7]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i969_3_lut (.I0(n1422), .I1(n1489), 
            .I2(n1455), .I3(GND_net), .O(n1521));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n79558_bdd_4_lut (.I0(n79558), .I1(duty[3]), .I2(n4927), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n79558_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5895));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5894));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4978_4_lut (.I0(n25771), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5856));
    defparam i4978_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut (.I0(n24_adj_5856), .I1(delay_counter[14]), .I2(delay_counter[12]), 
            .I3(delay_counter[13]), .O(n69799));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1921 (.I0(n69799), .I1(delay_counter[18]), .I2(n25773), 
            .I3(GND_net), .O(n69558));
    defparam i2_3_lut_adj_1921.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5893));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1570_23_lut (.I0(n78688), .I1(n2313), 
            .I2(VCC_net), .I3(n59549), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n59548), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5892));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_22 (.CI(n59548), .I0(n2314), 
            .I1(VCC_net), .CO(n59549));
    SB_LUT4 encoder0_position_30__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n59547), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5891));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_21 (.CI(n59547), .I0(n2315), 
            .I1(VCC_net), .CO(n59548));
    SB_LUT4 encoder0_position_30__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n59546), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1922 (.I0(delay_counter[23]), .I1(n69558), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7));
    defparam i2_4_lut_adj_1922.LUT_INIT = 16'heaaa;
    SB_CARRY encoder0_position_30__I_0_add_1570_20 (.CI(n59546), .I0(n2316), 
            .I1(VCC_net), .CO(n59547));
    SB_LUT4 encoder0_position_30__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n59545), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1923 (.I0(n7), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n25776), .O(n62));
    defparam i4_4_lut_adj_1923.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5917));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1924 (.I0(delay_counter[28]), .I1(n12_adj_5917), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n25776));
    defparam i6_4_lut_adj_1924.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1925 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n25773));
    defparam i2_3_lut_adj_1925.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5890));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_19 (.CI(n59545), .I0(n2317), 
            .I1(VCC_net), .CO(n59546));
    SB_LUT4 encoder0_position_30__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n59544), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5889));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5888));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_18 (.CI(n59544), .I0(n2318), 
            .I1(VCC_net), .CO(n59545));
    SB_LUT4 encoder0_position_30__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n59543), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1570_17 (.CI(n59543), .I0(n2319), 
            .I1(VCC_net), .CO(n59544));
    SB_LUT4 encoder0_position_30__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n59542), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1926 (.I0(delay_counter[5]), .I1(delay_counter[6]), 
            .I2(delay_counter[1]), .I3(delay_counter[2]), .O(n69884));
    defparam i3_4_lut_adj_1926.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1927 (.I0(n69884), .I1(delay_counter[8]), .I2(delay_counter[4]), 
            .I3(delay_counter[7]), .O(n10_adj_5939));
    defparam i4_4_lut_adj_1927.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1928 (.I0(delay_counter[3]), .I1(n10_adj_5939), 
            .I2(delay_counter[0]), .I3(GND_net), .O(n25771));
    defparam i5_3_lut_adj_1928.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1929 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5742));
    defparam i1_2_lut_adj_1929.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1930 (.I0(delay_counter[9]), .I1(n4_adj_5742), 
            .I2(delay_counter[10]), .I3(n25771), .O(n69651));
    defparam i2_4_lut_adj_1930.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1931 (.I0(n69651), .I1(n25773), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n69831));
    defparam i2_4_lut_adj_1931.LUT_INIT = 16'hffec;
    SB_CARRY encoder0_position_30__I_0_add_1570_16 (.CI(n59542), .I0(n2320), 
            .I1(VCC_net), .CO(n59543));
    SB_LUT4 encoder0_position_30__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n59541), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_15 (.CI(n59541), .I0(n2321), 
            .I1(VCC_net), .CO(n59542));
    SB_LUT4 encoder0_position_30__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n59540), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5887));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5886));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5907));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1932 (.I0(delay_counter[22]), .I1(n69831), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5908));
    defparam i2_4_lut_adj_1932.LUT_INIT = 16'ha8a0;
    SB_LUT4 i30714_4_lut (.I0(n7_adj_5908), .I1(delay_counter[31]), .I2(n25776), 
            .I3(n8_adj_5907), .O(n1319));   // verilog/TinyFPGA_B.v(380[14:38])
    defparam i30714_4_lut.LUT_INIT = 16'h3230;
    SB_CARRY encoder0_position_30__I_0_add_1570_14 (.CI(n59540), .I0(n2322), 
            .I1(VCC_net), .CO(n59541));
    SB_LUT4 encoder0_position_30__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n59539), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_13 (.CI(n59539), .I0(n2323), 
            .I1(VCC_net), .CO(n59540));
    SB_LUT4 encoder0_position_30__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n59538), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_12 (.CI(n59538), .I0(n2324), 
            .I1(VCC_net), .CO(n59539));
    SB_LUT4 encoder0_position_30__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n59537), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11851_bdd_4_lut_63621 (.I0(n11851), .I1(current[2]), .I2(duty[5]), 
            .I3(n11849), .O(n79552));
    defparam n11851_bdd_4_lut_63621.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1237_3_lut (.I0(n1818), .I1(n1885), 
            .I2(n1851), .I3(GND_net), .O(n1917));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5885));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_11 (.CI(n59537), .I0(n2325), 
            .I1(VCC_net), .CO(n59538));
    SB_LUT4 encoder0_position_30__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n59536), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_10 (.CI(n59536), .I0(n2326), 
            .I1(VCC_net), .CO(n59537));
    SB_LUT4 encoder0_position_30__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n59535), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_9 (.CI(n59535), .I0(n2327), 
            .I1(VCC_net), .CO(n59536));
    SB_LUT4 encoder0_position_30__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n59534), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5884));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_8 (.CI(n59534), .I0(n2328), 
            .I1(VCC_net), .CO(n59535));
    SB_LUT4 i15742_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_6047[1]), 
            .I2(r_SM_Main_adj_6047[2]), .I3(n6_adj_5955), .O(n29956));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i15742_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 encoder0_position_30__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n59533), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_7 (.CI(n59533), .I0(n2329), 
            .I1(GND_net), .CO(n59534));
    SB_LUT4 encoder0_position_30__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n59532), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_6 (.CI(n59532), .I0(n2330), 
            .I1(GND_net), .CO(n59533));
    SB_LUT4 n79552_bdd_4_lut (.I0(n79552), .I1(duty[2]), .I2(n4928), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n79552_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16265_4_lut_4_lut (.I0(n28194), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n30479));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16265_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 encoder0_position_30__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n59531), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_5 (.CI(n59531), .I0(n2331), 
            .I1(VCC_net), .CO(n59532));
    SB_LUT4 encoder0_position_30__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n59530), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_4 (.CI(n59530), .I0(n2332), 
            .I1(GND_net), .CO(n59531));
    SB_LUT4 encoder0_position_30__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n59529), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_3 (.CI(n59529), .I0(n2333), 
            .I1(VCC_net), .CO(n59530));
    SB_LUT4 encoder0_position_30__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1933 (.I0(ID[4]), .I1(ID[7]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_5940));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i6_4_lut_adj_1933.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1934 (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5941));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i5_4_lut_adj_1934.LUT_INIT = 16'hfffe;
    SB_LUT4 i30486_4_lut (.I0(n13_adj_5941), .I1(n70662), .I2(n14_adj_5940), 
            .I3(n34_adj_5961), .O(n44574));
    defparam i30486_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 i16808_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n31022));   // verilog/coms.v(130[12] 305[6])
    defparam i16808_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30709_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(366[12:35])
    defparam i30709_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5883));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5882));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n59529));
    SB_LUT4 i14964_4_lut (.I0(n28130), .I1(n1319), .I2(n75123), .I3(n44675), 
            .O(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i14964_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 mux_3812_i13_3_lut (.I0(encoder0_position[12]), .I1(n20_adj_5729), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5881));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5880));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_91[17]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5879));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5878));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5877));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5876));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1503_22_lut (.I0(GND_net), .I1(n2214), 
            .I2(VCC_net), .I3(n59509), .O(n2281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n59508), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_243_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_91[18]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i19_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_30__I_0_add_1503_21 (.CI(n59508), .I0(n2215), 
            .I1(VCC_net), .CO(n59509));
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28130), 
            .D(n1239), .R(n29178));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n59507), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1935 (.I0(n2316), .I1(n68498), .I2(n2317), .I3(n70854), 
            .O(n70860));
    defparam i1_4_lut_adj_1935.LUT_INIT = 16'hfffe;
    SB_LUT4 i62835_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n70860), 
            .O(n2346));
    defparam i62835_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1503_20 (.CI(n59507), .I0(n2216), 
            .I1(VCC_net), .CO(n59508));
    SB_LUT4 encoder0_position_30__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n59506), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_19 (.CI(n59506), .I0(n2217), 
            .I1(VCC_net), .CO(n59507));
    SB_LUT4 n11851_bdd_4_lut_63616 (.I0(n11851), .I1(current[1]), .I2(duty[4]), 
            .I3(n11849), .O(n79546));
    defparam n11851_bdd_4_lut_63616.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n59505), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_18 (.CI(n59505), .I0(n2218), 
            .I1(VCC_net), .CO(n59506));
    SB_LUT4 encoder0_position_30__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n59504), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_17 (.CI(n59504), .I0(n2219), 
            .I1(VCC_net), .CO(n59505));
    SB_LUT4 encoder0_position_30__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n59503), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_16 (.CI(n59503), .I0(n2220), 
            .I1(VCC_net), .CO(n59504));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n59502), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1503_15 (.CI(n59502), .I0(n2221), 
            .I1(VCC_net), .CO(n59503));
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position[25]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position[24]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n28051), .D(GHC_N_391), 
            .R(n29155));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n59501), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n28051), .D(GHB_N_377), 
            .R(n29155));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n28051), .D(GHA_N_355), 
            .R(n29155));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5970), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n28051), .D(GLA_N_372), 
            .R(n29155));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 mux_243_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_91[19]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i20_3_lut.LUT_INIT = 16'h3535;
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n28051), .D(GLB_N_386), 
            .R(n29155));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n28051), .D(GLC_N_400), 
            .R(n29155));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_30__I_0_add_1503_14 (.CI(n59501), .I0(n2222), 
            .I1(VCC_net), .CO(n59502));
    GND i1 (.Y(GND_net));
    SB_LUT4 encoder0_position_30__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n59500), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_13 (.CI(n59500), .I0(n2223), 
            .I1(VCC_net), .CO(n59501));
    SB_LUT4 encoder0_position_30__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n59499), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_12 (.CI(n59499), .I0(n2224), 
            .I1(VCC_net), .CO(n59500));
    SB_LUT4 encoder0_position_30__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n59498), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_11 (.CI(n59498), .I0(n2225), 
            .I1(VCC_net), .CO(n59499));
    SB_LUT4 encoder0_position_30__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n59497), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_10 (.CI(n59497), .I0(n2226), 
            .I1(VCC_net), .CO(n59498));
    SB_LUT4 encoder0_position_30__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n59496), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_9 (.CI(n59496), .I0(n2227), 
            .I1(VCC_net), .CO(n59497));
    SB_LUT4 encoder0_position_30__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n59495), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_8 (.CI(n59495), .I0(n2228), 
            .I1(VCC_net), .CO(n59496));
    SB_LUT4 i12_4_lut_adj_1936 (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(n11_adj_5952));
    defparam i12_4_lut_adj_1936.LUT_INIT = 16'h0aca;
    SB_LUT4 i13_3_lut (.I0(encoder0_position_scaled[20]), .I1(n11_adj_5952), 
            .I2(n15_adj_5793), .I3(GND_net), .O(n12_adj_5853));
    defparam i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n59494), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_7 (.CI(n59494), .I0(n2229), 
            .I1(GND_net), .CO(n59495));
    SB_LUT4 encoder0_position_30__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n59493), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_6 (.CI(n59493), .I0(n2230), 
            .I1(GND_net), .CO(n59494));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n59033), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n59492), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_5 (.CI(n59492), .I0(n2231), 
            .I1(VCC_net), .CO(n59493));
    SB_LUT4 encoder0_position_30__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n59491), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_4 (.CI(n59491), .I0(n2232), 
            .I1(GND_net), .CO(n59492));
    SB_LUT4 encoder0_position_30__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n59490), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_3 (.CI(n59490), .I0(n2233), 
            .I1(VCC_net), .CO(n59491));
    SB_LUT4 encoder0_position_30__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n59490));
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_91[21]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i22_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n59033), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n59034));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n59135), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n59134), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n59134), .I0(GND_net), .I1(n2), 
            .CO(n59135));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5712), 
            .I3(n59133), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n59032), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n59133), .I0(GND_net), .I1(n14_adj_5712), 
            .CO(n59134));
    SB_LUT4 mux_243_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_91[22]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1937 (.I0(n347), .I1(Ki[0]), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_5913));
    defparam i1_2_lut_adj_1937.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5713), 
            .I3(n59132), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n59132), .I0(GND_net), .I1(n15_adj_5713), 
            .CO(n59133));
    SB_LUT4 mux_245_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i24_3_lut (.I0(encoder0_position_scaled[23]), .I1(motor_state_23__N_91[23]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i24_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5714), 
            .I3(n59131), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n59032), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n59033));
    SB_LUT4 n79546_bdd_4_lut (.I0(n79546), .I1(duty[1]), .I2(n4929), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n79546_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24), .I3(n59031), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n59131), .I0(GND_net), .I1(n16_adj_5714), 
            .CO(n59132));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5715), 
            .I3(n59130), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1938 (.I0(n2419), .I1(n2422), .I2(n2423), .I3(n2425), 
            .O(n71206));
    defparam i1_4_lut_adj_1938.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n59130), .I0(GND_net), .I1(n17_adj_5715), 
            .CO(n59131));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5716), 
            .I3(n59129), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n59129), .I0(GND_net), .I1(n18_adj_5716), 
            .CO(n59130));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n59031), .I0(encoder0_position_scaled[1]), 
            .I1(n24), .CO(n59032));
    SB_LUT4 mux_245_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[0]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n11851_bdd_4_lut_63611 (.I0(n11851), .I1(current[0]), .I2(duty[3]), 
            .I3(n11849), .O(n79540));
    defparam n11851_bdd_4_lut_63611.LUT_INIT = 16'he4aa;
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n58878), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_243_i1_3_lut (.I0(encoder0_position_scaled[0]), .I1(motor_state_23__N_91[0]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5717), 
            .I3(n59128), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n59128), .I0(GND_net), .I1(n19_adj_5717), 
            .CO(n59129));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5718), 
            .I3(n59127), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n59127), .I0(GND_net), .I1(n20_adj_5718), 
            .CO(n59128));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25), .CO(n59031));
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i2_3_lut (.I0(encoder0_position_scaled[1]), .I1(motor_state_23__N_91[1]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5719), 
            .I3(n59126), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n59126), .I0(GND_net), .I1(n21_adj_5719), 
            .CO(n59127));
    SB_LUT4 mux_243_i3_3_lut (.I0(encoder0_position_scaled[2]), .I1(motor_state_23__N_91[2]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5720), 
            .I3(n59125), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_11 (.CI(n58885), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n58886));
    SB_CARRY unary_minus_16_add_3_5 (.CI(n59125), .I0(GND_net), .I1(n22_adj_5720), 
            .CO(n59126));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5721), 
            .I3(n59124), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5723));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n59124), .I0(GND_net), .I1(n23_adj_5721), 
            .CO(n59125));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5722), 
            .I3(n59123), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n59123), .I0(GND_net), .I1(n24_adj_5722), 
            .CO(n59124));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n45282), .I1(GND_net), .I2(n25_adj_5723), 
            .I3(VCC_net), .O(n75098)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1436_21_lut (.I0(n78778), .I1(n2115), 
            .I2(VCC_net), .I3(n59463), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5722));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n59462), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5723), 
            .CO(n59123));
    SB_CARRY encoder0_position_30__I_0_add_1436_20 (.CI(n59462), .I0(n2116), 
            .I1(VCC_net), .CO(n59463));
    SB_LUT4 encoder0_position_30__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n59461), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_19 (.CI(n59461), .I0(n2117), 
            .I1(VCC_net), .CO(n59462));
    SB_LUT4 encoder0_position_30__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n59460), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_18 (.CI(n59460), .I0(n2118), 
            .I1(VCC_net), .CO(n59461));
    SB_LUT4 encoder0_position_30__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n59459), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n79540_bdd_4_lut (.I0(n79540), .I1(duty[0]), .I2(n4930), .I3(n11849), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n79540_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1436_17 (.CI(n59459), .I0(n2119), 
            .I1(VCC_net), .CO(n59460));
    SB_LUT4 encoder0_position_30__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n59458), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_16 (.CI(n59458), .I0(n2120), 
            .I1(VCC_net), .CO(n59459));
    SB_LUT4 encoder0_position_30__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n59457), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_15 (.CI(n59457), .I0(n2121), 
            .I1(VCC_net), .CO(n59458));
    SB_LUT4 encoder0_position_30__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n59456), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_14 (.CI(n59456), .I0(n2122), 
            .I1(VCC_net), .CO(n59457));
    SB_LUT4 encoder0_position_30__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n59455), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_13 (.CI(n59455), .I0(n2123), 
            .I1(VCC_net), .CO(n59456));
    SB_LUT4 encoder0_position_30__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n59454), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_12 (.CI(n59454), .I0(n2124), 
            .I1(VCC_net), .CO(n59455));
    SB_LUT4 encoder0_position_30__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n59453), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_11 (.CI(n59453), .I0(n2125), 
            .I1(VCC_net), .CO(n59454));
    SB_LUT4 encoder0_position_30__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n59452), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_10 (.CI(n59452), .I0(n2126), 
            .I1(VCC_net), .CO(n59453));
    SB_LUT4 encoder0_position_30__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n59451), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_9 (.CI(n59451), .I0(n2127), 
            .I1(VCC_net), .CO(n59452));
    SB_LUT4 encoder0_position_30__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n59450), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_8 (.CI(n59450), .I0(n2128), 
            .I1(VCC_net), .CO(n59451));
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5721));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n59449), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(n16_adj_5786));
    defparam i17_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1436_7 (.CI(n59449), .I0(n2129), 
            .I1(GND_net), .CO(n59450));
    SB_LUT4 encoder0_position_30__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n59448), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_6 (.CI(n59448), .I0(n2130), 
            .I1(GND_net), .CO(n59449));
    SB_LUT4 encoder0_position_30__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n59447), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18_3_lut (.I0(encoder0_position_scaled[3]), .I1(n16_adj_5786), 
            .I2(n15_adj_5793), .I3(GND_net), .O(n17_adj_5954));
    defparam i18_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_30__I_0_add_1436_5 (.CI(n59447), .I0(n2131), 
            .I1(VCC_net), .CO(n59448));
    SB_LUT4 encoder0_position_30__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n59446), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_4 (.CI(n59446), .I0(n2132), 
            .I1(GND_net), .CO(n59447));
    SB_LUT4 encoder0_position_30__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n59445), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_3 (.CI(n59445), .I0(n2133), 
            .I1(VCC_net), .CO(n59446));
    SB_LUT4 encoder0_position_30__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n59445));
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5720));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5719));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5718));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5717));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n58907), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n58906), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51831_3_lut (.I0(n4_adj_5746), .I1(n7758), .I2(n67628), .I3(GND_net), 
            .O(n67631));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5716));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_243_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_91[8]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i9_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_151_32 (.CI(n58906), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n58907));
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5715));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51832_3_lut (.I0(encoder0_position[28]), .I1(n67631), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1369_20_lut (.I0(n78754), .I1(n2016), 
            .I2(VCC_net), .I3(n59427), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n59426), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_19 (.CI(n59426), .I0(n2017), 
            .I1(VCC_net), .CO(n59427));
    SB_LUT4 encoder0_position_30__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n59425), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5714));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1369_18 (.CI(n59425), .I0(n2018), 
            .I1(VCC_net), .CO(n59426));
    SB_LUT4 encoder0_position_30__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n59424), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_17 (.CI(n59424), .I0(n2019), 
            .I1(VCC_net), .CO(n59425));
    SB_LUT4 encoder0_position_30__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n59423), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31425_4_lut (.I0(n949), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n45520));
    defparam i31425_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5713));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1369_16 (.CI(n59423), .I0(n2020), 
            .I1(VCC_net), .CO(n59424));
    SB_LUT4 encoder0_position_30__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n59422), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_15 (.CI(n59422), .I0(n2021), 
            .I1(VCC_net), .CO(n59423));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n58905), .O(n1210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n59421), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_14 (.CI(n59421), .I0(n2022), 
            .I1(VCC_net), .CO(n59422));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n59420), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_13 (.CI(n59420), .I0(n2023), 
            .I1(VCC_net), .CO(n59421));
    SB_LUT4 encoder0_position_30__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n59419), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_12 (.CI(n59419), .I0(n2024), 
            .I1(VCC_net), .CO(n59420));
    SB_LUT4 encoder0_position_30__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n59418), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_11 (.CI(n59418), .I0(n2025), 
            .I1(VCC_net), .CO(n59419));
    SB_LUT4 encoder0_position_30__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n59417), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_10 (.CI(n59417), .I0(n2026), 
            .I1(VCC_net), .CO(n59418));
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5712));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n59416), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_9 (.CI(n59416), .I0(n2027), 
            .I1(VCC_net), .CO(n59417));
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n59415), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_8 (.CI(n59415), .I0(n2028), 
            .I1(VCC_net), .CO(n59416));
    SB_LUT4 encoder0_position_30__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n59414), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_7 (.CI(n59414), .I0(n2029), 
            .I1(GND_net), .CO(n59415));
    SB_LUT4 encoder0_position_30__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n59413), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_6 (.CI(n59413), .I0(n2030), 
            .I1(GND_net), .CO(n59414));
    SB_LUT4 encoder0_position_30__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n59412), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_5 (.CI(n59412), .I0(n2031), 
            .I1(VCC_net), .CO(n59413));
    SB_LUT4 encoder0_position_30__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n59411), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_4 (.CI(n59411), .I0(n2032), 
            .I1(GND_net), .CO(n59412));
    SB_LUT4 encoder0_position_30__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n59410), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_3 (.CI(n59410), .I0(n2033), 
            .I1(VCC_net), .CO(n59411));
    SB_LUT4 encoder0_position_30__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n59410));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5876), .I3(n59910), .O(n2_adj_5747)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5877), .I3(n59909), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_32 (.CI(n59909), 
            .I0(GND_net), .I1(n3_adj_5877), .CO(n59910));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5878), .I3(n59908), .O(n4_adj_5746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_31 (.CI(n59908), 
            .I0(GND_net), .I1(n4_adj_5878), .CO(n59909));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5879), .I3(n59907), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_30 (.CI(n59907), 
            .I0(GND_net), .I1(n5_adj_5879), .CO(n59908));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5880), .I3(n59906), .O(n6_adj_5745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_29 (.CI(n59906), 
            .I0(GND_net), .I1(n6_adj_5880), .CO(n59907));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5881), .I3(n59905), .O(n7_adj_5744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_28 (.CI(n59905), 
            .I0(GND_net), .I1(n7_adj_5881), .CO(n59906));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5882), .I3(n59904), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_27 (.CI(n59904), 
            .I0(GND_net), .I1(n8_adj_5882), .CO(n59905));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5883), .I3(n59903), .O(n9_adj_5741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_26 (.CI(n59903), 
            .I0(GND_net), .I1(n9_adj_5883), .CO(n59904));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5884), .I3(n59902), .O(n10_adj_5740)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_25 (.CI(n59902), 
            .I0(GND_net), .I1(n10_adj_5884), .CO(n59903));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5885), .I3(n59901), .O(n11_adj_5739)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_19_lut (.I0(n78373), .I1(n1917), 
            .I2(VCC_net), .I3(n59386), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n59385), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_24 (.CI(n59901), 
            .I0(GND_net), .I1(n11_adj_5885), .CO(n59902));
    SB_CARRY encoder0_position_30__I_0_add_1302_18 (.CI(n59385), .I0(n1918), 
            .I1(VCC_net), .CO(n59386));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5886), .I3(n59900), .O(n12_adj_5737)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n59384), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_17 (.CI(n59384), .I0(n1919), 
            .I1(VCC_net), .CO(n59385));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_23 (.CI(n59900), 
            .I0(GND_net), .I1(n12_adj_5886), .CO(n59901));
    SB_LUT4 encoder0_position_30__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n59383), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5887), .I3(n59899), .O(n13_adj_5736)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_16 (.CI(n59383), .I0(n1920), 
            .I1(VCC_net), .CO(n59384));
    SB_LUT4 encoder0_position_30__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n59382), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_22 (.CI(n59899), 
            .I0(GND_net), .I1(n13_adj_5887), .CO(n59900));
    SB_CARRY encoder0_position_30__I_0_add_1302_15 (.CI(n59382), .I0(n1921), 
            .I1(VCC_net), .CO(n59383));
    SB_LUT4 encoder0_position_30__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n59381), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5888), .I3(n59898), .O(n14_adj_5735)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_14 (.CI(n59381), .I0(n1922), 
            .I1(VCC_net), .CO(n59382));
    SB_LUT4 encoder0_position_30__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n59380), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_21 (.CI(n59898), 
            .I0(GND_net), .I1(n14_adj_5888), .CO(n59899));
    SB_CARRY encoder0_position_30__I_0_add_1302_13 (.CI(n59380), .I0(n1923), 
            .I1(VCC_net), .CO(n59381));
    SB_LUT4 encoder0_position_30__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n59379), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5889), .I3(n59897), .O(n15_adj_5734)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_12 (.CI(n59379), .I0(n1924), 
            .I1(VCC_net), .CO(n59380));
    SB_LUT4 encoder0_position_30__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n59378), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_20 (.CI(n59897), 
            .I0(GND_net), .I1(n15_adj_5889), .CO(n59898));
    SB_CARRY encoder0_position_30__I_0_add_1302_11 (.CI(n59378), .I0(n1925), 
            .I1(VCC_net), .CO(n59379));
    SB_LUT4 encoder0_position_30__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n59377), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5890), .I3(n59896), .O(n16_adj_5733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_10 (.CI(n59377), .I0(n1926), 
            .I1(VCC_net), .CO(n59378));
    SB_LUT4 encoder0_position_30__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n59376), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_19 (.CI(n59896), 
            .I0(GND_net), .I1(n16_adj_5890), .CO(n59897));
    SB_CARRY encoder0_position_30__I_0_add_1302_9 (.CI(n59376), .I0(n1927), 
            .I1(VCC_net), .CO(n59377));
    SB_LUT4 encoder0_position_30__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n59375), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5891), .I3(n59895), .O(n17_adj_5732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_8 (.CI(n59375), .I0(n1928), 
            .I1(VCC_net), .CO(n59376));
    SB_LUT4 encoder0_position_30__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n59374), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_18 (.CI(n59895), 
            .I0(GND_net), .I1(n17_adj_5891), .CO(n59896));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5892), .I3(n59894), .O(n18_adj_5731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_17 (.CI(n59894), 
            .I0(GND_net), .I1(n18_adj_5892), .CO(n59895));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5893), .I3(n59893), .O(n19_adj_5730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_16 (.CI(n59893), 
            .I0(GND_net), .I1(n19_adj_5893), .CO(n59894));
    SB_LUT4 i6661_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6661_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5894), .I3(n59892), .O(n20_adj_5729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_15 (.CI(n59892), 
            .I0(GND_net), .I1(n20_adj_5894), .CO(n59893));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5895), .I3(n59891), .O(n21_adj_5728)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_14 (.CI(n59891), 
            .I0(GND_net), .I1(n21_adj_5895), .CO(n59892));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5896), .I3(n59890), .O(n22_adj_5727)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_7 (.CI(n59374), .I0(n1929), 
            .I1(GND_net), .CO(n59375));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_13 (.CI(n59890), 
            .I0(GND_net), .I1(n22_adj_5896), .CO(n59891));
    SB_LUT4 encoder0_position_30__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n59373), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5897), .I3(n59889), .O(n23_adj_5726)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_6 (.CI(n59373), .I0(n1930), 
            .I1(GND_net), .CO(n59374));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_12 (.CI(n59889), 
            .I0(GND_net), .I1(n23_adj_5897), .CO(n59890));
    SB_LUT4 encoder0_position_30__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n59372), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5898), .I3(n59888), .O(n24_adj_5725)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_5 (.CI(n59372), .I0(n1931), 
            .I1(VCC_net), .CO(n59373));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_11 (.CI(n59888), 
            .I0(GND_net), .I1(n24_adj_5898), .CO(n59889));
    SB_LUT4 encoder0_position_30__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n59371), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5899), .I3(n59887), .O(n25_adj_5724)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_4 (.CI(n59371), .I0(n1932), 
            .I1(GND_net), .CO(n59372));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_10 (.CI(n59887), 
            .I0(GND_net), .I1(n25_adj_5899), .CO(n59888));
    SB_LUT4 encoder0_position_30__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n59370), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5900), .I3(n59886), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_9 (.CI(n59886), 
            .I0(GND_net), .I1(n26_adj_5900), .CO(n59887));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5901), .I3(n59885), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_8 (.CI(n59885), 
            .I0(GND_net), .I1(n27_adj_5901), .CO(n59886));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5902), .I3(n59884), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_7 (.CI(n59884), 
            .I0(GND_net), .I1(n28_adj_5902), .CO(n59885));
    SB_LUT4 i2_2_lut_adj_1939 (.I0(hall2), .I1(commutation_state_7__N_27[2]), 
            .I2(GND_net), .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_adj_1939.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5903), .I3(n59883), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_6 (.CI(n59883), 
            .I0(GND_net), .I1(n29_adj_5903), .CO(n59884));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5904), .I3(n59882), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_3 (.CI(n59370), .I0(n1933), 
            .I1(VCC_net), .CO(n59371));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_5 (.CI(n59882), 
            .I0(GND_net), .I1(n30_adj_5904), .CO(n59883));
    SB_LUT4 encoder0_position_30__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5905), .I3(n59881), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n59370));
    SB_LUT4 i1_3_lut_adj_1940 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1940.LUT_INIT = 16'h1414;
    SB_LUT4 i16659_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n30873));   // verilog/coms.v(130[12] 305[6])
    defparam i16659_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_4 (.CI(n59881), 
            .I0(GND_net), .I1(n31_adj_5905), .CO(n59882));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5906), .I3(n59880), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_3 (.CI(n59880), 
            .I0(GND_net), .I1(n32_adj_5906), .CO(n59881));
    SB_LUT4 i16832_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n31046));   // verilog/coms.v(130[12] 305[6])
    defparam i16832_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n59880));
    SB_LUT4 i6659_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6659_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 add_2634_25_lut (.I0(n78930), .I1(n2_adj_5876), .I2(n1059), 
            .I3(n59879), .O(encoder0_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2634_24_lut (.I0(n78869), .I1(n2_adj_5876), .I2(n1158), 
            .I3(n59878), .O(encoder0_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_24 (.CI(n59878), .I0(n2_adj_5876), .I1(n1158), .CO(n59879));
    SB_LUT4 i14935_2_lut (.I0(n28051), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29155));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14935_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_2634_23_lut (.I0(n78873), .I1(n2_adj_5876), .I2(n1257), 
            .I3(n59877), .O(encoder0_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_23 (.CI(n59877), .I0(n2_adj_5876), .I1(n1257), .CO(n59878));
    SB_LUT4 i62417_4_lut (.I0(commutation_state[1]), .I1(n23188), .I2(dti), 
            .I3(commutation_state[2]), .O(n28051));
    defparam i62417_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 add_2634_22_lut (.I0(n78888), .I1(n2_adj_5876), .I2(n1356), 
            .I3(n59876), .O(encoder0_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_22 (.CI(n59876), .I0(n2_adj_5876), .I1(n1356), .CO(n59877));
    SB_LUT4 i16691_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2874));   // verilog/coms.v(130[12] 305[6])
    defparam i16691_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2634_21_lut (.I0(n78917), .I1(n2_adj_5876), .I2(n1455), 
            .I3(n59875), .O(encoder0_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_21 (.CI(n59875), .I0(n2_adj_5876), .I1(n1455), .CO(n59876));
    SB_LUT4 add_2634_20_lut (.I0(n78848), .I1(n2_adj_5876), .I2(n1554), 
            .I3(n59874), .O(encoder0_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_20 (.CI(n59874), .I0(n2_adj_5876), .I1(n1554), .CO(n59875));
    SB_CARRY add_151_31 (.CI(n58905), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n58906));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n58904), .O(n1211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2634_19_lut (.I0(n78647), .I1(n2_adj_5876), .I2(n1653), 
            .I3(n59873), .O(encoder0_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_19 (.CI(n59873), .I0(n2_adj_5876), .I1(n1653), .CO(n59874));
    SB_LUT4 add_2634_18_lut (.I0(n78377), .I1(n2_adj_5876), .I2(n1752), 
            .I3(n59872), .O(encoder0_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_151_30 (.CI(n58904), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n58905));
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n58903), .O(n1212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2634_18 (.CI(n59872), .I0(n2_adj_5876), .I1(n1752), .CO(n59873));
    SB_LUT4 i31304_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n41637), .O(n45398));
    defparam i31304_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_2634_17_lut (.I0(n78490), .I1(n2_adj_5876), .I2(n1851), 
            .I3(n59871), .O(encoder0_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_17 (.CI(n59871), .I0(n2_adj_5876), .I1(n1851), .CO(n59872));
    SB_LUT4 add_2634_16_lut (.I0(n78373), .I1(n2_adj_5876), .I2(n1950), 
            .I3(n59870), .O(encoder0_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1190_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n58999), .O(n4907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n58884), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_29 (.CI(n58903), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n58904));
    SB_CARRY add_2634_16 (.CI(n59870), .I0(n2_adj_5876), .I1(n1950), .CO(n59871));
    SB_LUT4 add_2634_15_lut (.I0(n78754), .I1(n2_adj_5876), .I2(n2049), 
            .I3(n59869), .O(encoder0_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_15 (.CI(n59869), .I0(n2_adj_5876), .I1(n2049), .CO(n59870));
    SB_LUT4 add_2634_14_lut (.I0(n78778), .I1(n2_adj_5876), .I2(n2148), 
            .I3(n59868), .O(encoder0_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_14 (.CI(n59868), .I0(n2_adj_5876), .I1(n2148), .CO(n59869));
    SB_LUT4 add_2634_13_lut (.I0(n78728), .I1(n2_adj_5876), .I2(n2247), 
            .I3(n59867), .O(encoder0_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_13 (.CI(n59867), .I0(n2_adj_5876), .I1(n2247), .CO(n59868));
    SB_LUT4 add_2634_12_lut (.I0(n78688), .I1(n2_adj_5876), .I2(n2346), 
            .I3(n59866), .O(encoder0_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_12 (.CI(n59866), .I0(n2_adj_5876), .I1(n2346), .CO(n59867));
    SB_LUT4 add_2634_11_lut (.I0(n78517), .I1(n2_adj_5876), .I2(n2445), 
            .I3(n59865), .O(encoder0_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_11 (.CI(n59865), .I0(n2_adj_5876), .I1(n2445), .CO(n59866));
    SB_LUT4 add_2634_10_lut (.I0(n78616), .I1(n2_adj_5876), .I2(n2544), 
            .I3(n59864), .O(encoder0_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_10 (.CI(n59864), .I0(n2_adj_5876), .I1(n2544), .CO(n59865));
    SB_LUT4 add_1190_24_lut (.I0(GND_net), .I1(GND_net), .I2(n12450), 
            .I3(n58998), .O(n4908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1941 (.I0(state[0]), .I1(bit_ctr[3]), .I2(n44741), 
            .I3(bit_ctr[4]), .O(n4));   // verilog/neopixel.v(34[12] 113[6])
    defparam i1_2_lut_4_lut_adj_1941.LUT_INIT = 16'hd555;
    SB_LUT4 add_2634_9_lut (.I0(n78546), .I1(n2_adj_5876), .I2(n2643), 
            .I3(n59863), .O(encoder0_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1190_24 (.CI(n58998), .I0(GND_net), .I1(n12450), .CO(n58999));
    SB_CARRY add_2634_9 (.CI(n59863), .I0(n2_adj_5876), .I1(n2643), .CO(n59864));
    SB_LUT4 add_1190_23_lut (.I0(GND_net), .I1(GND_net), .I2(n12452), 
            .I3(n58997), .O(n4909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_4 (.CI(n58878), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n58879));
    SB_LUT4 add_2634_8_lut (.I0(n78463), .I1(n2_adj_5876), .I2(n2742), 
            .I3(n59862), .O(encoder0_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1190_23 (.CI(n58997), .I0(GND_net), .I1(n12452), .CO(n58998));
    SB_CARRY add_151_10 (.CI(n58884), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n58885));
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n58902), .O(n1213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2634_8 (.CI(n59862), .I0(n2_adj_5876), .I1(n2742), .CO(n59863));
    SB_LUT4 add_1190_22_lut (.I0(GND_net), .I1(GND_net), .I2(n12454), 
            .I3(n58996), .O(n4910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_28 (.CI(n58902), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n58903));
    SB_LUT4 add_2634_7_lut (.I0(n78580), .I1(n2_adj_5876), .I2(n2841), 
            .I3(n59861), .O(encoder0_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1190_22 (.CI(n58996), .I0(GND_net), .I1(n12454), .CO(n58997));
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n58901), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n58883), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2634_7 (.CI(n59861), .I0(n2_adj_5876), .I1(n2841), .CO(n59862));
    SB_LUT4 add_1190_21_lut (.I0(GND_net), .I1(GND_net), .I2(n12456), 
            .I3(n58995), .O(n4911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_27 (.CI(n58901), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n58902));
    SB_LUT4 add_2634_6_lut (.I0(n78612), .I1(n2_adj_5876), .I2(n2940), 
            .I3(n59860), .O(encoder0_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1190_21 (.CI(n58995), .I0(GND_net), .I1(n12456), .CO(n58996));
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n58877), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2634_6 (.CI(n59860), .I0(n2_adj_5876), .I1(n2940), .CO(n59861));
    SB_LUT4 add_1190_20_lut (.I0(GND_net), .I1(GND_net), .I2(n12458), 
            .I3(n58994), .O(n4912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_9 (.CI(n58883), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n58884));
    SB_LUT4 i15513_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n23094), .I3(GND_net), .O(n29727));   // verilog/coms.v(130[12] 305[6])
    defparam i15513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2634_5_lut (.I0(n78937), .I1(n2_adj_5876), .I2(n3039), 
            .I3(n59859), .O(encoder0_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_5 (.CI(n59859), .I0(n2_adj_5876), .I1(n3039), .CO(n59860));
    SB_LUT4 add_2634_4_lut (.I0(n78970), .I1(n2_adj_5876), .I2(n3138), 
            .I3(n59858), .O(encoder0_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_4 (.CI(n59858), .I0(n2_adj_5876), .I1(n3138), .CO(n59859));
    SB_LUT4 add_2634_3_lut (.I0(n79004), .I1(n2_adj_5876), .I2(n3237), 
            .I3(n59857), .O(encoder0_position_scaled_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_3 (.CI(n59857), .I0(n2_adj_5876), .I1(n3237), .CO(n59858));
    SB_LUT4 add_2634_2_lut (.I0(n78351), .I1(n2_adj_5876), .I2(n45484), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_2 (.CI(VCC_net), .I0(n2_adj_5876), .I1(n45484), 
            .CO(n59857));
    SB_LUT4 encoder0_position_30__I_0_add_2173_33_lut (.I0(n79004), .I1(n3204), 
            .I2(VCC_net), .I3(n59856), .O(n72039)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1190_20 (.CI(n58994), .I0(GND_net), .I1(n12458), .CO(n58995));
    SB_LUT4 encoder0_position_30__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n59855), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_19_lut (.I0(GND_net), .I1(GND_net), .I2(n12460), 
            .I3(n58993), .O(n4913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_32 (.CI(n59855), .I0(n3205), 
            .I1(VCC_net), .CO(n59856));
    SB_LUT4 encoder0_position_30__I_0_add_1235_18_lut (.I0(GND_net), .I1(n1818), 
            .I2(VCC_net), .I3(n59354), .O(n1885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_19 (.CI(n58993), .I0(GND_net), .I1(n12460), .CO(n58994));
    SB_LUT4 encoder0_position_30__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n59854), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_18_lut (.I0(GND_net), .I1(GND_net), .I2(n12462), 
            .I3(n58992), .O(n4914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_31 (.CI(n59854), .I0(n3206), 
            .I1(VCC_net), .CO(n59855));
    SB_LUT4 encoder0_position_30__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n59353), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_18 (.CI(n58992), .I0(GND_net), .I1(n12462), .CO(n58993));
    SB_LUT4 encoder0_position_30__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n59853), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_17_lut (.I0(GND_net), .I1(GND_net), .I2(n12464), 
            .I3(n58991), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_30 (.CI(n59853), .I0(n3207), 
            .I1(VCC_net), .CO(n59854));
    SB_CARRY encoder0_position_30__I_0_add_1235_17 (.CI(n59353), .I0(n1819), 
            .I1(VCC_net), .CO(n59354));
    SB_CARRY add_1190_17 (.CI(n58991), .I0(GND_net), .I1(n12464), .CO(n58992));
    SB_LUT4 encoder0_position_30__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n59852), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n59352), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_16_lut (.I0(GND_net), .I1(GND_net), .I2(n12466), 
            .I3(n58990), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n58900), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_26 (.CI(n58900), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n58901));
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(n3476), .I1(n89), .I2(reset), .I3(GND_net), 
            .O(n82));
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_CARRY encoder0_position_30__I_0_add_2173_29 (.CI(n59852), .I0(n3208), 
            .I1(VCC_net), .CO(n59853));
    SB_LUT4 encoder0_position_30__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n59851), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_28 (.CI(n59851), .I0(n3209), 
            .I1(VCC_net), .CO(n59852));
    SB_LUT4 encoder0_position_30__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n59850), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_27 (.CI(n59850), .I0(n3210), 
            .I1(VCC_net), .CO(n59851));
    SB_LUT4 encoder0_position_30__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n59849), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_26 (.CI(n59849), .I0(n3211), 
            .I1(VCC_net), .CO(n59850));
    SB_LUT4 encoder0_position_30__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n59848), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_25 (.CI(n59848), .I0(n3212), 
            .I1(VCC_net), .CO(n59849));
    SB_LUT4 encoder0_position_30__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n59847), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_16 (.CI(n59352), .I0(n1820), 
            .I1(VCC_net), .CO(n59353));
    SB_CARRY add_1190_16 (.CI(n58990), .I0(GND_net), .I1(n12466), .CO(n58991));
    SB_CARRY encoder0_position_30__I_0_add_2173_24 (.CI(n59847), .I0(n3213), 
            .I1(VCC_net), .CO(n59848));
    SB_LUT4 add_1190_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12468), 
            .I3(n58989), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n59846), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n59351), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_15 (.CI(n58989), .I0(GND_net), .I1(n12468), .CO(n58990));
    SB_CARRY encoder0_position_30__I_0_add_2173_23 (.CI(n59846), .I0(n3214), 
            .I1(VCC_net), .CO(n59847));
    SB_LUT4 add_1190_14_lut (.I0(GND_net), .I1(GND_net), .I2(n12470), 
            .I3(n58988), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n59845), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_15 (.CI(n59351), .I0(n1821), 
            .I1(VCC_net), .CO(n59352));
    SB_CARRY add_1190_14 (.CI(n58988), .I0(GND_net), .I1(n12470), .CO(n58989));
    SB_CARRY encoder0_position_30__I_0_add_2173_22 (.CI(n59845), .I0(n3215), 
            .I1(VCC_net), .CO(n59846));
    SB_LUT4 add_1190_13_lut (.I0(GND_net), .I1(GND_net), .I2(n12472), 
            .I3(n58987), .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n59844), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822_adj_5851), 
            .I2(VCC_net), .I3(n59350), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_21 (.CI(n59844), .I0(n3216), 
            .I1(VCC_net), .CO(n59845));
    SB_CARRY add_1190_13 (.CI(n58987), .I0(GND_net), .I1(n12472), .CO(n58988));
    SB_LUT4 encoder0_position_30__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n59843), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_12_lut (.I0(GND_net), .I1(GND_net), .I2(n12474), 
            .I3(n58986), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_20 (.CI(n59843), .I0(n3217), 
            .I1(VCC_net), .CO(n59844));
    SB_LUT4 encoder0_position_30__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n59842), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_19 (.CI(n59842), .I0(n3218), 
            .I1(VCC_net), .CO(n59843));
    SB_LUT4 encoder0_position_30__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n59841), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_18 (.CI(n59841), .I0(n3219), 
            .I1(VCC_net), .CO(n59842));
    SB_LUT4 encoder0_position_30__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n59840), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_17 (.CI(n59840), .I0(n3220), 
            .I1(VCC_net), .CO(n59841));
    SB_LUT4 encoder0_position_30__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n59839), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_14 (.CI(n59350), .I0(n1822_adj_5851), 
            .I1(VCC_net), .CO(n59351));
    SB_CARRY encoder0_position_30__I_0_add_2173_16 (.CI(n59839), .I0(n3221), 
            .I1(VCC_net), .CO(n59840));
    SB_LUT4 encoder0_position_30__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n59349), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_12 (.CI(n58986), .I0(GND_net), .I1(n12474), .CO(n58987));
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n58899), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_25 (.CI(n58899), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n58900));
    SB_LUT4 encoder0_position_30__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n59838), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_11_lut (.I0(GND_net), .I1(GND_net), .I2(n12476), 
            .I3(n58985), .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1942 (.I0(n2424), .I1(n2428), .I2(n2426), .I3(n2427), 
            .O(n71126));
    defparam i1_4_lut_adj_1942.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_2173_15 (.CI(n59838), .I0(n3222), 
            .I1(VCC_net), .CO(n59839));
    SB_CARRY encoder0_position_30__I_0_add_1235_13 (.CI(n59349), .I0(n1823), 
            .I1(VCC_net), .CO(n59350));
    SB_CARRY add_1190_11 (.CI(n58985), .I0(GND_net), .I1(n12476), .CO(n58986));
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n58898), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_24 (.CI(n58898), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n58899));
    SB_LUT4 encoder0_position_30__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n59837), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_10_lut (.I0(GND_net), .I1(GND_net), .I2(n12478), 
            .I3(n58984), .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n58882), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_14 (.CI(n59837), .I0(n3223), 
            .I1(VCC_net), .CO(n59838));
    SB_LUT4 encoder0_position_30__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824_adj_5852), 
            .I2(VCC_net), .I3(n59348), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_10 (.CI(n58984), .I0(GND_net), .I1(n12478), .CO(n58985));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n58897), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n59836), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_13 (.CI(n59836), .I0(n3224), 
            .I1(VCC_net), .CO(n59837));
    SB_CARRY add_151_3 (.CI(n58877), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n58878));
    SB_LUT4 encoder0_position_30__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n59835), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_9_lut (.I0(GND_net), .I1(GND_net), .I2(n12480), .I3(n58983), 
            .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_8 (.CI(n58882), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n58883));
    SB_CARRY add_151_23 (.CI(n58897), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n58898));
    SB_CARRY encoder0_position_30__I_0_add_1235_12 (.CI(n59348), .I0(n1824_adj_5852), 
            .I1(VCC_net), .CO(n59349));
    SB_CARRY encoder0_position_30__I_0_add_2173_12 (.CI(n59835), .I0(n3225), 
            .I1(VCC_net), .CO(n59836));
    SB_LUT4 encoder0_position_30__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n59347), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n58896), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n59834), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_11 (.CI(n59347), .I0(n1825), 
            .I1(VCC_net), .CO(n59348));
    SB_CARRY add_1190_9 (.CI(n58983), .I0(GND_net), .I1(n12480), .CO(n58984));
    SB_CARRY add_151_22 (.CI(n58896), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n58897));
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n58895), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_11 (.CI(n59834), .I0(n3226), 
            .I1(VCC_net), .CO(n59835));
    SB_LUT4 encoder0_position_30__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n59346), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_10 (.CI(n59346), .I0(n1826), 
            .I1(VCC_net), .CO(n59347));
    SB_LUT4 encoder0_position_30__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n59833), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_10 (.CI(n59833), .I0(n3227), 
            .I1(VCC_net), .CO(n59834));
    SB_LUT4 encoder0_position_30__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n59832), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_9 (.CI(n59832), .I0(n3228), 
            .I1(VCC_net), .CO(n59833));
    SB_LUT4 encoder0_position_30__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n59831), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_8 (.CI(n59831), .I0(n3229), 
            .I1(GND_net), .CO(n59832));
    SB_LUT4 encoder0_position_30__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n59830), .O(n75097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_7 (.CI(n59830), .I0(n3230), 
            .I1(GND_net), .CO(n59831));
    SB_LUT4 encoder0_position_30__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n59345), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_9 (.CI(n59345), .I0(n1827), 
            .I1(VCC_net), .CO(n59346));
    SB_LUT4 encoder0_position_30__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n59829), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_6 (.CI(n59829), .I0(n3231), 
            .I1(VCC_net), .CO(n59830));
    SB_LUT4 encoder0_position_30__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n59344), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_5_lut (.I0(n6_adj_5914), .I1(n3232), 
            .I2(GND_net), .I3(n59828), .O(n75094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_30__I_0_add_1235_8 (.CI(n59344), .I0(n1828), 
            .I1(VCC_net), .CO(n59345));
    SB_CARRY encoder0_position_30__I_0_add_2173_5 (.CI(n59828), .I0(n3232), 
            .I1(GND_net), .CO(n59829));
    SB_LUT4 add_1190_8_lut (.I0(GND_net), .I1(GND_net), .I2(n12482), .I3(n58982), 
            .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_4_lut (.I0(n3301), .I1(n3233), 
            .I2(VCC_net), .I3(n59827), .O(n6_adj_5914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n59343), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1943 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n71380));
    defparam i1_2_lut_adj_1943.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_30__I_0_add_2173_4 (.CI(n59827), .I0(n3233), 
            .I1(VCC_net), .CO(n59828));
    SB_LUT4 encoder0_position_30__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n59826), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_7 (.CI(n59343), .I0(n1829), 
            .I1(GND_net), .CO(n59344));
    SB_CARRY encoder0_position_30__I_0_add_2173_3 (.CI(n59826), .I0(n957), 
            .I1(GND_net), .CO(n59827));
    SB_LUT4 encoder0_position_30__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n59342), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_8 (.CI(n58982), .I0(GND_net), .I1(n12482), .CO(n58983));
    SB_CARRY encoder0_position_30__I_0_add_2173_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n59826));
    SB_LUT4 add_1190_7_lut (.I0(GND_net), .I1(GND_net), .I2(n12484), .I3(n58981), 
            .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2106_31_lut (.I0(n78970), .I1(n3105), 
            .I2(VCC_net), .I3(n59825), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1235_6 (.CI(n59342), .I0(n1830), 
            .I1(GND_net), .CO(n59343));
    SB_CARRY add_1190_7 (.CI(n58981), .I0(GND_net), .I1(n12484), .CO(n58982));
    SB_LUT4 encoder0_position_30__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n59824), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_6_lut (.I0(GND_net), .I1(GND_net), .I2(n12486), .I3(n58980), 
            .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_30 (.CI(n59824), .I0(n3106), 
            .I1(VCC_net), .CO(n59825));
    SB_LUT4 i16825_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n31039));   // verilog/coms.v(130[12] 305[6])
    defparam i16825_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n59823), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n59341), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_6 (.CI(n58980), .I0(GND_net), .I1(n12486), .CO(n58981));
    SB_CARRY add_151_21 (.CI(n58895), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n58896));
    SB_CARRY encoder0_position_30__I_0_add_2106_29 (.CI(n59823), .I0(n3107), 
            .I1(VCC_net), .CO(n59824));
    SB_LUT4 add_1190_5_lut (.I0(GND_net), .I1(GND_net), .I2(n12488), .I3(n58979), 
            .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n58894), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n58881), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n59822), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_28 (.CI(n59822), .I0(n3108), 
            .I1(VCC_net), .CO(n59823));
    SB_CARRY encoder0_position_30__I_0_add_1235_5 (.CI(n59341), .I0(n1831), 
            .I1(VCC_net), .CO(n59342));
    SB_LUT4 encoder0_position_30__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n59340), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n59821), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_4 (.CI(n59340), .I0(n1832), 
            .I1(GND_net), .CO(n59341));
    SB_CARRY add_1190_5 (.CI(n58979), .I0(GND_net), .I1(n12488), .CO(n58980));
    SB_CARRY add_151_20 (.CI(n58894), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n58895));
    SB_CARRY encoder0_position_30__I_0_add_2106_27 (.CI(n59821), .I0(n3109), 
            .I1(VCC_net), .CO(n59822));
    SB_LUT4 encoder0_position_30__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n59339), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_3 (.CI(n59339), .I0(n1833), 
            .I1(VCC_net), .CO(n59340));
    SB_LUT4 encoder0_position_30__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n59820), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_26 (.CI(n59820), .I0(n3110), 
            .I1(VCC_net), .CO(n59821));
    SB_CARRY encoder0_position_30__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n59339));
    SB_LUT4 encoder0_position_30__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n59819), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_25 (.CI(n59819), .I0(n3111), 
            .I1(VCC_net), .CO(n59820));
    SB_LUT4 encoder0_position_30__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n59818), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_24 (.CI(n59818), .I0(n3112), 
            .I1(VCC_net), .CO(n59819));
    SB_LUT4 encoder0_position_30__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n59817), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_23 (.CI(n59817), .I0(n3113), 
            .I1(VCC_net), .CO(n59818));
    SB_LUT4 encoder0_position_30__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n59816), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1944 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[12] [5]), .I3(\data_in_frame[12] [6]), .O(n67578));
    defparam i1_2_lut_4_lut_adj_1944.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_30__I_0_add_2106_22 (.CI(n59816), .I0(n3114), 
            .I1(VCC_net), .CO(n59817));
    SB_LUT4 add_1190_4_lut (.I0(GND_net), .I1(GND_net), .I2(n12490), .I3(n58978), 
            .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_4 (.CI(n58978), .I0(GND_net), .I1(n12490), .CO(n58979));
    SB_LUT4 encoder0_position_30__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n59815), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1945 (.I0(n2421), .I1(n71380), .I2(n71126), .I3(n45520), 
            .O(n71130));
    defparam i1_4_lut_adj_1945.LUT_INIT = 16'hfefa;
    SB_CARRY encoder0_position_30__I_0_add_2106_21 (.CI(n59815), .I0(n3115), 
            .I1(VCC_net), .CO(n59816));
    SB_LUT4 encoder0_position_30__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n59814), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[9] [5]), .I3(GND_net), .O(n66979));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n66744));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 add_1190_3_lut (.I0(GND_net), .I1(GND_net), .I2(n12492), .I3(n58977), 
            .O(n4929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_20 (.CI(n59814), .I0(n3116), 
            .I1(VCC_net), .CO(n59815));
    SB_CARRY add_1190_3 (.CI(n58977), .I0(GND_net), .I1(n12492), .CO(n58978));
    SB_LUT4 encoder0_position_30__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n59813), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_2_lut (.I0(GND_net), .I1(GND_net), .I2(n11914), .I3(VCC_net), 
            .O(n4930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_19 (.CI(n59813), .I0(n3117), 
            .I1(VCC_net), .CO(n59814));
    SB_CARRY add_1190_2 (.CI(VCC_net), .I0(GND_net), .I1(n11914), .CO(n58977));
    SB_LUT4 encoder0_position_30__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n59812), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n66703));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226_adj_5838));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2106_18 (.CI(n59812), .I0(n3118), 
            .I1(VCC_net), .CO(n59813));
    SB_LUT4 encoder0_position_30__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n59811), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_17 (.CI(n59811), .I0(n3119), 
            .I1(VCC_net), .CO(n59812));
    SB_LUT4 encoder0_position_30__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n59810), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n29359));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2106_16 (.CI(n59810), .I0(n3120), 
            .I1(VCC_net), .CO(n59811));
    SB_LUT4 encoder0_position_30__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n59809), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_15 (.CI(n59809), .I0(n3121), 
            .I1(VCC_net), .CO(n59810));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1948 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n66700));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1948.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n59808), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_14 (.CI(n59808), .I0(n3122), 
            .I1(VCC_net), .CO(n59809));
    SB_LUT4 encoder0_position_30__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n59807), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_13 (.CI(n59807), .I0(n3123), 
            .I1(VCC_net), .CO(n59808));
    SB_LUT4 encoder0_position_30__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n59806), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_12 (.CI(n59806), .I0(n3124), 
            .I1(VCC_net), .CO(n59807));
    SB_LUT4 encoder0_position_30__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n59805), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n66699));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1168_17_lut (.I0(n78377), .I1(n1719), 
            .I2(VCC_net), .I3(n59318), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2106_11 (.CI(n59805), .I0(n3125), 
            .I1(VCC_net), .CO(n59806));
    SB_LUT4 encoder0_position_30__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n59317), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_16 (.CI(n59317), .I0(n1720), 
            .I1(VCC_net), .CO(n59318));
    SB_LUT4 encoder0_position_30__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n59804), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n59316), .O(n1788_adj_5846)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_15 (.CI(n59316), .I0(n1721), 
            .I1(VCC_net), .CO(n59317));
    SB_CARRY encoder0_position_30__I_0_add_2106_10 (.CI(n59804), .I0(n3126), 
            .I1(VCC_net), .CO(n59805));
    SB_LUT4 encoder0_position_30__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n59315), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1950 (.I0(n2415), .I1(n2416), .I2(n2418), .I3(n71206), 
            .O(n71212));
    defparam i1_4_lut_adj_1950.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1168_14 (.CI(n59315), .I0(n1722), 
            .I1(VCC_net), .CO(n59316));
    SB_LUT4 encoder0_position_30__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n59803), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n59314), .O(n1790_adj_5847)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_13 (.CI(n59314), .I0(n1723), 
            .I1(VCC_net), .CO(n59315));
    SB_CARRY encoder0_position_30__I_0_add_2106_9 (.CI(n59803), .I0(n3127), 
            .I1(VCC_net), .CO(n59804));
    SB_LUT4 encoder0_position_30__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n59313), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n59802), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_12 (.CI(n59313), .I0(n1724), 
            .I1(VCC_net), .CO(n59314));
    SB_CARRY encoder0_position_30__I_0_add_2106_8 (.CI(n59802), .I0(n3128), 
            .I1(VCC_net), .CO(n59803));
    SB_LUT4 encoder0_position_30__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n59312), .O(n1792_adj_5848)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n59801), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_11 (.CI(n59312), .I0(n1725), 
            .I1(VCC_net), .CO(n59313));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n66577));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2106_7 (.CI(n59801), .I0(n3129), 
            .I1(GND_net), .CO(n59802));
    SB_LUT4 encoder0_position_30__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n59311), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n59800), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_10 (.CI(n59311), .I0(n1726), 
            .I1(VCC_net), .CO(n59312));
    SB_CARRY encoder0_position_30__I_0_add_2106_6 (.CI(n59800), .I0(n3130), 
            .I1(GND_net), .CO(n59801));
    SB_LUT4 encoder0_position_30__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n59310), .O(n1794_adj_5849)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n59799), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_9 (.CI(n59310), .I0(n1727), 
            .I1(VCC_net), .CO(n59311));
    SB_CARRY encoder0_position_30__I_0_add_2106_5 (.CI(n59799), .I0(n3131), 
            .I1(VCC_net), .CO(n59800));
    SB_LUT4 encoder0_position_30__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n59309), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_8 (.CI(n59309), .I0(n1728), 
            .I1(VCC_net), .CO(n59310));
    SB_LUT4 encoder0_position_30__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n59798), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n59308), .O(n1796_adj_5850)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15541_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n23094), .I3(GND_net), .O(n29755));   // verilog/coms.v(130[12] 305[6])
    defparam i15541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n66698));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [6]), .I3(\data_out_frame[9] [6]), .O(n67599));   // verilog/coms.v(100[12:26])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_30__I_0_add_1168_7 (.CI(n59308), .I0(n1729), 
            .I1(GND_net), .CO(n59309));
    SB_CARRY encoder0_position_30__I_0_add_2106_4 (.CI(n59798), .I0(n3132), 
            .I1(GND_net), .CO(n59799));
    SB_LUT4 encoder0_position_30__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n59307), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_6 (.CI(n59307), .I0(n1730), 
            .I1(GND_net), .CO(n59308));
    SB_LUT4 encoder0_position_30__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n59797), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n59306), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_3 (.CI(n59797), .I0(n3133), 
            .I1(VCC_net), .CO(n59798));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n66697));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n58893), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_5 (.CI(n59306), .I0(n1731), 
            .I1(VCC_net), .CO(n59307));
    SB_LUT4 encoder0_position_30__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n59305), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n59797));
    SB_CARRY encoder0_position_30__I_0_add_1168_4 (.CI(n59305), .I0(n1732), 
            .I1(GND_net), .CO(n59306));
    SB_LUT4 encoder0_position_30__I_0_add_2039_30_lut (.I0(n78937), .I1(n3006), 
            .I2(VCC_net), .I3(n59796), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n59304), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_3 (.CI(n59304), .I0(n1733), 
            .I1(VCC_net), .CO(n59305));
    SB_LUT4 encoder0_position_30__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n59795), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n59304));
    SB_CARRY encoder0_position_30__I_0_add_2039_29 (.CI(n59795), .I0(n3007), 
            .I1(VCC_net), .CO(n59796));
    SB_LUT4 encoder0_position_30__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n59794), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_28 (.CI(n59794), .I0(n3008), 
            .I1(VCC_net), .CO(n59795));
    SB_LUT4 encoder0_position_30__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n59793), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_19 (.CI(n58893), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n58894));
    SB_CARRY encoder0_position_30__I_0_add_2039_27 (.CI(n59793), .I0(n3009), 
            .I1(VCC_net), .CO(n59794));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n66696));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n59792), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_26 (.CI(n59792), .I0(n3010), 
            .I1(VCC_net), .CO(n59793));
    SB_LUT4 encoder0_position_30__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n59791), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n66695));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2039_25 (.CI(n59791), .I0(n3011), 
            .I1(VCC_net), .CO(n59792));
    SB_LUT4 encoder0_position_30__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n59790), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_24 (.CI(n59790), .I0(n3012), 
            .I1(VCC_net), .CO(n59791));
    SB_LUT4 encoder0_position_30__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n59789), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_23 (.CI(n59789), .I0(n3013), 
            .I1(VCC_net), .CO(n59790));
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 encoder0_position_30__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n59788), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_22 (.CI(n59788), .I0(n3014), 
            .I1(VCC_net), .CO(n59789));
    SB_LUT4 encoder0_position_30__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n59787), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n66694));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2039_21 (.CI(n59787), .I0(n3015), 
            .I1(VCC_net), .CO(n59788));
    SB_LUT4 encoder0_position_30__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n59786), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_7 (.CI(n58881), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n58882));
    SB_CARRY encoder0_position_30__I_0_add_2039_20 (.CI(n59786), .I0(n3016), 
            .I1(VCC_net), .CO(n59787));
    SB_LUT4 encoder0_position_30__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n59785), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_19 (.CI(n59785), .I0(n3017), 
            .I1(VCC_net), .CO(n59786));
    SB_LUT4 encoder0_position_30__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n59784), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n27_adj_5910));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2039_18 (.CI(n59784), .I0(n3018), 
            .I1(VCC_net), .CO(n59785));
    SB_LUT4 encoder0_position_30__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n59783), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_17 (.CI(n59783), .I0(n3019), 
            .I1(VCC_net), .CO(n59784));
    SB_LUT4 encoder0_position_30__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n59782), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_16 (.CI(n59782), .I0(n3020), 
            .I1(VCC_net), .CO(n59783));
    SB_LUT4 encoder0_position_30__I_0_add_1101_16_lut (.I0(n78647), .I1(n1620), 
            .I2(VCC_net), .I3(n59290), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n58892), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n59289), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n59781), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_15 (.CI(n59289), .I0(n1621), 
            .I1(VCC_net), .CO(n59290));
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_18 (.CI(n58892), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n58893));
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n58880), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n59288), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_15 (.CI(n59781), .I0(n3021), 
            .I1(VCC_net), .CO(n59782));
    SB_CARRY encoder0_position_30__I_0_add_1101_14 (.CI(n59288), .I0(n1622), 
            .I1(VCC_net), .CO(n59289));
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n58891), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_17 (.CI(n58891), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n58892));
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n58890), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n59287), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n59780), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_13 (.CI(n59287), .I0(n1623), 
            .I1(VCC_net), .CO(n59288));
    SB_CARRY add_151_16 (.CI(n58890), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n58891));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n58889), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n59286), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1505_3_lut (.I0(n2214), .I1(n2281), 
            .I2(n2247), .I3(GND_net), .O(n2313));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1505_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2039_14 (.CI(n59780), .I0(n3022), 
            .I1(VCC_net), .CO(n59781));
    SB_CARRY encoder0_position_30__I_0_add_1101_12 (.CI(n59286), .I0(n1624), 
            .I1(VCC_net), .CO(n59287));
    SB_CARRY add_151_6 (.CI(n58880), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n58881));
    SB_LUT4 encoder0_position_30__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n59285), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n59779), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_11 (.CI(n59285), .I0(n1625), 
            .I1(VCC_net), .CO(n59286));
    SB_CARRY add_151_15 (.CI(n58889), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n58890));
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n58888), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n59284), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_13 (.CI(n59779), .I0(n3023), 
            .I1(VCC_net), .CO(n59780));
    SB_CARRY encoder0_position_30__I_0_add_1101_10 (.CI(n59284), .I0(n1626), 
            .I1(VCC_net), .CO(n59285));
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n58877));
    SB_LUT4 encoder0_position_30__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n59283), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n59778), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_9 (.CI(n59283), .I0(n1627), 
            .I1(VCC_net), .CO(n59284));
    SB_LUT4 encoder0_position_30__I_0_i837_3_lut (.I0(n1226_adj_5838), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n66693));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n59282), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_12 (.CI(n59778), .I0(n3024), 
            .I1(VCC_net), .CO(n59779));
    SB_CARRY encoder0_position_30__I_0_add_1101_8 (.CI(n59282), .I0(n1628), 
            .I1(VCC_net), .CO(n59283));
    SB_LUT4 encoder0_position_30__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n59777), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n59281), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_11 (.CI(n59777), .I0(n3025), 
            .I1(VCC_net), .CO(n59778));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n66692));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1101_7 (.CI(n59281), .I0(n1629), 
            .I1(GND_net), .CO(n59282));
    SB_LUT4 encoder0_position_30__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n59776), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n59280), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_10 (.CI(n59776), .I0(n3026), 
            .I1(VCC_net), .CO(n59777));
    SB_CARRY encoder0_position_30__I_0_add_1101_6 (.CI(n59280), .I0(n1630), 
            .I1(GND_net), .CO(n59281));
    SB_LUT4 encoder0_position_30__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n59775), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n59279), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_9 (.CI(n59775), .I0(n3027), 
            .I1(VCC_net), .CO(n59776));
    SB_CARRY encoder0_position_30__I_0_add_1101_5 (.CI(n59279), .I0(n1631), 
            .I1(VCC_net), .CO(n59280));
    SB_LUT4 encoder0_position_30__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n59774), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n59278), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_8 (.CI(n59774), .I0(n3028), 
            .I1(VCC_net), .CO(n59775));
    SB_CARRY encoder0_position_30__I_0_add_1101_4 (.CI(n59278), .I0(n1632), 
            .I1(GND_net), .CO(n59279));
    SB_LUT4 encoder0_position_30__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n59277), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3812_i23_3_lut (.I0(encoder0_position[22]), .I1(n10_adj_5740), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n935));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n59773), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_3 (.CI(n59277), .I0(n1633), 
            .I1(VCC_net), .CO(n59278));
    SB_CARRY encoder0_position_30__I_0_add_2039_7 (.CI(n59773), .I0(n3029), 
            .I1(GND_net), .CO(n59774));
    SB_LUT4 encoder0_position_30__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n59277));
    SB_LUT4 encoder0_position_30__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n59772), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_6 (.CI(n59772), .I0(n3030), 
            .I1(GND_net), .CO(n59773));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n66691));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n66690));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n66689));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n66688));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n66687));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i709_3_lut (.I0(n935), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232_adj_5844));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i843_3_lut (.I0(n1232_adj_5844), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n66686));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1178_3_lut (.I0(n1727), .I1(n1794_adj_5849), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n66685));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n66684));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n66683));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n66682));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n66681));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n66680));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n66679));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n66678));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n66677));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n66676));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 i15955_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n66866), 
            .I3(GND_net), .O(n30169));   // verilog/coms.v(130[12] 305[6])
    defparam i15955_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n66675));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 mux_3812_i27_3_lut (.I0(encoder0_position[26]), .I1(n6_adj_5745), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n66674));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 mux_3812_i28_3_lut (.I0(encoder0_position[27]), .I1(n5), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n291_adj_5806));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_2_lut (.I0(pwm_setpoint[19]), .I1(pwm_counter[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/pwm.v(11[19:30])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_2_lut_adj_1978 (.I0(pwm_setpoint[20]), .I1(pwm_counter[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(11[19:30])
    defparam i10_2_lut_adj_1978.LUT_INIT = 16'h6666;
    SB_LUT4 i11_2_lut_adj_1979 (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5859));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i11_2_lut_adj_1979.LUT_INIT = 16'h6666;
    SB_LUT4 mux_3812_i29_3_lut (.I0(encoder0_position[28]), .I1(n4_adj_5746), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n66673));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n66672));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 i9_2_lut_adj_1982 (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5858));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i9_2_lut_adj_1982.LUT_INIT = 16'h6666;
    SB_LUT4 i12_2_lut_adj_1983 (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5857));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i12_2_lut_adj_1983.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n66671));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1985 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n66670));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1985.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n66669));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n66668));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n66667));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i16824_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n31038));   // verilog/coms.v(130[12] 305[6])
    defparam i16824_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n66666));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n66665));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n66664));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_3_lut_adj_1992 (.I0(reset), .I1(n41637), .I2(n8_adj_5835), 
            .I3(GND_net), .O(n28713));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut_adj_1992.LUT_INIT = 16'h0404;
    SB_LUT4 i23431_3_lut (.I0(n32_adj_5860), .I1(pwm_counter[16]), .I2(pwm_setpoint[16]), 
            .I3(GND_net), .O(n34));   // verilog/pwm.v(11[19:30])
    defparam i23431_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 mux_3812_i30_3_lut (.I0(encoder0_position[29]), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6167_2_lut (.I0(n2_adj_5747), .I1(encoder0_position[30]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i6167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1993 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n66663));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1993.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n66662));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n66661));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1996 (.I0(n2413), .I1(n2417), .I2(n2420), .I3(n71130), 
            .O(n71136));
    defparam i1_4_lut_adj_1996.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n66660));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i62664_4_lut (.I0(n71136), .I1(n2412), .I2(n71212), .I3(n2414), 
            .O(n2445));
    defparam i62664_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1172_3_lut (.I0(n1721), .I1(n1788_adj_5846), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1998 (.I0(n2524), .I1(n2528), .I2(n2523), .I3(n2520), 
            .O(n71232));
    defparam i1_4_lut_adj_1998.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i10_3_lut (.I0(encoder0_position[9]), .I1(n23_adj_5726), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31351_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n45446));
    defparam i31351_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1999 (.I0(n2525), .I1(n2521), .I2(GND_net), .I3(GND_net), 
            .O(n70766));
    defparam i1_2_lut_adj_1999.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2000 (.I0(n2519), .I1(n71232), .I2(n2527), .I3(n2526), 
            .O(n71236));
    defparam i1_4_lut_adj_2000.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2001 (.I0(n2529), .I1(n45446), .I2(n2530), .I3(n2531), 
            .O(n68507));
    defparam i1_4_lut_adj_2001.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2002 (.I0(n68507), .I1(n71236), .I2(n70766), 
            .I3(n2517), .O(n70770));
    defparam i1_4_lut_adj_2002.LUT_INIT = 16'hfffe;
    SB_LUT4 i15958_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n66862), 
            .I3(GND_net), .O(n30172));   // verilog/coms.v(130[12] 305[6])
    defparam i15958_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n66659));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n66658));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2005 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n66657));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2005.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2006 (.I0(n2516), .I1(n2518), .I2(n2522), .I3(GND_net), 
            .O(n71058));
    defparam i1_3_lut_adj_2006.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n66656));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2008 (.I0(n71058), .I1(n2514), .I2(n70770), .I3(n2515), 
            .O(n70774));
    defparam i1_4_lut_adj_2008.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n66655));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n66654));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62787_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n70774), 
            .O(n2544));
    defparam i62787_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i51835_3_lut (.I0(n6_adj_5745), .I1(n7760), .I2(n67628), .I3(GND_net), 
            .O(n67635));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2011 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n66653));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2011.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2012 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n66652));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2012.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n66651));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2014 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n66650));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2014.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_3_lut_adj_2015 (.I0(reset), .I1(n41637), .I2(n8_adj_5748), 
            .I3(GND_net), .O(n28717));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut_adj_2015.LUT_INIT = 16'h0404;
    SB_LUT4 i1_4_lut_adj_2016 (.I0(n67238), .I1(n67584), .I2(Kp_23__N_1389), 
            .I3(\data_in_frame[13] [7]), .O(n71574));
    defparam i1_4_lut_adj_2016.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2017 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n66649));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2017.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2018 (.I0(n67194), .I1(n16_adj_5752), .I2(n71574), 
            .I3(n69065), .O(n71578));
    defparam i1_4_lut_adj_2018.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2019 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n66648));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2019.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2020 (.I0(n27203), .I1(n67135), .I2(n25590), 
            .I3(n71578), .O(n67500));
    defparam i1_4_lut_adj_2020.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_2021 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n71716));
    defparam i1_2_lut_adj_2021.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_2022 (.I0(n67235), .I1(\data_in_frame[17] [5]), 
            .I2(n71716), .I3(\data_in_frame[14] [6]), .O(n71722));
    defparam i1_4_lut_adj_2022.LUT_INIT = 16'h6996;
    SB_LUT4 i51836_3_lut (.I0(encoder0_position[26]), .I1(n67635), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2023 (.I0(n66945), .I1(n67596), .I2(n67578), 
            .I3(n71722), .O(n71728));
    defparam i1_4_lut_adj_2023.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2024 (.I0(n67213), .I1(n67500), .I2(n61396), 
            .I3(n71728), .O(n69485));
    defparam i1_4_lut_adj_2024.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2025 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n66647));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2025.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2026 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n66646));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2026.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2027 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n66645));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2027.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2028 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n66644));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2028.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_adj_2029 (.I0(n5_adj_5956), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n71200));
    defparam i1_3_lut_adj_2029.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_30__I_0_i500_4_lut (.I0(n2_adj_5747), .I1(n7756), 
            .I2(n71200), .I3(encoder0_position[30]), .O(n828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2030 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n66643));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2030.LUT_INIT = 16'h2300;
    SB_LUT4 i14_2_lut (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5749));   // verilog/coms.v(99[12:25])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2031 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n66642));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2031.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n66641));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_2033 (.I0(\data_in_frame[14] [5]), .I1(n26875), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5937));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_2033.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_2034 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [4]), 
            .I2(n27243), .I3(n6_adj_5937), .O(n61396));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut_adj_2034.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2035 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n66580));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2035.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2036 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n66581));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2036.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2037 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n66582));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2037.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2038 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n66583));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2038.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2039 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n66584));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2039.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2040 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n66585));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2040.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut_adj_2041 (.I0(\data_in_frame[14] [4]), .I1(n69463), 
            .I2(\data_in_frame[12] [3]), .I3(n67243), .O(n26760));
    defparam i3_4_lut_adj_2041.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n66586));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2043 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n66588));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2043.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2044 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n29288));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2044.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2045 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n66589));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2045.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2046 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n66590));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2046.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2047 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n66591));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2047.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2048 (.I0(n2622), .I1(n2624), .I2(n2626), .I3(n2628), 
            .O(n71088));
    defparam i1_4_lut_adj_2048.LUT_INIT = 16'hfffe;
    SB_LUT4 i31421_4_lut (.I0(n951), .I1(n2631), .I2(n2632), .I3(n2633), 
            .O(n45516));
    defparam i31421_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_2049 (.I0(n2625), .I1(n2627), .I2(n2623), .I3(GND_net), 
            .O(n71066));
    defparam i1_3_lut_adj_2049.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228_adj_5840));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2050 (.I0(n2629), .I1(n2630), .I2(GND_net), .I3(GND_net), 
            .O(n71386));
    defparam i1_2_lut_adj_2050.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2051 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n66592));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2051.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2052 (.I0(n2619), .I1(n71386), .I2(n71066), .I3(n45516), 
            .O(n71070));
    defparam i1_4_lut_adj_2052.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2053 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n66593));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2053.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i839_3_lut (.I0(n1228_adj_5840), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2054 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n66594));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2054.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2055 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n66595));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2055.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2056 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n66596));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2056.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2057 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n66578));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2057.LUT_INIT = 16'h2300;
    SB_LUT4 i15561_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(n359), 
            .I2(n28076), .I3(GND_net), .O(n29775));   // verilog/motorControl.v(42[14] 73[8])
    defparam i15561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2058 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n29278));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2058.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2059 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n66597));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2059.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2060 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n66598));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2060.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2061 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n66599));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2061.LUT_INIT = 16'h2300;
    SB_LUT4 i16572_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n23094), .I3(GND_net), .O(n30786));   // verilog/coms.v(130[12] 305[6])
    defparam i16572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2062 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n66600));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2062.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2063 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n66601));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2063.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2064 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n66602));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2064.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2065 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n29271));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2065.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2066 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n66603));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2066.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2067 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n66604));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2067.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2068 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n66605));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2068.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2069 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n66606));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2069.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2070 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n66607));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2070.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2071 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n66576));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2071.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2072 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n66608));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2072.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2073 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n29263));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2073.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2074 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n66609));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2074.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2075 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n29261));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2075.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2076 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n66610));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2076.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2077 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n66611));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2077.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2078 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n66612));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2078.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2079 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n66613));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2079.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2080 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n66614));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2080.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2081 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n66615));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2081.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2082 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n66616));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2082.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2083 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n29253));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2083.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2084 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n66617));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2084.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2085 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n29251));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2085.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2086 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n66618));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2086.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2087 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n66619));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2087.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2088 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n66620));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2088.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2089 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n66621));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2089.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2090 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n66743));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2090.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2091 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n66742));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2091.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2092 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n66741));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2092.LUT_INIT = 16'h2300;
    SB_LUT4 i30471_2_lut (.I0(n23188), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n44559));
    defparam i30471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1174_3_lut (.I0(n1723), .I1(n1790_adj_5847), 
            .I2(n1752), .I3(GND_net), .O(n1822_adj_5851));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1241_3_lut (.I0(n1822_adj_5851), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2093 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n66740));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2093.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2094 (.I0(n2615), .I1(n2616), .I2(n2617), .I3(n71070), 
            .O(n71076));
    defparam i1_4_lut_adj_2094.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2095 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n66739));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2095.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2096 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n66738));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2096.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2097 (.I0(n2618), .I1(n2620), .I2(n2621), .I3(n71088), 
            .O(n71094));
    defparam i1_4_lut_adj_2097.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2098 (.I0(n2612), .I1(n2613), .I2(n2614), .I3(n71076), 
            .O(n71082));
    defparam i1_4_lut_adj_2098.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62693_4_lut (.I0(n2611), .I1(n71082), .I2(n71094), .I3(n2610), 
            .O(n2643));
    defparam i62693_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2099 (.I0(n2724), .I1(n2718), .I2(n2723), .I3(n2728), 
            .O(n70922));
    defparam i1_4_lut_adj_2099.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2100 (.I0(n2726), .I1(n2722), .I2(n2720), .I3(n2725), 
            .O(n70924));
    defparam i1_4_lut_adj_2100.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n44574), .O(n65060));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb1f1;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2101 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n66737));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2101.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2102 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n66736));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2102.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2103 (.I0(n70922), .I1(n2717), .I2(n2727), .I3(GND_net), 
            .O(n70926));
    defparam i1_3_lut_adj_2103.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2104 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n66735));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2104.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2105 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n66734));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2105.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2106 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n66733));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2106.LUT_INIT = 16'h2300;
    SB_LUT4 i15658_3_lut (.I0(\data_in_frame[23] [7]), .I1(rx_data[7]), 
            .I2(n28703), .I3(GND_net), .O(n29872));   // verilog/coms.v(130[12] 305[6])
    defparam i15658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2107 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n66732));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2107.LUT_INIT = 16'h2300;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[23] [6]), .I1(n45398), .I2(n28703), 
            .I3(rx_data[6]), .O(n65962));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2108 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n66731));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2108.LUT_INIT = 16'h2300;
    SB_LUT4 i11_4_lut_adj_2109 (.I0(\data_in_frame[23] [5]), .I1(n45398), 
            .I2(n28703), .I3(rx_data[5]), .O(n65964));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut_adj_2109.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2110 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n66730));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2110.LUT_INIT = 16'h2300;
    SB_LUT4 i31419_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n45514));
    defparam i31419_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i25_3_lut (.I0(encoder0_position[24]), .I1(n8), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2111 (.I0(n2715), .I1(n70926), .I2(n2716), .I3(n70924), 
            .O(n70932));
    defparam i1_4_lut_adj_2111.LUT_INIT = 16'hfffe;
    SB_LUT4 i15649_3_lut (.I0(\data_in_frame[23] [4]), .I1(rx_data[4]), 
            .I2(n28703), .I3(GND_net), .O(n29863));   // verilog/coms.v(130[12] 305[6])
    defparam i15649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2112 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n66729));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2112.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2113 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n66728));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2113.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2114 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n66727));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2114.LUT_INIT = 16'h2300;
    SB_LUT4 i59852_2_lut (.I0(n79), .I1(n45283), .I2(GND_net), .I3(GND_net), 
            .O(n75251));   // verilog/coms.v(94[13:20])
    defparam i59852_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2115 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n66726));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2115.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2116 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n66725));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2116.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2117 (.I0(n2729), .I1(n70932), .I2(n45514), .I3(n2730), 
            .O(n70934));
    defparam i1_4_lut_adj_2117.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2118 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n66724));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2118.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2119 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n66723));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2119.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2120 (.I0(n2711), .I1(n2713), .I2(n70934), .I3(n2714), 
            .O(n70940));
    defparam i1_4_lut_adj_2120.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_2121 (.I0(n2712), .I1(n2721), .I2(n2719), .I3(GND_net), 
            .O(n70946));
    defparam i1_3_lut_adj_2121.LUT_INIT = 16'hfefe;
    SB_LUT4 i27521_4_lut (.I0(n75251), .I1(n75250), .I2(rx_data[3]), .I3(\data_in_frame[23] [3]), 
            .O(n41654));   // verilog/coms.v(94[13:20])
    defparam i27521_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i27522_3_lut (.I0(n41654), .I1(\data_in_frame[23] [3]), .I2(reset), 
            .I3(GND_net), .O(n30469));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_2122 (.I0(\data_in_frame[23] [2]), .I1(n45398), 
            .I2(n28703), .I3(rx_data[2]), .O(n65966));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut_adj_2122.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2123 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n29387));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2123.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2124 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n66722));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2124.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62610_4_lut (.I0(n2709), .I1(n70946), .I2(n70940), .I3(n2710), 
            .O(n2742));
    defparam i62610_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230_adj_5842));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2125 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n66721));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2125.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2126 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n66720));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2126.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2127 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n66719));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2127.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2128 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n66718));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2128.LUT_INIT = 16'h2300;
    SB_LUT4 i44548_3_lut_4_lut (.I0(n37307), .I1(Ki[3]), .I2(n4_adj_5738), 
            .I3(n20467), .O(n6));
    defparam i44548_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2129 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n66717));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2129.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2130 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n66716));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2130.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_4_lut (.I0(n37307), .I1(Ki[3]), .I2(n4_adj_5738), 
            .I3(n20467), .O(n20421));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 encoder0_position_30__I_0_i841_3_lut (.I0(n1230_adj_5842), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2131 (.I0(n2823), .I1(n2827), .I2(n2826), .I3(n2825), 
            .O(n71170));
    defparam i1_4_lut_adj_2131.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2132 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n66715));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2132.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n6_adj_5743));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_2133 (.I0(n2814), .I1(n2815), .I2(n2824), .I3(n2828), 
            .O(n71144));
    defparam i1_4_lut_adj_2133.LUT_INIT = 16'hfffe;
    SB_LUT4 i15631_3_lut (.I0(\data_in_frame[23] [1]), .I1(rx_data[1]), 
            .I2(n28703), .I3(GND_net), .O(n29845));   // verilog/coms.v(130[12] 305[6])
    defparam i15631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(n61795), .I3(\data_out_frame[18] [5]), .O(n62302));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_2134 (.I0(\data_out_frame[17] [7]), .I1(n27184), 
            .I2(n67259), .I3(n62277), .O(n8_adj_5950));   // verilog/coms.v(100[12:26])
    defparam i3_3_lut_4_lut_adj_2134.LUT_INIT = 16'h9669;
    SB_LUT4 encoder0_position_30__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i56248_2_lut (.I0(color_bit_N_502[2]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n72094));
    defparam i56248_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2135 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n66714));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2135.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2136 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n66713));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2136.LUT_INIT = 16'h2300;
    SB_LUT4 i31367_3_lut (.I0(n953), .I1(n2832), .I2(n2833), .I3(GND_net), 
            .O(n45462));
    defparam i31367_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2137 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n66712));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2137.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_2138 (.I0(\data_out_frame[17] [7]), .I1(n27184), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n67425));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_2138.LUT_INIT = 16'h9696;
    SB_LUT4 i59672_4_lut (.I0(n72094), .I1(n61457), .I2(n61432), .I3(color_bit_N_502[1]), 
            .O(n75301));   // verilog/neopixel.v(34[12] 113[6])
    defparam i59672_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i1_4_lut_adj_2139 (.I0(n2820), .I1(n2821_adj_5854), .I2(n2822), 
            .I3(n71170), .O(n71176));
    defparam i1_4_lut_adj_2139.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1176_3_lut (.I0(n1725), .I1(n1792_adj_5848), 
            .I2(n1752), .I3(GND_net), .O(n1824_adj_5852));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2140 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n66711));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2140.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2141 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n29374));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2141.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1178_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5927));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59679_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n75535));   // verilog/uart_rx.v(119[17:57])
    defparam i59679_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_2142 (.I0(n2829), .I1(n45462), .I2(n2830), .I3(n2831), 
            .O(n68558));
    defparam i1_4_lut_adj_2142.LUT_INIT = 16'ha080;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2143 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n66710));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2143.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2144 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n66622));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2144.LUT_INIT = 16'h2300;
    SB_LUT4 i26_4_lut (.I0(n25406), .I1(n75301), .I2(state[1]), .I3(n4), 
            .O(n65800));   // verilog/neopixel.v(34[12] 113[6])
    defparam i26_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 encoder0_position_30__I_0_i1243_3_lut (.I0(n1824_adj_5852), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2145 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n66623));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2145.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2146 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n29244));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2146.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2147 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n29243));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2147.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2148 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n66624));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2148.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16879_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n31093));   // verilog/coms.v(130[12] 305[6])
    defparam i16879_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2149 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n66625));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2149.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2150 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n66626));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2150.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2151 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n66627));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2151.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2152 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n66628));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2152.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2153 (.I0(n2818), .I1(n2819), .I2(n68558), .I3(n71176), 
            .O(n71182));
    defparam i1_4_lut_adj_2153.LUT_INIT = 16'hfffe;
    SB_LUT4 i15628_3_lut (.I0(\data_in_frame[23] [0]), .I1(rx_data[0]), 
            .I2(n28703), .I3(GND_net), .O(n29842));   // verilog/coms.v(130[12] 305[6])
    defparam i15628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2154 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n66629));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2154.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2155 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n71144), 
            .O(n71150));
    defparam i1_4_lut_adj_2155.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16267_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n336), 
            .I2(n28076), .I3(GND_net), .O(n30481));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_2156 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n66790));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_2156.LUT_INIT = 16'h2222;
    SB_LUT4 i15625_3_lut (.I0(\data_in_frame[22] [7]), .I1(rx_data[7]), 
            .I2(n66853), .I3(GND_net), .O(n29839));   // verilog/coms.v(130[12] 305[6])
    defparam i15625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15622_3_lut (.I0(\data_in_frame[22] [6]), .I1(rx_data[6]), 
            .I2(n66853), .I3(GND_net), .O(n29836));   // verilog/coms.v(130[12] 305[6])
    defparam i15622_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_2157 (.I0(hall1), .I1(hall2), .I2(n21154), 
            .I3(GND_net), .O(n4_adj_5962));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut_adj_2157.LUT_INIT = 16'hf2f2;
    SB_LUT4 i15619_3_lut (.I0(\data_in_frame[22] [5]), .I1(rx_data[5]), 
            .I2(n66853), .I3(GND_net), .O(n29833));   // verilog/coms.v(130[12] 305[6])
    defparam i15619_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2158 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n29236));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2158.LUT_INIT = 16'h2300;
    SB_LUT4 i15616_3_lut (.I0(\data_in_frame[22] [4]), .I1(rx_data[4]), 
            .I2(n66853), .I3(GND_net), .O(n29830));   // verilog/coms.v(130[12] 305[6])
    defparam i15616_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2159 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n29235));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2159.LUT_INIT = 16'h2300;
    SB_LUT4 i16275_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(n337), 
            .I2(n28076), .I3(GND_net), .O(n30489));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n37117), .I2(n28076), 
            .I3(GND_net), .O(n30490));
    defparam i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2160 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n66587));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2160.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2161 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n66630));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2161.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2162 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n29232));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2162.LUT_INIT = 16'h2300;
    SB_LUT4 i15613_3_lut (.I0(\data_in_frame[22] [3]), .I1(rx_data[3]), 
            .I2(n66853), .I3(GND_net), .O(n29827));   // verilog/coms.v(130[12] 305[6])
    defparam i15613_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2163 (.I0(n2809), .I1(n2816), .I2(n2817), .I3(n71182), 
            .O(n71188));
    defparam i1_4_lut_adj_2163.LUT_INIT = 16'hfffe;
    SB_LUT4 i16281_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(n339), 
            .I2(n28076), .I3(GND_net), .O(n30495));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16282_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n340), 
            .I2(n28076), .I3(GND_net), .O(n30496));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2164 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n66709));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2164.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n37307), .I2(n28076), 
            .I3(GND_net), .O(n30497));
    defparam i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2165 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n66708));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2165.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2166 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n66707));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2166.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2167 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n29369));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2167.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2168 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n29231));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2168.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16284_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n342), 
            .I2(n28076), .I3(GND_net), .O(n30498));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_2169 (.I0(n37307), .I1(Ki[2]), .I2(n58586), 
            .I3(n20468), .O(n20422));
    defparam i1_3_lut_4_lut_adj_2169.LUT_INIT = 16'h8778;
    SB_LUT4 i44540_3_lut_4_lut (.I0(n37307), .I1(Ki[2]), .I2(n58586), 
            .I3(n20468), .O(n4_adj_5738));
    defparam i44540_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_2_lut_3_lut_adj_2170 (.I0(n69502), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[22] [5]), .I3(GND_net), .O(n67203));
    defparam i1_2_lut_3_lut_adj_2170.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2171 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n66631));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2171.LUT_INIT = 16'h2300;
    SB_LUT4 i62727_4_lut (.I0(n2810), .I1(n71188), .I2(n71150), .I3(n2808), 
            .O(n2841));
    defparam i62727_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_2172 (.I0(n69502), .I1(\data_out_frame[20] [3]), 
            .I2(n67274), .I3(GND_net), .O(n24045));
    defparam i1_2_lut_3_lut_adj_2172.LUT_INIT = 16'h6969;
    SB_LUT4 encoder0_position_30__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2173 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n66632));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2173.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2174 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n66633));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2174.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2175 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n66634));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2175.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2176 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n66635));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2176.LUT_INIT = 16'h2300;
    SB_LUT4 i16285_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n343), 
            .I2(n28076), .I3(GND_net), .O(n30499));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2177 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n66636));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2177.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16286_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n344), 
            .I2(n28076), .I3(GND_net), .O(n30500));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2178 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n29224));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2178.LUT_INIT = 16'h2300;
    SB_LUT4 mux_3812_i11_3_lut (.I0(encoder0_position[10]), .I1(n22_adj_5727), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2179 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n66579));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2179.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16287_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n345), 
            .I2(n28076), .I3(GND_net), .O(n30501));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16288_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n346), 
            .I2(n28076), .I3(GND_net), .O(n30502));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i8_3_lut (.I0(encoder0_position[7]), .I1(n25_adj_5724), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2180 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n66637));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2180.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22621_3_lut (.I0(n322), .I1(IntegralLimit[12]), .I2(n258), 
            .I3(GND_net), .O(n347));
    defparam i22621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2181 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n66638));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2181.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_1181_i15_2_lut (.I0(r_Clock_Count_adj_6048[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5925));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2182 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n66639));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2182.LUT_INIT = 16'h2300;
    SB_LUT4 i22622_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(n347), 
            .I2(n28076), .I3(GND_net), .O(n30503));
    defparam i22622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2183 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n66640));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2183.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2184 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n66706));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2184.LUT_INIT = 16'h2300;
    SB_LUT4 i15610_3_lut (.I0(\data_in_frame[22] [2]), .I1(rx_data[2]), 
            .I2(n66853), .I3(GND_net), .O(n29824));   // verilog/coms.v(130[12] 305[6])
    defparam i15610_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2185 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n29367));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2185.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2186 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n29366));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2186.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1181_i9_2_lut (.I0(r_Clock_Count_adj_6048[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5921));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2187 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n66705));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2187.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1181_i13_2_lut (.I0(r_Clock_Count_adj_6048[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5923));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i11_2_lut (.I0(r_Clock_Count_adj_6048[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5922));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2188 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n66704));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2188.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2189 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n66702));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2189.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2190 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [0]), 
            .O(n66701));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2190.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1181_i4_4_lut (.I0(r_Clock_Count_adj_6048[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_6048[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5918));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61828_3_lut (.I0(n4_adj_5918), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5922), 
            .I3(GND_net), .O(n77684));   // verilog/uart_tx.v(117[17:57])
    defparam i61828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61829_3_lut (.I0(n77684), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5923), 
            .I3(GND_net), .O(n77685));   // verilog/uart_tx.v(117[17:57])
    defparam i61829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i9_3_lut (.I0(encoder0_position[8]), .I1(n24_adj_5725), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60670_4_lut (.I0(n13_adj_5923), .I1(n11_adj_5922), .I2(n9_adj_5921), 
            .I3(n75544), .O(n76526));
    defparam i60670_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1181_i8_3_lut (.I0(n6_adj_5919), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5921), .I3(GND_net), .O(n8_adj_5920));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_2191 (.I0(n2921), .I1(n2927), .I2(n2926), .I3(GND_net), 
            .O(n71000));
    defparam i1_3_lut_adj_2191.LUT_INIT = 16'hfefe;
    SB_LUT4 i15692_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n70340), 
            .I3(n27_adj_5855), .O(n29906));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15692_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61732_3_lut (.I0(n77685), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5925), 
            .I3(GND_net), .O(n14_adj_5924));   // verilog/uart_tx.v(117[17:57])
    defparam i61732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61359_4_lut (.I0(n14_adj_5924), .I1(n8_adj_5920), .I2(n15_adj_5925), 
            .I3(n76526), .O(n77215));   // verilog/uart_tx.v(117[17:57])
    defparam i61359_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61360_3_lut (.I0(n77215), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_6048[8]), 
            .I3(GND_net), .O(n5220));   // verilog/uart_tx.v(117[17:57])
    defparam i61360_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16291_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n348), 
            .I2(n28076), .I3(GND_net), .O(n30505));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15607_3_lut (.I0(\data_in_frame[22] [1]), .I1(rx_data[1]), 
            .I2(n66853), .I3(GND_net), .O(n29821));   // verilog/coms.v(130[12] 305[6])
    defparam i15607_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51923_2_lut (.I0(r_SM_Main_adj_6047[2]), .I1(r_SM_Main_adj_6047[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67730));
    defparam i51923_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2192 (.I0(n2923), .I1(n2919), .I2(n2924), .I3(n2928), 
            .O(n71002));
    defparam i1_4_lut_adj_2192.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15696_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n70356), 
            .I3(n27_adj_5855), .O(n29910));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15696_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2193 (.I0(n2917), .I1(n2922), .I2(n2918), .I3(n2920), 
            .O(n71004));
    defparam i1_4_lut_adj_2193.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_3812_i12_3_lut (.I0(encoder0_position[11]), .I1(n21_adj_5728), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31369_3_lut (.I0(n954), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n45464));
    defparam i31369_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i22668_3_lut (.I0(n247), .I1(n299_adj_5790), .I2(n284), .I3(GND_net), 
            .O(n36832));
    defparam i22668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22669_3_lut (.I0(n36832), .I1(IntegralLimit[10]), .I2(n258), 
            .I3(GND_net), .O(n349));
    defparam i22669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15700_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n70276), 
            .I3(n27_adj_5855), .O(n29914));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15700_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2194 (.I0(n2914), .I1(n71004), .I2(n71002), .I3(n71000), 
            .O(n71010));
    defparam i1_4_lut_adj_2194.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16293_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(n349), 
            .I2(n28076), .I3(GND_net), .O(n30507));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i7_3_lut (.I0(encoder0_position[6]), .I1(n26), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2195 (.I0(n2929), .I1(n45464), .I2(n2930), .I3(n2931), 
            .O(n68527));
    defparam i1_4_lut_adj_2195.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2196 (.I0(n2916), .I1(n2915), .I2(n2925), .I3(GND_net), 
            .O(n70754));
    defparam i1_3_lut_adj_2196.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2197 (.I0(n68527), .I1(n2910), .I2(n2912), .I3(n71010), 
            .O(n69567));
    defparam i1_4_lut_adj_2197.LUT_INIT = 16'hfffe;
    SB_LUT4 i15701_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n70324), 
            .I3(n27_adj_5855), .O(n29915));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15701_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6653_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6653_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i6651_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6651_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i15720_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n70308), 
            .I3(n27_adj_5855), .O(n29934));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15720_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5750), .I3(n15_adj_5816), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_91[9]), 
            .I2(n15_adj_5793), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16294_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n350), 
            .I2(n28076), .I3(GND_net), .O(n30508));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6655_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i6655_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i15722_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n70388), 
            .I3(n27_adj_5855), .O(n29936));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15722_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16295_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(n351), 
            .I2(n28076), .I3(GND_net), .O(n30509));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15723_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n70372), 
            .I3(n27_adj_5855), .O(n29937));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15723_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16296_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n352), 
            .I2(n28076), .I3(GND_net), .O(n30510));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63437 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [4]), .I2(\data_out_frame[23] [4]), 
            .I3(byte_transmit_counter[1]), .O(n79240));
    defparam byte_transmit_counter_0__bdd_4_lut_63437.LUT_INIT = 16'he4aa;
    SB_LUT4 i59688_3_lut_4_lut (.I0(r_Clock_Count_adj_6048[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_6048[2]), .O(n75544));   // verilog/uart_tx.v(117[17:57])
    defparam i59688_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i6657_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i6657_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 LessThan_1181_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_6048[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5919));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i15727_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n23025), .I3(GND_net), .O(n29941));   // verilog/coms.v(130[12] 305[6])
    defparam i15727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16297_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n353), 
            .I2(n28076), .I3(GND_net), .O(n30511));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15729_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n23094), .I3(GND_net), .O(n29943));   // verilog/coms.v(130[12] 305[6])
    defparam i15729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16298_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(n354), 
            .I2(n28076), .I3(GND_net), .O(n30512));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16299_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(n355), 
            .I2(n28076), .I3(GND_net), .O(n30513));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16300_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(n356), 
            .I2(n28076), .I3(GND_net), .O(n30514));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16820_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n31034));   // verilog/coms.v(130[12] 305[6])
    defparam i16820_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16301_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(n357), 
            .I2(n28076), .I3(GND_net), .O(n30515));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15733_3_lut (.I0(current[0]), .I1(data_adj_6031[0]), .I2(n28099), 
            .I3(GND_net), .O(n29947));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16302_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(n358), 
            .I2(n28076), .I3(GND_net), .O(n30516));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16303_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n23025), .I3(GND_net), .O(n30517));   // verilog/coms.v(130[12] 305[6])
    defparam i16303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2198 (.I0(\data_in_frame[17] [4]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[4]), .O(n65990));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2198.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2199 (.I0(\data_in_frame[17] [3]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[3]), .O(n65994));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2199.LUT_INIT = 16'h3a0a;
    SB_LUT4 n79240_bdd_4_lut (.I0(n79240), .I1(\data_out_frame[21] [4]), 
            .I2(\data_out_frame[20] [4]), .I3(byte_transmit_counter[1]), 
            .O(n79243));
    defparam n79240_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15961_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n66862), 
            .I3(GND_net), .O(n30175));   // verilog/coms.v(130[12] 305[6])
    defparam i15961_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62469_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n44574), .I3(GND_net), .O(n28130));
    defparam i62469_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 mux_3812_i14_3_lut (.I0(encoder0_position[13]), .I1(n19_adj_5730), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59632_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n75123));
    defparam i59632_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 encoder0_position_30__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30586_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n44574), .I3(GND_net), .O(n44675));
    defparam i30586_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 encoder0_position_30__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2200 (.I0(n8_adj_5834), .I1(n41637), .I2(GND_net), 
            .I3(GND_net), .O(n28662));
    defparam i1_2_lut_adj_2200.LUT_INIT = 16'hbbbb;
    SB_LUT4 mux_3812_i15_3_lut (.I0(encoder0_position[14]), .I1(n18_adj_5731), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_2201 (.I0(\data_in_frame[17] [2]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[2]), .O(n65998));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2201.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16244_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n28715), .I3(GND_net), .O(n30458));   // verilog/coms.v(130[12] 305[6])
    defparam i16244_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(0)_U0  quad_counter0 (.\a_new[1] (a_new[1]), .\b_new[1] (b_new[1]), 
            .debounce_cnt_N_3833(debounce_cnt_N_3833), .a_prev(a_prev), 
            .b_prev(b_prev), .position_31__N_3836(position_31__N_3836), 
            .GND_net(GND_net), .ENCODER0_B_N_keep(ENCODER0_B_N), .n1779(clk16MHz), 
            .ENCODER0_A_N_keep(ENCODER0_A_N), .n30012(n30012), .n1742(n1742), 
            .n30008(n30008), .n29986(n29986), .n1744(n1744), .\encoder0_position[30] (encoder0_position[30]), 
            .\encoder0_position[29] (encoder0_position[29]), .\encoder0_position[28] (encoder0_position[28]), 
            .\encoder0_position[27] (encoder0_position[27]), .\encoder0_position[26] (encoder0_position[26]), 
            .\encoder0_position[25] (encoder0_position[25]), .\encoder0_position[24] (encoder0_position[24]), 
            .\encoder0_position[23] (encoder0_position[23]), .\encoder0_position[22] (encoder0_position[22]), 
            .\encoder0_position[21] (encoder0_position[21]), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(305[27] 311[6])
    SB_LUT4 mux_3812_i16_3_lut (.I0(encoder0_position[15]), .I1(n17_adj_5732), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), .I2(n28715), 
            .I3(GND_net), .O(n65960));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15745_3_lut (.I0(b_prev_adj_5797), .I1(b_new_adj_6011[1]), 
            .I2(debounce_cnt_N_3833_adj_5798), .I3(GND_net), .O(n29959));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15745_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15746_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[1]), 
            .I2(n10_adj_5953), .I3(n25932), .O(n29960));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15746_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_2202 (.I0(\data_in_frame[16] [7]), .I1(n28664), 
            .I2(n28717), .I3(rx_data[7]), .O(n65866));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2202.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15747_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[2]), 
            .I2(n4_adj_5787), .I3(n25890), .O(n29961));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15747_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15751_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[3]), 
            .I2(n4_adj_5787), .I3(n25932), .O(n29965));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15751_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15752_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[4]), 
            .I2(n4_adj_5788), .I3(n25890), .O(n29966));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15752_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15753_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[5]), 
            .I2(n4_adj_5788), .I3(n25932), .O(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15753_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_adj_2203 (.I0(n37307), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_2203.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_2204 (.I0(\data_in_frame[16] [4]), .I1(n28664), 
            .I2(n28717), .I3(rx_data[4]), .O(n65842));
    defparam i12_4_lut_adj_2204.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_4_lut_adj_2205 (.I0(n2909), .I1(n2911), .I2(n2913), .I3(n70754), 
            .O(n70760));
    defparam i1_4_lut_adj_2205.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_3812_i17_3_lut (.I0(encoder0_position[16]), .I1(n16_adj_5733), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63501 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[21] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(byte_transmit_counter[0]), .O(n79234));
    defparam byte_transmit_counter_1__bdd_4_lut_63501.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_2206 (.I0(\data_in_frame[16] [3]), .I1(n28664), 
            .I2(n28717), .I3(rx_data[3]), .O(n65870));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2206.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15754_3_lut (.I0(t0[0]), .I1(timer[0]), .I2(n3165), .I3(GND_net), 
            .O(n29968));   // verilog/neopixel.v(34[12] 113[6])
    defparam i15754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62759_4_lut (.I0(n2908), .I1(n2907), .I2(n70760), .I3(n69567), 
            .O(n2940));
    defparam i62759_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i12_4_lut_adj_2207 (.I0(\data_in_frame[16] [2]), .I1(n28664), 
            .I2(n28717), .I3(rx_data[2]), .O(n65874));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2207.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15755_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[6]), 
            .I2(n44782), .I3(n25890), .O(n29969));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15755_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16218_3_lut (.I0(\data_in_frame[16] [1]), .I1(rx_data[1]), 
            .I2(n28717), .I3(GND_net), .O(n30432));   // verilog/coms.v(130[12] 305[6])
    defparam i16218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_2208 (.I0(n8_adj_5748), .I1(n41637), .I2(GND_net), 
            .I3(GND_net), .O(n28664));
    defparam i1_2_lut_adj_2208.LUT_INIT = 16'hbbbb;
    SB_LUT4 i12_4_lut_adj_2209 (.I0(\data_in_frame[16] [0]), .I1(n28664), 
            .I2(n28717), .I3(rx_data[0]), .O(n65878));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2209.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15756_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6024[7]), 
            .I2(n44782), .I3(n25932), .O(n29970));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15756_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7583_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n21154));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i7583_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8841_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i8841_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51825_3_lut (.I0(n4_adj_5962), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n67625));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i51825_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 encoder0_position_30__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i18_3_lut (.I0(encoder0_position[17]), .I1(n15_adj_5734), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n940));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15758_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n23094), .I3(GND_net), .O(n29972));   // verilog/coms.v(130[12] 305[6])
    defparam i15758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15759_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n23094), .I3(GND_net), .O(n29973));   // verilog/coms.v(130[12] 305[6])
    defparam i15759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15760_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n23094), .I3(GND_net), .O(n29974));   // verilog/coms.v(130[12] 305[6])
    defparam i15760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15761_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n23094), .I3(GND_net), .O(n29975));   // verilog/coms.v(130[12] 305[6])
    defparam i15761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n79234_bdd_4_lut (.I0(n79234), .I1(\data_out_frame[22] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(byte_transmit_counter[0]), 
            .O(n79237));
    defparam n79234_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15762_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n23094), .I3(GND_net), .O(n29976));   // verilog/coms.v(130[12] 305[6])
    defparam i15762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_2210 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n69981));
    defparam i3_4_lut_adj_2210.LUT_INIT = 16'h0004;
    SB_LUT4 encoder0_position_30__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21136_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n23094), .I3(GND_net), .O(n29979));
    defparam i21136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15769_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n23094), .I3(GND_net), .O(n29983));   // verilog/coms.v(130[12] 305[6])
    defparam i15769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15770_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n23094), .I3(GND_net), .O(n29984));   // verilog/coms.v(130[12] 305[6])
    defparam i15770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15772_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29986));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15773_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n23094), .I3(GND_net), .O(n29987));   // verilog/coms.v(130[12] 305[6])
    defparam i15773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15774_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n23094), .I3(GND_net), .O(n29988));   // verilog/coms.v(130[12] 305[6])
    defparam i15774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15775_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n23094), .I3(GND_net), .O(n29989));   // verilog/coms.v(130[12] 305[6])
    defparam i15775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i26_3_lut (.I0(encoder0_position[25]), .I1(n7_adj_5744), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2211 (.I0(n4_adj_5746), .I1(n5), .I2(n731), .I3(n6_adj_5745), 
            .O(n5_adj_5956));
    defparam i1_4_lut_adj_2211.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_2212 (.I0(n3), .I1(n2_adj_5747), .I2(n5_adj_5956), 
            .I3(GND_net), .O(n67628));
    defparam i1_3_lut_adj_2212.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_30__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15776_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n23025), .I3(GND_net), .O(n29990));   // verilog/coms.v(130[12] 305[6])
    defparam i15776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30336_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n23025), .I3(GND_net), .O(n29991));
    defparam i30336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51833_3_lut (.I0(n5), .I1(n7759), .I2(n67628), .I3(GND_net), 
            .O(n67633));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821_adj_5854));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1920_3_lut (.I0(n2821_adj_5854), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i19_3_lut (.I0(encoder0_position[18]), .I1(n14_adj_5735), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51834_3_lut (.I0(encoder0_position[27]), .I1(n67633), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16184_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n66869), .I3(GND_net), .O(n30398));   // verilog/coms.v(130[12] 305[6])
    defparam i16184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16181_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n66869), .I3(GND_net), .O(n30395));   // verilog/coms.v(130[12] 305[6])
    defparam i16181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16178_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n66869), .I3(GND_net), .O(n30392));   // verilog/coms.v(130[12] 305[6])
    defparam i16178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i20_3_lut (.I0(encoder0_position[19]), .I1(n13_adj_5736), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n938));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59792_2_lut (.I0(n79447), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n75275));
    defparam i59792_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227_adj_5839));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16174_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n66869), .I3(GND_net), .O(n30388));   // verilog/coms.v(130[12] 305[6])
    defparam i16174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i21_3_lut (.I0(encoder0_position[20]), .I1(n12_adj_5737), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n937));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1180_3_lut (.I0(n1729), .I1(n1796_adj_5850), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i838_3_lut (.I0(n1227_adj_5839), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1178_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5929));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16168_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n66869), .I3(GND_net), .O(n30382));   // verilog/coms.v(130[12] 305[6])
    defparam i16168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1178_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5926));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_1178_i8_3_lut (.I0(n6_adj_5927), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5929), .I3(GND_net), .O(n8_adj_5928));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62239_4_lut (.I0(n8_adj_5928), .I1(n4_adj_5926), .I2(n9_adj_5929), 
            .I3(n75535), .O(n78095));   // verilog/uart_rx.v(119[17:57])
    defparam i62239_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i56527_3_lut (.I0(n4910), .I1(duty[20]), .I2(n11851), .I3(GND_net), 
            .O(n72383));
    defparam i56527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62240_3_lut (.I0(n78095), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n78096));   // verilog/uart_rx.v(119[17:57])
    defparam i62240_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62009_3_lut (.I0(n78096), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n77865));   // verilog/uart_rx.v(119[17:57])
    defparam i62009_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61999_3_lut (.I0(n77865), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n5217));   // verilog/uart_rx.v(119[17:57])
    defparam i61999_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i56529_3_lut (.I0(n72383), .I1(n72378), .I2(n11849), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i56529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56524_3_lut (.I0(n4909), .I1(duty[21]), .I2(n11851), .I3(GND_net), 
            .O(n72380));
    defparam i56524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56526_3_lut (.I0(n72380), .I1(n72378), .I2(n11849), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i56526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56522_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n11851), 
            .I3(GND_net), .O(n72378));
    defparam i56522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56521_3_lut (.I0(n4908), .I1(duty[22]), .I2(n11851), .I3(GND_net), 
            .O(n72377));
    defparam i56521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56523_3_lut (.I0(n72377), .I1(n72378), .I2(n11849), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i56523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15964_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n66862), 
            .I3(GND_net), .O(n30178));   // verilog/coms.v(130[12] 305[6])
    defparam i15964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15967_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n66862), 
            .I3(GND_net), .O(n30181));   // verilog/coms.v(130[12] 305[6])
    defparam i15967_3_lut.LUT_INIT = 16'hacac;
    motorControl control (.GND_net(GND_net), .IntegralLimit({IntegralLimit}), 
            .\Kp[4] (Kp[4]), .n20421(n20421), .\Kp[5] (Kp[5]), .PWMLimit({PWMLimit}), 
            .n284(n284), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[7] (Kp[7]), 
            .\Kp[6] (Kp[6]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .n258(n258), .n356(n356), 
            .\Ki[1] (Ki[1]), .n357(n357), .\Ki[0] (Ki[0]), .n339(n339), 
            .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .n239(n239), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Kp[15] (Kp[15]), 
            .\Ki[6] (Ki[6]), .n346(n346), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .n358(n358), 
            .n20422(n20422), .n299(n299_adj_5790), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .n56(n56), 
            .setpoint({setpoint}), .\motor_state[9] (motor_state[9]), .n340(n340), 
            .VCC_net(VCC_net), .\motor_state[8] (motor_state[8]), .n359(n359), 
            .\motor_state[7] (motor_state[7]), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .n336(n336), .\motor_state[6] (motor_state[6]), .\motor_state[5] (motor_state[5]), 
            .n21(n21_adj_5868), .n460(n460), .n461(n461), .n467(n467), 
            .n475(n475), .n462(n462), .n247(n247), .n37(n37_adj_5869), 
            .n9(n9_adj_5862), .n16(n16_adj_5863), .n34689(n34689), .n20(n20_adj_5864), 
            .n291(n291), .n25(n25_adj_5866), .n35(n35), .n33(n33), .n37_adj_27(n37), 
            .n41(n41_adj_5867), .n22(n22_adj_5865), .n105(n105), .n35782(n35782), 
            .n24(n24_adj_5875), .n36147(n36147), .n36361(n36361), .\motor_state[4] (motor_state[4]), 
            .n25921(n25921), .n4(n4_adj_5861), .n342(n342), .n337(n337), 
            .n37307(n37307), .n37117(n37117), .n137(n137), .n347(n347_adj_5909), 
            .n6(n6), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .deadband({deadband}), 
            .n8(n8_adj_5870), .n25_adj_28(n25_adj_5872), .n343(n343), 
            .n10(n10_adj_5871), .n34(n34_adj_5873), .n38(n38_adj_5874), 
            .n40(n40), .n38_adj_29(n38), .n36(n36), .n75815(n75815), 
            .n24_adj_30(n24_adj_5916), .n30516(n30516), .n30515(n30515), 
            .n30514(n30514), .n30513(n30513), .n30512(n30512), .n30511(n30511), 
            .n30510(n30510), .n30509(n30509), .n30508(n30508), .n30507(n30507), 
            .n30505(n30505), .n30503(n30503), .n30502(n30502), .n30501(n30501), 
            .n30500(n30500), .n30499(n30499), .n30498(n30498), .n30497(n30497), 
            .n30496(n30496), .n30495(n30495), .n30490(n30490), .n30489(n30489), 
            .n30481(n30481), .n29775(n29775), .n347_adj_31(n347), .\control_mode[0] (control_mode[0]), 
            .n53108(n53108), .\control_mode[1] (control_mode[1]), .n28076(n28076), 
            .n344(n344), .n348(n348), .n17(n17_adj_5954), .n45282(n45282), 
            .\motor_state[2] (motor_state[2]), .\motor_state[1] (motor_state[1]), 
            .\motor_state[0] (motor_state[0]), .n349(n349), .\motor_state[23] (motor_state[23]), 
            .n38_adj_32(n38_adj_5913), .\motor_state[22] (motor_state[22]), 
            .n350(n350), .\motor_state[21] (motor_state[21]), .n345(n345), 
            .n12(n12_adj_5853), .\motor_state[19] (motor_state[19]), .\motor_state[18] (motor_state[18]), 
            .\motor_state[17] (motor_state[17]), .n486(n486), .n351(n351), 
            .n110(n110), .\motor_state[16] (motor_state[16]), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .\motor_state[13] (motor_state[13]), 
            .n10_adj_33(n10_adj_5911), .n42994(n42994), .\motor_state[10] (motor_state[10]), 
            .n352(n352), .n353(n353), .n354(n354), .n58586(n58586), 
            .n322(n322), .n20467(n20467), .n20468(n20468), .n355(n355), 
            .n313(n313)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 303[4])
    SB_LUT4 i7290_3_lut (.I0(n4907), .I1(current[15]), .I2(n11849), .I3(GND_net), 
            .O(n21158));
    defparam i7290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15970_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n66862), 
            .I3(GND_net), .O(n30184));   // verilog/coms.v(130[12] 305[6])
    defparam i15970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7291_3_lut (.I0(n21158), .I1(duty[23]), .I2(n11851), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i7291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15779_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n23025), .I3(GND_net), .O(n29993));   // verilog/coms.v(130[12] 305[6])
    defparam i15779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15973_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n66862), 
            .I3(GND_net), .O(n30187));   // verilog/coms.v(130[12] 305[6])
    defparam i15973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15976_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n66862), 
            .I3(GND_net), .O(n30190));   // verilog/coms.v(130[12] 305[6])
    defparam i15976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15780_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n23025), .I3(GND_net), .O(n29994));   // verilog/coms.v(130[12] 305[6])
    defparam i15780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15979_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n66862), 
            .I3(GND_net), .O(n30193));   // verilog/coms.v(130[12] 305[6])
    defparam i15979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16161_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n66869), .I3(GND_net), .O(n30375));   // verilog/coms.v(130[12] 305[6])
    defparam i16161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16158_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n66872), .I3(GND_net), .O(n30372));   // verilog/coms.v(130[12] 305[6])
    defparam i16158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15781_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n23025), .I3(GND_net), .O(n29995));   // verilog/coms.v(130[12] 305[6])
    defparam i15781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16154_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n66872), .I3(GND_net), .O(n30368));   // verilog/coms.v(130[12] 305[6])
    defparam i16154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15782_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n23025), .I3(GND_net), .O(n29996));   // verilog/coms.v(130[12] 305[6])
    defparam i15782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15783_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n23025), .I3(GND_net), .O(n29997));   // verilog/coms.v(130[12] 305[6])
    defparam i15783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15784_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n23025), .I3(GND_net), .O(n29998));   // verilog/coms.v(130[12] 305[6])
    defparam i15784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16151_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n66872), .I3(GND_net), .O(n30365));   // verilog/coms.v(130[12] 305[6])
    defparam i16151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30335_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n23025), .I3(GND_net), .O(n29999));
    defparam i30335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15786_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n23025), .I3(GND_net), .O(n30000));   // verilog/coms.v(130[12] 305[6])
    defparam i15786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15787_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n23025), .I3(GND_net), .O(n30001));   // verilog/coms.v(130[12] 305[6])
    defparam i15787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_2213 (.I0(data_ready), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5965));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i2_3_lut_4_lut_adj_2213.LUT_INIT = 16'h080c;
    SB_LUT4 i15788_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n23025), .I3(GND_net), .O(n30002));   // verilog/coms.v(130[12] 305[6])
    defparam i15788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16148_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n66872), .I3(GND_net), .O(n30362));   // verilog/coms.v(130[12] 305[6])
    defparam i16148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5771));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5783));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5781));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5775));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_2214 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n44574), .O(n24_adj_5959));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_adj_2214.LUT_INIT = 16'hffbf;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5774));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5773));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5779));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5778));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n28117), .O(n62510));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5777));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5761));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5762));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31399_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n45494));
    defparam i31399_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i16141_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n66872), .I3(GND_net), .O(n30355));   // verilog/coms.v(130[12] 305[6])
    defparam i16141_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5758));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5759));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31517_4_lut (.I0(n829), .I1(n828), .I2(n45494), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i31517_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i51837_3_lut (.I0(n7_adj_5744), .I1(n7761), .I2(n67628), .I3(GND_net), 
            .O(n67637));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i3_3_lut (.I0(encoder0_position[2]), .I1(n30), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51838_3_lut (.I0(encoder0_position[25]), .I1(n67637), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5766));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5764));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_3812_i4_3_lut (.I0(encoder0_position[3]), .I1(n29), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31405_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n45500));
    defparam i31405_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_2215 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n70950));
    defparam i1_2_lut_adj_2215.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5763));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2216 (.I0(n927), .I1(n70950), .I2(n928), .I3(n45500), 
            .O(n960));
    defparam i1_4_lut_adj_2216.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_30__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5768));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59941_4_lut (.I0(n11_adj_5763), .I1(n9_adj_5764), .I2(n7_adj_5766), 
            .I3(n5_adj_5768), .O(n75797));
    defparam i59941_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31337_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n45432));
    defparam i31337_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_3812_i5_3_lut (.I0(encoder0_position[4]), .I1(n28), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5765), .I1(current_limit[9]), 
            .I2(n19_adj_5758), .I3(GND_net), .O(n16_adj_5760));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16341_3_lut (.I0(t0[10]), .I1(timer[10]), .I2(n3165), .I3(GND_net), 
            .O(n30555));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5769));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i61477_3_lut (.I0(n4_adj_5769), .I1(current_limit[5]), .I2(n11_adj_5763), 
            .I3(GND_net), .O(n77333));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i61477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61478_3_lut (.I0(n77333), .I1(current_limit[6]), .I2(n13_adj_5762), 
            .I3(GND_net), .O(n77334));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i61478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2217 (.I0(n1029), .I1(n45432), .I2(n1030), .I3(n1031), 
            .O(n68436));
    defparam i1_4_lut_adj_2217.LUT_INIT = 16'ha080;
    SB_LUT4 i59871_4_lut (.I0(n17_adj_5759), .I1(n15_adj_5761), .I2(n13_adj_5762), 
            .I3(n75797), .O(n75727));
    defparam i59871_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61677_4_lut (.I0(n16_adj_5760), .I1(n6_adj_5767), .I2(n19_adj_5758), 
            .I3(n75719), .O(n77533));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i61677_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i63077_4_lut (.I0(n1026), .I1(n68436), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i63077_4_lut.LUT_INIT = 16'h0001;
    \quadrature_decoder(0)  quad_counter1 (.\a_new[1] (a_new_adj_6010[1]), 
            .\b_new[1] (b_new_adj_6011[1]), .debounce_cnt_N_3833(debounce_cnt_N_3833_adj_5798), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1779(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .b_prev(b_prev_adj_5797), .GND_net(GND_net), .n1786(n1786), 
            .n1788(n1788), .n1790(n1790), .n1792(n1792), .n1794(n1794), 
            .n1796(n1796), .\encoder1_position[25] (encoder1_position[25]), 
            .\encoder1_position[24] (encoder1_position[24]), .\encoder1_position[23] (encoder1_position[23]), 
            .\encoder1_position[22] (encoder1_position[22]), .\encoder1_position[21] (encoder1_position[21]), 
            .\encoder1_position[20] (encoder1_position[20]), .\encoder1_position[19] (encoder1_position[19]), 
            .\encoder1_position[18] (encoder1_position[18]), .\encoder1_position[17] (encoder1_position[17]), 
            .\encoder1_position[16] (encoder1_position[16]), .\encoder1_position[15] (encoder1_position[15]), 
            .\encoder1_position[14] (encoder1_position[14]), .\encoder1_position[13] (encoder1_position[13]), 
            .\encoder1_position[12] (encoder1_position[12]), .\encoder1_position[11] (encoder1_position[11]), 
            .\encoder1_position[10] (encoder1_position[10]), .\encoder1_position[9] (encoder1_position[9]), 
            .\encoder1_position[8] (encoder1_position[8]), .\encoder1_position[7] (encoder1_position[7]), 
            .\encoder1_position[6] (encoder1_position[6]), .\encoder1_position[5] (encoder1_position[5]), 
            .\encoder1_position[4] (encoder1_position[4]), .\encoder1_position[3] (encoder1_position[3]), 
            .\encoder1_position[2] (encoder1_position[2]), .n1822(n1822), 
            .n1824(n1824), .VCC_net(VCC_net), .n30013(n30013), .a_prev(a_prev_adj_5796), 
            .n29959(n29959), .n29958(n29958), .n1784(n1784), .position_31__N_3836(position_31__N_3836_adj_5799)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(313[27] 319[6])
    SB_LUT4 i60539_3_lut (.I0(n77334), .I1(current_limit[7]), .I2(n15_adj_5761), 
            .I3(GND_net), .O(n76395));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i60539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62178_4_lut (.I0(n76395), .I1(n77533), .I2(n19_adj_5758), 
            .I3(n75727), .O(n78034));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i62178_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62179_3_lut (.I0(n78034), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n22_adj_5757));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i62179_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_2218 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5966));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_2218.LUT_INIT = 16'h7bde;
    SB_LUT4 encoder0_position_30__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16135_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n66872), .I3(GND_net), .O(n30349));   // verilog/coms.v(130[12] 305[6])
    defparam i16135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11851_bdd_4_lut_63606 (.I0(n11851), .I1(current[15]), .I2(duty[22]), 
            .I3(n11849), .O(n79150));
    defparam n11851_bdd_4_lut_63606.LUT_INIT = 16'he4aa;
    SB_LUT4 n79150_bdd_4_lut (.I0(n79150), .I1(duty[19]), .I2(n4911), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[19]));
    defparam n79150_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229_adj_5841));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i840_3_lut (.I0(n1229_adj_5841), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_2219 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [2]), .I3(\data_out_frame[20] [1]), 
            .O(n26999));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_2219.LUT_INIT = 16'h6996;
    SB_LUT4 n11851_bdd_4_lut_63287 (.I0(n11851), .I1(current[15]), .I2(duty[21]), 
            .I3(n11849), .O(n79126));
    defparam n11851_bdd_4_lut_63287.LUT_INIT = 16'he4aa;
    SB_LUT4 n79126_bdd_4_lut (.I0(n79126), .I1(duty[18]), .I2(n4912), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[18]));
    defparam n79126_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5707));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i63250_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5970));
    defparam i63250_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 encoder0_position_30__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5753));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n11851_bdd_4_lut_63268 (.I0(n11851), .I1(current[15]), .I2(duty[20]), 
            .I3(n11849), .O(n79120));
    defparam n11851_bdd_4_lut_63268.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15798_3_lut_4_lut (.I0(n1742), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3836), .O(n30012));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15798_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5755));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59714_4_lut (.I0(n11), .I1(n9), .I2(n7_adj_5753), .I3(n5_adj_5755), 
            .O(n75570));
    defparam i59714_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1956_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n44574), .O(n6903));   // verilog/TinyFPGA_B.v(362[5] 388[12])
    defparam i1956_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i15793_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n30007));   // verilog/coms.v(130[12] 305[6])
    defparam i15793_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17), .I3(GND_net), 
            .O(n8_adj_5751));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n79120_bdd_4_lut (.I0(n79120), .I1(duty[17]), .I2(n4913), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[17]));
    defparam n79120_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7_adj_5753), 
            .I3(GND_net), .O(n6_adj_5754));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11851_bdd_4_lut_63263 (.I0(n11851), .I1(current[15]), .I2(duty[19]), 
            .I3(n11849), .O(n79114));
    defparam n11851_bdd_4_lut_63263.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5751), .I1(n301), .I2(n19_adj_5707), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_2220 (.I0(duty[17]), .I1(duty[22]), .I2(n294), 
            .I3(GND_net), .O(n8_adj_5936));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i2_3_lut_adj_2220.LUT_INIT = 16'h7e7e;
    SB_LUT4 i4_4_lut_adj_2221 (.I0(duty[21]), .I1(n8_adj_5936), .I2(duty[15]), 
            .I3(n294), .O(n10_adj_5935));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i4_4_lut_adj_2221.LUT_INIT = 16'hdffe;
    SB_LUT4 i5_4_lut_adj_2222 (.I0(duty[14]), .I1(n10_adj_5935), .I2(duty[18]), 
            .I3(n294), .O(n69858));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i5_4_lut_adj_2222.LUT_INIT = 16'hdffe;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n305), .I1(n304), .I2(n13), .I3(GND_net), 
            .O(n10));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n75098), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5756));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    coms neopxl_color_23__I_0 (.VCC_net(VCC_net), .clk16MHz(clk16MHz), .\Kp[6] (Kp[6]), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), 
         .encoder0_position_scaled({encoder0_position_scaled}), .byte_transmit_counter({Open_3, 
         Open_4, Open_5, Open_6, Open_7, byte_transmit_counter[2:0]}), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n2874(n2874), .\data_out_frame[8] ({\data_out_frame[8] }), .n66744(n66744), 
         .n66703(n66703), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .reset(reset), .rx_data({rx_data}), .\data_in_frame[11] ({\data_in_frame[11] [7], 
         Open_8, Open_9, Open_10, Open_11, Open_12, Open_13, Open_14}), 
         .\Kp[5] (Kp[5]), .GND_net(GND_net), .\Kp[4] (Kp[4]), .\data_out_frame[1][6] (\data_out_frame[1] [6]), 
         .\data_out_frame[3][6] (\data_out_frame[3] [6]), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .n67085(n67085), 
         .n79(n79), .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\Kp[3] (Kp[3]), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n25419(n25419), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n67203(n67203), .n26999(n26999), .\Kp[2] (Kp[2]), .displacement({displacement}), 
         .DE_c(DE_c), .\Kp[1] (Kp[1]), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .pwm_setpoint({pwm_setpoint}), .IntegralLimit({IntegralLimit}), 
         .n24045(n24045), .LED_c(LED_c), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .n30193(n30193), .\data_in_frame[6] ({\data_in_frame[6] }), .n30190(n30190), 
         .n30187(n30187), .n30184(n30184), .n30181(n30181), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n30178(n30178), .n26619(n26619), .\data_out_frame[1][3] (\data_out_frame[1] [3]), 
         .n69502(n69502), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .setpoint({setpoint}), .n62277(n62277), .n62302(n62302), .n30175(n30175), 
         .n29359(n29359), .\data_in_frame[12][6] (\data_in_frame[12] [6]), 
         .\data_in_frame[19] ({Open_15, Open_16, Open_17, Open_18, Open_19, 
         Open_20, Open_21, \data_in_frame[19] [0]}), .\data_in_frame[16] ({Open_22, 
         Open_23, Open_24, \data_in_frame[16] [4:1], Open_25}), .deadband({deadband}), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n66700(n66700), 
         .n30172(n30172), .n8(n8_adj_5950), .n67425(n67425), .\data_in_frame[16][7] (\data_in_frame[16] [7]), 
         .\data_out_frame[1][7] (\data_out_frame[1] [7]), .\data_out_frame[3][7] (\data_out_frame[3] [7]), 
         .n28392(n28392), .n30169(n30169), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n66699(n66699), .n72460(n72460), .n72458(n72458), .n66577(n66577), 
         .n66698(n66698), .\data_out_frame[9] ({\data_out_frame[9] }), .n66697(n66697), 
         .n66696(n66696), .n66695(n66695), .n66694(n66694), .n27(n27_adj_5910), 
         .n66693(n66693), .n66692(n66692), .n66691(n66691), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n66690(n66690), .n66689(n66689), .n66688(n66688), .n66687(n66687), 
         .n66686(n66686), .n66685(n66685), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n66684(n66684), .n66683(n66683), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .n66682(n66682), .n66681(n66681), .n66680(n66680), .n66679(n66679), 
         .n66678(n66678), .n66677(n66677), .n66676(n66676), .n66675(n66675), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .n66674(n66674), 
         .n66673(n66673), .n66672(n66672), .n66671(n66671), .n66670(n66670), 
         .n66669(n66669), .\data_in_frame[15][5] (\data_in_frame[15] [5]), 
         .n66668(n66668), .n30166(n30166), .n66667(n66667), .\FRAME_MATCHER.i[1] (\FRAME_MATCHER.i [1]), 
         .\data_in_frame[14] ({Open_26, Open_27, Open_28, Open_29, Open_30, 
         Open_31, Open_32, \data_in_frame[14] [0]}), .\FRAME_MATCHER.i[2] (\FRAME_MATCHER.i [2]), 
         .n66666(n66666), .n25421(n25421), .n30163(n30163), .n30160(n30160), 
         .n30157(n30157), .n30154(n30154), .\data_in_frame[14][2] (\data_in_frame[14] [2]), 
         .n30151(n30151), .n66665(n66665), .n67274(n67274), .n30148(n30148), 
         .\FRAME_MATCHER.i[0] (\FRAME_MATCHER.i [0]), .n62281(n62281), .\data_in_frame[14][4] (\data_in_frame[14] [4]), 
         .n69075(n69075), .\data_in_frame[14][5] (\data_in_frame[14] [5]), 
         .\data_in_frame[14][6] (\data_in_frame[14] [6]), .\data_in_frame[14][7] (\data_in_frame[14] [7]), 
         .\data_in_frame[13][2] (\data_in_frame[13] [2]), .n66664(n66664), 
         .\data_in_frame[13][4] (\data_in_frame[13] [4]), .n30145(n30145), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[13][5] (\data_in_frame[13] [5]), 
         .\data_in_frame[13][6] (\data_in_frame[13] [6]), .n30141(n30141), 
         .n30138(n30138), .n8_adj_5(n8_adj_5748), .n30135(n30135), .\data_in_frame[13][7] (\data_in_frame[13] [7]), 
         .n30132(n30132), .n23094(n23094), .n30129(n30129), .n67599(n67599), 
         .n30126(n30126), .n30123(n30123), .n67361(n67361), .\data_in_frame[12][2] (\data_in_frame[12] [2]), 
         .\data_in_frame[12][3] (\data_in_frame[12] [3]), .PWMLimit({PWMLimit}), 
         .n35(n35), .\data_in_frame[12][5] (\data_in_frame[12] [5]), .n462(n462), 
         .n36361(n36361), .\data_in_frame[12][4] (\data_in_frame[12] [4]), 
         .n105(n105), .control_mode({Open_33, Open_34, Open_35, Open_36, 
         control_mode[3:0]}), .control_update(control_update), .n24(n24_adj_5916), 
         .n30(n30_adj_5912), .n27184(n27184), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .\data_out_frame[3][4] (\data_out_frame[3] [4]), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n66663(n66663), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .\data_out_frame[3][3] (\data_out_frame[3] [3]), .n66662(n66662), 
         .n66661(n66661), .n66660(n66660), .n66659(n66659), .n66658(n66658), 
         .n66657(n66657), .n66656(n66656), .n66655(n66655), .n66654(n66654), 
         .n66653(n66653), .n66652(n66652), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .\data_out_frame[3][1] (\data_out_frame[3] [1]), .n66651(n66651), 
         .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .n66650(n66650), 
         .n66649(n66649), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), 
         .n66648(n66648), .n66647(n66647), .n66646(n66646), .\Kp[13] (Kp[13]), 
         .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), 
         .\Ki[3] (Ki[3]), .n66645(n66645), .n66644(n66644), .n66643(n66643), 
         .n66642(n66642), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .n66641(n66641), 
         .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .n66580(n66580), .n66581(n66581), 
         .n66582(n66582), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
         .n66583(n66583), .\Ki[11] (Ki[11]), .n66584(n66584), .n66585(n66585), 
         .n66586(n66586), .\Ki[12] (Ki[12]), .n66588(n66588), .n30873(n30873), 
         .n29288(n29288), .n66589(n66589), .n66590(n66590), .\Ki[13] (Ki[13]), 
         .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .n66591(n66591), .n66592(n66592), 
         .n66593(n66593), .n66594(n66594), .n66595(n66595), .n66596(n66596), 
         .n66578(n66578), .n30883(n30883), .n29278(n29278), .n30007(n30007), 
         .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n30003(n30003), .neopxl_color({neopxl_color}), .n30002(n30002), 
         .n30001(n30001), .n30000(n30000), .n29999(n29999), .n29998(n29998), 
         .n29997(n29997), .n29996(n29996), .n29995(n29995), .n29994(n29994), 
         .n29993(n29993), .n75275(n75275), .n29991(n29991), .n29990(n29990), 
         .n29989(n29989), .n29988(n29988), .n29987(n29987), .n29984(n29984), 
         .\control_mode[5] (control_mode[5]), .n29983(n29983), .\control_mode[6] (control_mode[6]), 
         .n29979(n29979), .\control_mode[7] (control_mode[7]), .n29976(n29976), 
         .\current_limit[1] (current_limit[1]), .n29975(n29975), .\current_limit[2] (current_limit[2]), 
         .n29974(n29974), .\current_limit[3] (current_limit[3]), .n29973(n29973), 
         .\current_limit[4] (current_limit[4]), .n29972(n29972), .\current_limit[5] (current_limit[5]), 
         .n29943(n29943), .\current_limit[0] (current_limit[0]), .n29941(n29941), 
         .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .n66597(n66597), .n66598(n66598), 
         .n66599(n66599), .n66600(n66600), .n66601(n66601), .n66602(n66602), 
         .n29271(n29271), .n66603(n66603), .n66604(n66604), .n66605(n66605), 
         .n66606(n66606), .n66607(n66607), .n66576(n66576), .n66608(n66608), 
         .n29263(n29263), .n66609(n66609), .n29261(n29261), .n66610(n66610), 
         .n66611(n66611), .n66612(n66612), .n66613(n66613), .n66614(n66614), 
         .n66615(n66615), .n66616(n66616), .n29253(n29253), .n66617(n66617), 
         .n29251(n29251), .n66618(n66618), .n66619(n66619), .n66620(n66620), 
         .n66621(n66621), .n66743(n66743), .n66742(n66742), .n66741(n66741), 
         .n38(n38_adj_5874), .n460(n460), .n486(n486), .n40(n40), .n41637(n41637), 
         .n66852(n66852), .n34(n34_adj_5873), .n36(n36), .n66740(n66740), 
         .n66739(n66739), .n30786(n30786), .\current_limit[8] (current_limit[8]), 
         .n45283(n45283), .encoder1_position_scaled({encoder1_position_scaled}), 
         .n53108(n53108), .n42994(n42994), .n30785(n30785), .\current_limit[9] (current_limit[9]), 
         .n30781(n30781), .\current_limit[10] (current_limit[10]), .n30779(n30779), 
         .\current_limit[12] (current_limit[12]), .n65900(n65900), .\data_in_frame[18] ({\data_in_frame[18] }), 
         .n65896(n65896), .n65892(n65892), .n65888(n65888), .\motor_state_23__N_91[12] (motor_state_23__N_91[12]), 
         .n15(n15_adj_5793), .n10(n10_adj_5911), .n29731(n29731), .n29734(n29734), 
         .n30740(n30740), .n65884(n65884), .n29740(n29740), .n30734(n30734), 
         .n29746(n29746), .\data_in_frame[19][2] (\data_in_frame[19] [2]), 
         .n30727(n30727), .\data_in_frame[17] ({\data_in_frame[17] }), .n29749(n29749), 
         .\data_in_frame[19][3] (\data_in_frame[19] [3]), .n29752(n29752), 
         .\data_in_frame[19][4] (\data_in_frame[19] [4]), .n29756(n29756), 
         .\data_in_frame[19][5] (\data_in_frame[19] [5]), .n30678(n30678), 
         .n30666(n30666), .\data_in_frame[9] ({\data_in_frame[9] }), .n66738(n66738), 
         .n30632(n30632), .n30249(n30249), .n29759(n29759), .\data_in_frame[19][6] (\data_in_frame[19] [6]), 
         .n30252(n30252), .n30255(n30255), .n29763(n29763), .\data_in_frame[19][7] (\data_in_frame[19] [7]), 
         .n30258(n30258), .n30261(n30261), .n30264(n30264), .n30619(n30619), 
         .n30616(n30616), .n66737(n66737), .\data_in_frame[20][0] (\data_in_frame[20] [0]), 
         .\data_in_frame[20][1] (\data_in_frame[20] [1]), .\data_in_frame[20][2] (\data_in_frame[20] [2]), 
         .\data_in_frame[20][4] (\data_in_frame[20] [4]), .n29794(n29794), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .n29797(n29797), .n30267(n30267), 
         .n30603(n30603), .n29800(n29800), .n29803(n29803), .n30593(n30593), 
         .n29806(n29806), .n30589(n30589), .n30588(n30588), .n29809(n29809), 
         .n30585(n30585), .n29812(n29812), .n29815(n29815), .n29818(n29818), 
         .\data_in_frame[22] ({\data_in_frame[22] }), .n66142(n66142), .n30349(n30349), 
         .\data_in_frame[13][0] (\data_in_frame[13] [0]), .n30355(n30355), 
         .n30362(n30362), .n30365(n30365), .n30368(n30368), .n30372(n30372), 
         .n30375(n30375), .n66736(n66736), .n66735(n66735), .n30382(n30382), 
         .n30388(n30388), .n30392(n30392), .n30395(n30395), .n30398(n30398), 
         .n65878(n65878), .\data_in_frame[16][0] (\data_in_frame[16] [0]), 
         .n30432(n30432), .n65874(n65874), .n65870(n65870), .n65842(n65842), 
         .n65866(n65866), .n65960(n65960), .n30458(n30458), .n65998(n65998), 
         .n65994(n65994), .n65990(n65990), .n30517(n30517), .n66734(n66734), 
         .n29821(n29821), .n29824(n29824), .n29827(n29827), .n29830(n29830), 
         .n29833(n29833), .n29836(n29836), .n29839(n29839), .n29842(n29842), 
         .\data_in_frame[23] ({\data_in_frame[23] }), .n29845(n29845), .n65966(n65966), 
         .n30469(n30469), .n29863(n29863), .n65964(n65964), .n65962(n65962), 
         .n29872(n29872), .n26875(n26875), .\data_in_frame[1][1] (\data_in_frame[1] [1]), 
         .\data_in_frame[1][2] (\data_in_frame[1] [2]), .\data_in_frame[1][3] (\data_in_frame[1] [3]), 
         .\data_in_frame[1][5] (\data_in_frame[1] [5]), .\data_in_frame[1][6] (\data_in_frame[1] [6]), 
         .\data_in_frame[1][7] (\data_in_frame[1] [7]), .n66733(n66733), 
         .n66732(n66732), .n66731(n66731), .n66730(n66730), .n66729(n66729), 
         .n66728(n66728), .n66727(n66727), .n66726(n66726), .n26311(n26311), 
         .n66725(n66725), .n66724(n66724), .n66723(n66723), .n26475(n26475), 
         .n29387(n29387), .n66722(n66722), .n66721(n66721), .n66720(n66720), 
         .n66719(n66719), .n66718(n66718), .n66717(n66717), .n66716(n66716), 
         .n66715(n66715), .n66714(n66714), .n66713(n66713), .n66712(n66712), 
         .n66711(n66711), .n29374(n29374), .n66710(n66710), .n66622(n66622), 
         .n66623(n66623), .n29755(n29755), .\current_limit[6] (current_limit[6]), 
         .n31022(n31022), .n29244(n29244), .n31023(n31023), .n29243(n29243), 
         .n66624(n66624), .n66625(n66625), .n66626(n66626), .n66627(n66627), 
         .n66628(n66628), .n66629(n66629), .n29236(n29236), .n31031(n31031), 
         .n29235(n29235), .n66587(n66587), .n66630(n66630), .n31034(n31034), 
         .n29232(n29232), .n66709(n66709), .n82(n82), .n28703(n28703), 
         .n28672(n28672), .n66708(n66708), .n66707(n66707), .n31038(n31038), 
         .n29369(n29369), .n31039(n31039), .n29231(n29231), .n66631(n66631), 
         .n66632(n66632), .n66633(n66633), .n66634(n66634), .n66635(n66635), 
         .n66636(n66636), .n31046(n31046), .n29224(n29224), .n66579(n66579), 
         .n66637(n66637), .n66638(n66638), .n66639(n66639), .n66640(n66640), 
         .n61795(n61795), .n66706(n66706), .n31088(n31088), .n29367(n29367), 
         .n29727(n29727), .\current_limit[7] (current_limit[7]), .n31093(n31093), 
         .n29366(n29366), .n66705(n66705), .n66704(n66704), .n66702(n66702), 
         .n66701(n66701), .n15_adj_6(n15_adj_5816), .rx_data_ready(rx_data_ready), 
         .n15_adj_7(n15_adj_5750), .\motor_state_23__N_91[8] (motor_state_23__N_91[8]), 
         .n25590(n25590), .n66867(n66867), .n66869(n66869), .n66862(n66862), 
         .\current[7] (current[7]), .\current[6] (current[6]), .\current[5] (current[5]), 
         .n67584(n67584), .\current[4] (current[4]), .n461(n461), .n38_adj_8(n38), 
         .n75815(n75815), .n6(n6_adj_5934), .n3476(n3476), .n66945(n66945), 
         .ID({ID}), .n79417(n79417), .n79243(n79243), .n1(n1), .n5(n5_adj_5951), 
         .n67259(n67259), .n27089(n27089), .n69485(n69485), .n67194(n67194), 
         .n6_adj_9(n6_adj_5749), .n69065(n69065), .n16(n16_adj_5752), 
         .n67500(n67500), .n67135(n67135), .n69463(n69463), .n27243(n27243), 
         .n26760(n26760), .n61396(n61396), .n67238(n67238), .n67596(n67596), 
         .n67235(n67235), .n89(n89), .n4(n4_adj_5861), .Kp_23__N_1389(Kp_23__N_1389), 
         .n25921(n25921), .\current[3] (current[3]), .\current[2] (current[2]), 
         .\current[1] (current[1]), .\current[0] (current[0]), .\current[15] (current[15]), 
         .n8_adj_10(n8_adj_5834), .n67578(n67578), .n8_adj_11(n8_adj_5835), 
         .n67243(n67243), .n61406(n61406), .n67213(n67213), .n28715(n28715), 
         .n75246(n75246), .n27203(n27203), .n66853(n66853), .\current[11] (current[11]), 
         .\current[10] (current[10]), .\current[9] (current[9]), .\current[8] (current[8]), 
         .n28730(n28730), .n75250(n75250), .n28717(n28717), .n10_adj_12(n10_adj_5960), 
         .n66872(n66872), .n66866(n66866), .n79237(n79237), .tx_active(tx_active), 
         .n23025(n23025), .n79447(n79447), .n51(n51), .n22(n22_adj_5757), 
         .n260(n260), .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_6047}), .n29956(n29956), 
         .r_Clock_Count({r_Clock_Count_adj_6048}), .n5220(n5220), .n27_adj_13(n27_adj_5855), 
         .n67730(n67730), .n6_adj_14(n6_adj_5955), .tx_enable(tx_enable), 
         .r_Clock_Count_adj_26({r_Clock_Count}), .baudrate({baudrate}), 
         .n28240(n28240), .n67800(n67800), .\r_SM_Main[2]_adj_23 (r_SM_Main[2]), 
         .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), 
         .n5217(n5217), .n66790(n66790), .\r_SM_Main[1]_adj_24 (r_SM_Main[1]), 
         .n28117(n28117), .n70292(n70292), .n29937(n29937), .n29936(n29936), 
         .n29934(n29934), .n29915(n29915), .n29914(n29914), .n29910(n29910), 
         .n29906(n29906), .n30762(n30762), .n62510(n62510), .n30758(n30758), 
         .\r_Bit_Index[0] (r_Bit_Index[0]), .n70662(n70662), .n34_adj_25(n34_adj_5961), 
         .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), 
         .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), 
         .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), 
         .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), 
         .n70340(n70340), .n70356(n70356), .n70276(n70276), .n70324(n70324), 
         .n70308(n70308), .n70388(n70388), .n70372(n70372)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i1_4_lut_4_lut_adj_2223 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2821), .O(n25_adj_5958));   // verilog/TinyFPGA_B.v(377[7:11])
    defparam i1_4_lut_4_lut_adj_2223.LUT_INIT = 16'h5450;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n10), .I1(n303), .I2(n15), .I3(GND_net), 
            .O(n12));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n79114_bdd_4_lut (.I0(n79114), .I1(duty[16]), .I2(n4914), 
            .I3(n11849), .O(pwm_setpoint_23__N_3[16]));
    defparam n79114_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i59708_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n75570), 
            .O(n75564));
    defparam i59708_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(reset), .I1(rx_data[3]), .I2(\data_in_frame[12] [3]), 
            .I3(n28672), .O(n66142));   // verilog/coms.v(94[13:20])
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hf0e4;
    SB_LUT4 i62166_4_lut (.I0(n16), .I1(n6_adj_5754), .I2(n19_adj_5707), 
            .I3(n75562), .O(n78022));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i62166_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61675_4_lut (.I0(n12), .I1(n4_adj_5756), .I2(n15), .I3(n75568), 
            .O(n77531));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61675_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62295_4_lut (.I0(n77531), .I1(n78022), .I2(n19_adj_5707), 
            .I3(n75564), .O(n78151));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i62295_4_lut.LUT_INIT = 16'hccca;
    TLI4970 tli (.GND_net(GND_net), .VCC_net(VCC_net), .n5(n5_adj_5791), 
            .n5_adj_3(n5_adj_5817), .n5_adj_4(n5_adj_5807), .state_7__N_4319(state_7__N_4319), 
            .n44711(n44711), .clk16MHz(clk16MHz), .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), 
            .n30119(n30119), .\data[15] (data_adj_6031[15]), .n30118(n30118), 
            .\data[12] (data_adj_6031[12]), .n30117(n30117), .\data[11] (data_adj_6031[11]), 
            .n30116(n30116), .\data[10] (data_adj_6031[10]), .n30115(n30115), 
            .\data[9] (data_adj_6031[9]), .n30114(n30114), .\data[8] (data_adj_6031[8]), 
            .n30113(n30113), .\data[7] (data_adj_6031[7]), .n30112(n30112), 
            .\data[6] (data_adj_6031[6]), .n30111(n30111), .\data[5] (data_adj_6031[5]), 
            .n30110(n30110), .\data[4] (data_adj_6031[4]), .n30109(n30109), 
            .\data[3] (data_adj_6031[3]), .n30108(n30108), .\data[2] (data_adj_6031[2]), 
            .n30107(n30107), .\data[1] (data_adj_6031[1]), .n29947(n29947), 
            .\current[0] (current[0]), .n30767(n30767), .\data[0] (data_adj_6031[0]), 
            .n30677(n30677), .\current[1] (current[1]), .n30676(n30676), 
            .\current[2] (current[2]), .n30675(n30675), .\current[3] (current[3]), 
            .n30674(n30674), .\current[4] (current[4]), .n30673(n30673), 
            .\current[5] (current[5]), .n30672(n30672), .\current[6] (current[6]), 
            .n30671(n30671), .\current[7] (current[7]), .n30670(n30670), 
            .\current[8] (current[8]), .n30669(n30669), .\current[9] (current[9]), 
            .n30668(n30668), .\current[10] (current[10]), .n30667(n30667), 
            .\current[11] (current[11]), .n28099(n28099), .\current[15] (current[15]), 
            .n25895(n25895), .n11(n11_adj_5792), .n25912(n25912), .n25869(n25869), 
            .n25885(n25885)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(405[11] 411[4])
    SB_LUT4 i62296_3_lut (.I0(n78151), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n78152));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i62296_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62246_3_lut (.I0(n78152), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n78102));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i62246_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_2224 (.I0(duty[16]), .I1(duty[13]), .I2(n294), 
            .I3(n69858), .O(n8_adj_5967));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i3_4_lut_adj_2224.LUT_INIT = 16'hff7e;
    SB_LUT4 i2_3_lut_adj_2225 (.I0(duty[20]), .I1(duty[19]), .I2(n294), 
            .I3(GND_net), .O(n7_adj_5968));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i2_3_lut_adj_2225.LUT_INIT = 16'h7e7e;
    SB_LUT4 i61719_3_lut (.I0(n78102), .I1(n298), .I2(duty[12]), .I3(GND_net), 
            .O(n77575));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61719_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61720_4_lut (.I0(n77575), .I1(n294), .I2(n7_adj_5968), .I3(n8_adj_5967), 
            .O(n77576));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61720_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_adj_2226 (.I0(n37117), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n137));
    defparam i1_2_lut_adj_2226.LUT_INIT = 16'h8888;
    SB_LUT4 i52039_4_lut (.I0(n260), .I1(duty[23]), .I2(n294), .I3(n77576), 
            .O(n11849));
    defparam i52039_4_lut.LUT_INIT = 16'h1151;
    SB_LUT4 i60664_3_lut (.I0(n15_adj_5777), .I1(n13_adj_5778), .I2(n11_adj_5779), 
            .I3(GND_net), .O(n76520));
    defparam i60664_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5784));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60468_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n76520), .O(n76324));
    defparam i60468_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i59581_4_lut (.I0(n21_adj_5773), .I1(n19_adj_5774), .I2(n17_adj_5775), 
            .I3(n9_adj_5781), .O(n75437));
    defparam i59581_4_lut.LUT_INIT = 16'haaab;
    pwm PWM (.n2874(n2874), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .\pwm_counter[7] (pwm_counter[7]), 
        .GND_net(GND_net), .\pwm_counter[16] (pwm_counter[16]), .\pwm_counter[20] (pwm_counter[20]), 
        .\pwm_counter[19] (pwm_counter[19]), .\pwm_counter[12] (pwm_counter[12]), 
        .\pwm_setpoint[18] (pwm_setpoint[18]), .\pwm_setpoint[17] (pwm_setpoint[17]), 
        .\pwm_counter[4] (pwm_counter[4]), .VCC_net(VCC_net), .reset(reset), 
        .\pwm_setpoint[22] (pwm_setpoint[22]), .\pwm_setpoint[21] (pwm_setpoint[21]), 
        .\pwm_setpoint[11] (pwm_setpoint[11]), .\pwm_setpoint[10] (pwm_setpoint[10]), 
        .\pwm_setpoint[9] (pwm_setpoint[9]), .\pwm_setpoint[6] (pwm_setpoint[6]), 
        .\pwm_setpoint[8] (pwm_setpoint[8]), .\pwm_setpoint[3] (pwm_setpoint[3]), 
        .\pwm_setpoint[5] (pwm_setpoint[5]), .\pwm_setpoint[2] (pwm_setpoint[2]), 
        .n9(n9_adj_5857), .n15(n15_adj_5858), .\pwm_setpoint[1] (pwm_setpoint[1]), 
        .\pwm_setpoint[0] (pwm_setpoint[0]), .\pwm_setpoint[7] (pwm_setpoint[7]), 
        .\pwm_setpoint[12] (pwm_setpoint[12]), .n25(n25_adj_5859), .\pwm_setpoint[13] (pwm_setpoint[13]), 
        .\pwm_setpoint[14] (pwm_setpoint[14]), .\pwm_setpoint[15] (pwm_setpoint[15]), 
        .n32(n32_adj_5860), .n34(n34), .\pwm_setpoint[20] (pwm_setpoint[20]), 
        .n41(n41), .n39(n39), .\pwm_setpoint[19] (pwm_setpoint[19]), .\pwm_setpoint[23] (pwm_setpoint[23]), 
        .\pwm_setpoint[4] (pwm_setpoint[4])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    SB_LUT4 encoder0_position_30__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22956_3_lut (.I0(n313), .I1(IntegralLimit[21]), .I2(n258), 
            .I3(GND_net), .O(n37117));
    defparam i22956_3_lut.LUT_INIT = 16'hcaca;
    EEPROM eeprom (.GND_net(GND_net), .enable_slow_N_4213(enable_slow_N_4213), 
           .clk16MHz(clk16MHz), .data({data_adj_6024}), .baudrate({baudrate}), 
           .n28272(n28272), .\state_7__N_3918[0] (state_7__N_3918[0]), .data_ready(data_ready), 
           .ID({ID}), .n30714(n30714), .n30713(n30713), .n30712(n30712), 
           .n30711(n30711), .n30710(n30710), .n30709(n30709), .n30708(n30708), 
           .n30707(n30707), .n30697(n30697), .n30696(n30696), .n30695(n30695), 
           .n30694(n30694), .n30693(n30693), .n30692(n30692), .n30691(n30691), 
           .n30690(n30690), .\state[0] (state_adj_6057[0]), .n28274(n28274), 
           .\state_7__N_4110[0] (state_7__N_4110[0]), .scl_enable(scl_enable), 
           .sda_enable(sda_enable), .sda_out(sda_out), .n29970(n29970), 
           .n29969(n29969), .n29967(n29967), .n29966(n29966), .n29965(n29965), 
           .n29961(n29961), .n29960(n29960), .n6707(n6707), .n30751(n30751), 
           .n8(n8_adj_5969), .VCC_net(VCC_net), .n11(n11_adj_5789), .\state_7__N_4126[3] (state_7__N_4126[3]), 
           .n44639(n44639), .n10(n10_adj_5953), .n4(n4_adj_5787), .n4_adj_2(n4_adj_5788), 
           .n25890(n25890), .n25932(n25932), .n44782(n44782), .scl(scl)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(391[10] 403[6])
    SB_LUT4 i15604_3_lut (.I0(\data_in_frame[22] [0]), .I1(rx_data[0]), 
            .I2(n66853), .I3(GND_net), .O(n29818));   // verilog/coms.v(130[12] 305[6])
    defparam i15604_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i60825_4_lut (.I0(n9_adj_5781), .I1(n7_adj_5783), .I2(current[2]), 
            .I3(duty[2]), .O(n76681));
    defparam i60825_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5780));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, bit_ctr, \color_bit_N_502[1] , 
            GND_net, neopxl_color, timer, state, n29968, t0, n28194, 
            \bit_ctr[3] , \bit_ctr[4] , VCC_net, n30584, n30583, n30582, 
            n30581, n30580, n30579, n30578, n30577, n30576, n30555, 
            n30479, n65800, NEOPXL_c, n61457, n61432, \color_bit_N_502[2] , 
            n44741, n25406, LED_c, n3165) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output [4:0]bit_ctr;
    output \color_bit_N_502[1] ;
    input GND_net;
    input [23:0]neopxl_color;
    output [10:0]timer;
    output [1:0]state;
    input n29968;
    output [10:0]t0;
    output n28194;
    output \bit_ctr[3] ;
    output \bit_ctr[4] ;
    input VCC_net;
    input n30584;
    input n30583;
    input n30582;
    input n30581;
    input n30580;
    input n30579;
    input n30578;
    input n30577;
    input n30576;
    input n30555;
    input n30479;
    input n65800;
    output NEOPXL_c;
    output n61457;
    output n61432;
    output \color_bit_N_502[2] ;
    output n44741;
    output n25406;
    input LED_c;
    output n3165;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [10:0]t1_10__N_432;
    wire [10:0]t1;   // verilog/neopixel.v(11[12:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n68956, \neo_pixel_transmitter.done , 
        start_N_507, n66036, start, n79378, n79381, n72530, n72531, 
        n72534, n72533, n72572, n72573, n72609, n72608;
    wire [10:0]n49;
    
    wire n60164, n60163, n60162, n60161, n60160, n60159, n15, 
        n15_adj_5703, n32, n25906, n60158, n22994, n60157, n60156;
    wire [31:0]n149;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(20[11:18])
    
    wire n29446, n60155;
    wire [10:0]n1;
    
    wire n59167, n59166, n59165, n59164, n59163, n59162, n59161, 
        n59160, n59159, n59158, n20530, n28184, n29160;
    wire [1:0]state_1__N_451;
    
    wire n28198, n29448, one_wire_N_499, n44, n69044, n25908, n75333, 
        n68710, n68, n67830, n68958, n53_adj_5704, n44678, n67738, 
        n66803, n72540, n72539, n79255, n72541, n72543, n72544, 
        n81, n79195, n73769, n67802, n25903, n22, n66845, n25, 
        n67826, n8_adj_5705, n45412, n7193, n79252, n67736, n45236, 
        n25863, n28, n75325, n79192, n6_adj_5706, n70003;
    
    SB_DFF t1_i0 (.Q(t1[0]), .C(clk16MHz), .D(t1_10__N_432[0]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n68956), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n66036), .D(start_N_507));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i2201_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(\color_bit_N_502[1] ));   // verilog/neopixel.v(65[23:32])
    defparam i2201_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n79378_bdd_4_lut (.I0(n79378), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(\color_bit_N_502[1] ), .O(n79381));
    defparam n79378_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i56674_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n72530));
    defparam i56674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56675_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n72531));
    defparam i56675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56678_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n72534));
    defparam i56678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56677_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n72533));
    defparam i56677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56716_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n72572));
    defparam i56716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56717_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n72573));
    defparam i56717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56753_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n72609));
    defparam i56753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56752_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n72608));
    defparam i56752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2039_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n60164), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2039_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n60163), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_11 (.CI(n60163), .I0(GND_net), .I1(timer[9]), 
            .CO(n60164));
    SB_LUT4 timer_2039_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n60162), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_10 (.CI(n60162), .I0(GND_net), .I1(timer[8]), 
            .CO(n60163));
    SB_LUT4 timer_2039_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n60161), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_9 (.CI(n60161), .I0(GND_net), .I1(timer[7]), 
            .CO(n60162));
    SB_LUT4 timer_2039_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n60160), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_8 (.CI(n60160), .I0(GND_net), .I1(timer[6]), 
            .CO(n60161));
    SB_LUT4 timer_2039_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n60159), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_4_lut (.I0(n15), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(n15_adj_5703), .O(n32));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h14d7;
    SB_CARRY timer_2039_add_4_7 (.CI(n60159), .I0(GND_net), .I1(timer[5]), 
            .CO(n60160));
    SB_LUT4 i2_3_lut_4_lut (.I0(t1[1]), .I1(t1[0]), .I2(t1[4]), .I3(t1[3]), 
            .O(n25906));   // verilog/neopixel.v(60[15:45])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF timer_2039__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(14[12:21])
    SB_LUT4 timer_2039_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n60158), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_6 (.CI(n60158), .I0(GND_net), .I1(timer[4]), 
            .CO(n60159));
    SB_LUT4 i8808_3_lut_4_lut (.I0(n15), .I1(t1[2]), .I2(n25906), .I3(state[0]), 
            .O(n22994));   // verilog/neopixel.v(35[4] 112[11])
    defparam i8808_3_lut_4_lut.LUT_INIT = 16'hf3aa;
    SB_LUT4 timer_2039_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n60157), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF t0_i0_i0 (.Q(t0[0]), .C(clk16MHz), .D(n29968));   // verilog/neopixel.v(34[12] 113[6])
    SB_CARRY timer_2039_add_4_5 (.CI(n60157), .I0(GND_net), .I1(timer[3]), 
            .CO(n60158));
    SB_LUT4 timer_2039_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n60156), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_4 (.CI(n60156), .I0(GND_net), .I1(timer[2]), 
            .CO(n60157));
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n28194), 
            .D(n149[2]), .R(n29446));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i3 (.Q(\bit_ctr[3] ), .C(clk16MHz), .E(n28194), 
            .D(n149[3]), .R(n29446));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i4 (.Q(\bit_ctr[4] ), .C(clk16MHz), .E(n28194), 
            .D(n149[4]), .R(n29446));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 timer_2039_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n60155), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_3 (.CI(n60155), .I0(GND_net), .I1(timer[1]), 
            .CO(n60156));
    SB_LUT4 timer_2039_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF timer_2039__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(14[12:21])
    SB_CARRY timer_2039_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n60155));
    SB_DFF t0_i0_i1 (.Q(t0[1]), .C(clk16MHz), .D(n30584));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i2 (.Q(t0[2]), .C(clk16MHz), .D(n30583));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i3 (.Q(t0[3]), .C(clk16MHz), .D(n30582));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i4 (.Q(t0[4]), .C(clk16MHz), .D(n30581));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i5 (.Q(t0[5]), .C(clk16MHz), .D(n30580));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i6 (.Q(t0[6]), .C(clk16MHz), .D(n30579));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i7 (.Q(t0[7]), .C(clk16MHz), .D(n30578));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i8 (.Q(t0[8]), .C(clk16MHz), .D(n30577));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i9 (.Q(t0[9]), .C(clk16MHz), .D(n30576));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i10 (.Q(t0[10]), .C(clk16MHz), .D(n30555));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .D(n30479));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n65800));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i2215_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), 
            .I2(bit_ctr[0]), .I3(\bit_ctr[3] ), .O(n149[3]));   // verilog/neopixel.v(65[23:32])
    defparam i2215_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 timer_10__I_0_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n59167), .O(t1_10__N_432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_10__I_0_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n59166), .O(t1_10__N_432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_11 (.CI(n59166), .I0(timer[9]), .I1(n1[9]), 
            .CO(n59167));
    SB_LUT4 timer_10__I_0_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n59165), .O(t1_10__N_432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_10 (.CI(n59165), .I0(timer[8]), .I1(n1[8]), 
            .CO(n59166));
    SB_LUT4 timer_10__I_0_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n59164), .O(t1_10__N_432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_9 (.CI(n59164), .I0(timer[7]), .I1(n1[7]), 
            .CO(n59165));
    SB_LUT4 timer_10__I_0_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n59163), .O(t1_10__N_432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_8 (.CI(n59163), .I0(timer[6]), .I1(n1[6]), 
            .CO(n59164));
    SB_LUT4 timer_10__I_0_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n59162), .O(t1_10__N_432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_7 (.CI(n59162), .I0(timer[5]), .I1(n1[5]), 
            .CO(n59163));
    SB_LUT4 timer_10__I_0_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n59161), .O(t1_10__N_432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_6 (.CI(n59161), .I0(timer[4]), .I1(n1[4]), 
            .CO(n59162));
    SB_LUT4 timer_10__I_0_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n59160), .O(t1_10__N_432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_5 (.CI(n59160), .I0(timer[3]), .I1(n1[3]), 
            .CO(n59161));
    SB_LUT4 timer_10__I_0_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n59159), .O(t1_10__N_432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_4 (.CI(n59159), .I0(timer[2]), .I1(n1[2]), 
            .CO(n59160));
    SB_LUT4 timer_10__I_0_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n1[1]), 
            .I3(n59158), .O(t1_10__N_432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_3 (.CI(n59158), .I0(timer[1]), .I1(n1[1]), 
            .CO(n59159));
    SB_LUT4 timer_10__I_0_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(t1_10__N_432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n59158));
    SB_DFF t1_i10 (.Q(t1[10]), .C(clk16MHz), .D(t1_10__N_432[10]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i9 (.Q(t1[9]), .C(clk16MHz), .D(t1_10__N_432[9]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i8 (.Q(t1[8]), .C(clk16MHz), .D(t1_10__N_432[8]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i7 (.Q(t1[7]), .C(clk16MHz), .D(t1_10__N_432[7]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i6 (.Q(t1[6]), .C(clk16MHz), .D(t1_10__N_432[6]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i5 (.Q(t1[5]), .C(clk16MHz), .D(t1_10__N_432[5]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i4 (.Q(t1[4]), .C(clk16MHz), .D(t1_10__N_432[4]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i3 (.Q(t1[3]), .C(clk16MHz), .D(t1_10__N_432[3]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i2 (.Q(t1[2]), .C(clk16MHz), .D(t1_10__N_432[2]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i1 (.Q(t1[1]), .C(clk16MHz), .D(t1_10__N_432[1]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n28184), .D(n20530), 
            .R(n29160));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n28198), .D(state_1__N_451[0]), 
            .S(n29448));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n44), .D(one_wire_N_499), 
            .R(n69044));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i60402_3_lut (.I0(n25908), .I1(state[0]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n75333));
    defparam i60402_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i72_4_lut (.I0(n68710), .I1(n75333), .I2(state[1]), .I3(start), 
            .O(n68));
    defparam i72_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i63248_4_lut (.I0(n67830), .I1(n68), .I2(n68958), .I3(n53_adj_5704), 
            .O(n44));
    defparam i63248_4_lut.LUT_INIT = 16'h2223;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(one_wire_N_499));
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30589_2_lut (.I0(n25908), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n44678));
    defparam i30589_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut (.I0(start), .I1(n67738), .I2(state[1]), .I3(n66803), 
            .O(n29448));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i56684_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n72540));
    defparam i56684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56683_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n72539));
    defparam i56683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56685_4_lut (.I0(n72540), .I1(n79255), .I2(n61457), .I3(n61432), 
            .O(n72541));
    defparam i56685_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i56687_4_lut (.I0(n72541), .I1(n72539), .I2(n61457), .I3(\color_bit_N_502[1] ), 
            .O(n72543));
    defparam i56687_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i56688_4_lut (.I0(n72543), .I1(n79381), .I2(n61457), .I3(\color_bit_N_502[2] ), 
            .O(n72544));
    defparam i56688_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i30488_4_lut (.I0(n72544), .I1(n81), .I2(n79195), .I3(n73769), 
            .O(state_1__N_451[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i30488_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2208_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n149[2]));   // verilog/neopixel.v(65[23:32])
    defparam i2208_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 timer_10__I_0_inv_0_i1_1_lut (.I0(t0[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_3_lut_4_lut (.I0(t1[6]), .I1(t1[7]), .I2(t1[5]), .I3(t1[8]), 
            .O(n67802));   // verilog/neopixel.v(100[14:42])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_4_lut_adj_1805 (.I0(t1[6]), .I1(t1[7]), .I2(t1[5]), 
            .I3(t1[9]), .O(n25903));   // verilog/neopixel.v(100[14:42])
    defparam i3_3_lut_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i47_3_lut_4_lut_3_lut (.I0(t1[1]), .I1(t1[3]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n22));
    defparam i47_3_lut_4_lut_3_lut.LUT_INIT = 16'h8181;
    SB_LUT4 i3_3_lut_4_lut_adj_1806 (.I0(t1[1]), .I1(t1[3]), .I2(t1[2]), 
            .I3(n66845), .O(n15));
    defparam i3_3_lut_4_lut_adj_1806.LUT_INIT = 16'hff7f;
    SB_LUT4 i46_3_lut_4_lut_3_lut (.I0(t1[1]), .I1(t1[3]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n25));
    defparam i46_3_lut_4_lut_3_lut.LUT_INIT = 16'h1818;
    SB_LUT4 timer_10__I_0_inv_0_i2_1_lut (.I0(t0[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i3_1_lut (.I0(t0[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1807 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n25908), .I3(state[1]), .O(n69044));
    defparam i2_3_lut_4_lut_adj_1807.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_1808 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n67830), .I3(n15_adj_5703), .O(n68710));
    defparam i2_3_lut_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 i52018_2_lut_3_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n25908), .I3(GND_net), .O(n67826));
    defparam i52018_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 timer_10__I_0_inv_0_i4_1_lut (.I0(t0[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i5_1_lut (.I0(t0[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i6_1_lut (.I0(t0[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i7_1_lut (.I0(t0[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i8_1_lut (.I0(t0[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i9_1_lut (.I0(t0[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i10_1_lut (.I0(t0[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i11_1_lut (.I0(t0[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(\bit_ctr[3] ), .I1(n44741), .I2(GND_net), .I3(GND_net), 
            .O(n61432));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut (.I0(\color_bit_N_502[2] ), .I1(n61457), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n8_adj_5705));
    defparam i3_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1174_4_lut (.I0(\color_bit_N_502[1] ), .I1(n45412), .I2(n8_adj_5705), 
            .I3(n61432), .O(n81));   // verilog/neopixel.v(24[26:38])
    defparam i1174_4_lut.LUT_INIT = 16'h3233;
    SB_LUT4 i2203_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n7193));   // verilog/neopixel.v(65[23:32])
    defparam i2203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15233_2_lut (.I0(n28194), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n29446));   // verilog/neopixel.v(34[12] 113[6])
    defparam i15233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(\color_bit_N_502[1] ), .I1(n72608), 
            .I2(n72609), .I3(\color_bit_N_502[2] ), .O(n79252));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n79252_bdd_4_lut (.I0(n79252), .I1(n72573), .I2(n72572), .I3(\color_bit_N_502[2] ), 
            .O(n79255));
    defparam n79252_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i57913_2_lut_3_lut (.I0(n61457), .I1(\bit_ctr[3] ), .I2(n44741), 
            .I3(GND_net), .O(n73769));   // verilog/neopixel.v(24[26:38])
    defparam i57913_2_lut_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i51931_2_lut_3_lut (.I0(n25908), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n67738));
    defparam i51931_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1809 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(t1[2]), .I3(n25906), .O(n68958));
    defparam i2_3_lut_4_lut_adj_1809.LUT_INIT = 16'h0080;
    SB_LUT4 i52022_2_lut_3_lut (.I0(t1[10]), .I1(t1[9]), .I2(n67802), 
            .I3(GND_net), .O(n67830));
    defparam i52022_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_4_lut_adj_1810 (.I0(n25406), .I1(state[1]), .I2(n44678), 
            .I3(state[0]), .O(n28198));
    defparam i1_4_lut_4_lut_adj_1810.LUT_INIT = 16'hee2e;
    SB_LUT4 i1_2_lut_3_lut (.I0(n25406), .I1(state[1]), .I2(n28184), .I3(GND_net), 
            .O(n28194));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n28184));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h20ff;
    SB_LUT4 i51929_2_lut (.I0(t1[10]), .I1(t1[9]), .I2(GND_net), .I3(GND_net), 
            .O(n67736));
    defparam i51929_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i31147_2_lut (.I0(state[1]), .I1(t1[0]), .I2(GND_net), .I3(GND_net), 
            .O(n45236));
    defparam i31147_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14946_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n29160));   // verilog/neopixel.v(35[4] 112[11])
    defparam i14946_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i6672_3_lut_4_lut (.I0(start), .I1(n25863), .I2(n22994), .I3(bit_ctr[0]), 
            .O(n20530));
    defparam i6672_3_lut_4_lut.LUT_INIT = 16'hfb04;
    SB_LUT4 i1_4_lut (.I0(n45236), .I1(n25), .I2(state[0]), .I3(n22), 
            .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h4540;
    SB_LUT4 i60269_4_lut (.I0(n67802), .I1(t1[2]), .I2(n28), .I3(t1[4]), 
            .O(n75325));
    defparam i60269_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_3_lut_adj_1811 (.I0(start), .I1(n25863), .I2(n22994), 
            .I3(GND_net), .O(n25406));
    defparam i1_2_lut_3_lut_adj_1811.LUT_INIT = 16'h0404;
    SB_LUT4 i45_4_lut (.I0(n75325), .I1(state[1]), .I2(start), .I3(n67736), 
            .O(n3165));
    defparam i45_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i1_2_lut_3_lut_adj_1812 (.I0(\bit_ctr[3] ), .I1(n44741), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n61457));
    defparam i1_2_lut_3_lut_adj_1812.LUT_INIT = 16'h7878;
    SB_LUT4 i31318_2_lut_3_lut (.I0(\bit_ctr[3] ), .I1(n44741), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n45412));
    defparam i31318_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i30652_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n44741));
    defparam i30652_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1813 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(\color_bit_N_502[2] ));
    defparam i1_2_lut_3_lut_adj_1813.LUT_INIT = 16'h1e1e;
    SB_LUT4 i2222_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n7193), .I2(\bit_ctr[3] ), 
            .I3(\bit_ctr[4] ), .O(n149[4]));   // verilog/neopixel.v(65[23:32])
    defparam i2222_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_63368 (.I0(\color_bit_N_502[1] ), 
            .I1(n72533), .I2(n72534), .I3(\color_bit_N_502[2] ), .O(n79192));
    defparam color_bit_N_502_1__bdd_4_lut_63368.LUT_INIT = 16'he4aa;
    SB_LUT4 n79192_bdd_4_lut (.I0(n79192), .I1(n72531), .I2(n72530), .I3(\color_bit_N_502[2] ), 
            .O(n79195));
    defparam n79192_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n79378));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i3_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n25903), .I2(t1[10]), 
            .I3(t1[8]), .O(n25863));
    defparam i3_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_adj_1814 (.I0(n22994), .I1(n25863), .I2(GND_net), 
            .I3(GND_net), .O(n66803));   // verilog/neopixel.v(34[12] 113[6])
    defparam i1_2_lut_adj_1814.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1815 (.I0(n25903), .I1(t1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5706));   // verilog/neopixel.v(100[14:42])
    defparam i1_2_lut_adj_1815.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut (.I0(t1[10]), .I1(n25906), .I2(t1[2]), .I3(n6_adj_5706), 
            .O(n25908));   // verilog/neopixel.v(100[14:42])
    defparam i4_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i22_4_lut (.I0(n66803), .I1(n67826), .I2(state[1]), .I3(start), 
            .O(n66036));
    defparam i22_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i62446_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 112[11])
    defparam i62446_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1816 (.I0(t1[0]), .I1(t1[4]), .I2(GND_net), .I3(GND_net), 
            .O(n66845));
    defparam i1_2_lut_adj_1816.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1817 (.I0(t1[2]), .I1(n25906), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5703));   // verilog/neopixel.v(60[15:45])
    defparam i1_2_lut_adj_1817.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(n15), .I1(\neo_pixel_transmitter.done ), .I2(state[0]), 
            .I3(GND_net), .O(n53_adj_5704));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i3_4_lut_adj_1818 (.I0(n25903), .I1(n32), .I2(t1[10]), .I3(t1[8]), 
            .O(n70003));
    defparam i3_4_lut_adj_1818.LUT_INIT = 16'h0004;
    SB_LUT4 i2_3_lut (.I0(state[1]), .I1(n70003), .I2(start), .I3(GND_net), 
            .O(n68956));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 state_1__I_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(35[4] 112[11])
    defparam state_1__I_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (\a_new[1] , \b_new[1] , debounce_cnt_N_3833, 
            a_prev, b_prev, position_31__N_3836, GND_net, ENCODER0_B_N_keep, 
            n1779, ENCODER0_A_N_keep, n30012, n1742, n30008, n29986, 
            n1744, \encoder0_position[30] , \encoder0_position[29] , \encoder0_position[28] , 
            \encoder0_position[27] , \encoder0_position[26] , \encoder0_position[25] , 
            \encoder0_position[24] , \encoder0_position[23] , \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            \encoder0_position[18] , \encoder0_position[17] , \encoder0_position[16] , 
            \encoder0_position[15] , \encoder0_position[14] , \encoder0_position[13] , 
            \encoder0_position[12] , \encoder0_position[11] , \encoder0_position[10] , 
            \encoder0_position[9] , \encoder0_position[8] , \encoder0_position[7] , 
            \encoder0_position[6] , \encoder0_position[5] , \encoder0_position[4] , 
            \encoder0_position[3] , \encoder0_position[2] , \encoder0_position[1] , 
            \encoder0_position[0] , VCC_net) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    output \b_new[1] ;
    output debounce_cnt_N_3833;
    output a_prev;
    output b_prev;
    output position_31__N_3836;
    input GND_net;
    input ENCODER0_B_N_keep;
    input n1779;
    input ENCODER0_A_N_keep;
    input n30012;
    output n1742;
    input n30008;
    input n29986;
    output n1744;
    output \encoder0_position[30] ;
    output \encoder0_position[29] ;
    output \encoder0_position[28] ;
    output \encoder0_position[27] ;
    output \encoder0_position[26] ;
    output \encoder0_position[25] ;
    output \encoder0_position[24] ;
    output \encoder0_position[23] ;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire direction_N_3840;
    wire [31:0]n133;
    
    wire n60320, n60319, n60318, n60317, n60316, n60315, n60314, 
        n60313, n60312, n60311, n60310, n60309, n60308, n60307, 
        n60306, n60305, n60304, n60303, n60302, n60301, n60300, 
        n60299, n60298, n60297, n60296, n60295, n60294, n60293, 
        n60292, n60291, n60290;
    
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1742), .C(n1779), .D(n30012));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n30008));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29986));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2054__i31 (.Q(n1744), .C(n1779), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i30 (.Q(\encoder0_position[30] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i29 (.Q(\encoder0_position[29] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i28 (.Q(\encoder0_position[28] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i27 (.Q(\encoder0_position[27] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i26 (.Q(\encoder0_position[26] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i25 (.Q(\encoder0_position[25] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i24 (.Q(\encoder0_position[24] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i23 (.Q(\encoder0_position[23] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i22 (.Q(\encoder0_position[22] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i21 (.Q(\encoder0_position[21] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i20 (.Q(\encoder0_position[20] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i19 (.Q(\encoder0_position[19] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i18 (.Q(\encoder0_position[18] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i17 (.Q(\encoder0_position[17] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i16 (.Q(\encoder0_position[16] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i15 (.Q(\encoder0_position[15] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i14 (.Q(\encoder0_position[14] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i13 (.Q(\encoder0_position[13] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i12 (.Q(\encoder0_position[12] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i11 (.Q(\encoder0_position[11] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i10 (.Q(\encoder0_position[10] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i9 (.Q(\encoder0_position[9] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i8 (.Q(\encoder0_position[8] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i7 (.Q(\encoder0_position[7] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i6 (.Q(\encoder0_position[6] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i5 (.Q(\encoder0_position[5] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i4 (.Q(\encoder0_position[4] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i3 (.Q(\encoder0_position[3] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i2 (.Q(\encoder0_position[2] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i1 (.Q(\encoder0_position[1] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i0 (.Q(\encoder0_position[0] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2054_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1744), .I3(n60320), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2054_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[30] ), .I3(n60319), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_32 (.CI(n60319), .I0(direction_N_3840), 
            .I1(\encoder0_position[30] ), .CO(n60320));
    SB_LUT4 position_2054_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[29] ), .I3(n60318), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_31 (.CI(n60318), .I0(direction_N_3840), 
            .I1(\encoder0_position[29] ), .CO(n60319));
    SB_LUT4 position_2054_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[28] ), .I3(n60317), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_30 (.CI(n60317), .I0(direction_N_3840), 
            .I1(\encoder0_position[28] ), .CO(n60318));
    SB_LUT4 position_2054_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[27] ), .I3(n60316), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_29 (.CI(n60316), .I0(direction_N_3840), 
            .I1(\encoder0_position[27] ), .CO(n60317));
    SB_LUT4 position_2054_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[26] ), .I3(n60315), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_28 (.CI(n60315), .I0(direction_N_3840), 
            .I1(\encoder0_position[26] ), .CO(n60316));
    SB_LUT4 position_2054_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[25] ), .I3(n60314), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_27 (.CI(n60314), .I0(direction_N_3840), 
            .I1(\encoder0_position[25] ), .CO(n60315));
    SB_LUT4 position_2054_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[24] ), .I3(n60313), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_26 (.CI(n60313), .I0(direction_N_3840), 
            .I1(\encoder0_position[24] ), .CO(n60314));
    SB_LUT4 position_2054_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[23] ), .I3(n60312), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_25 (.CI(n60312), .I0(direction_N_3840), 
            .I1(\encoder0_position[23] ), .CO(n60313));
    SB_LUT4 position_2054_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[22] ), .I3(n60311), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_24 (.CI(n60311), .I0(direction_N_3840), 
            .I1(\encoder0_position[22] ), .CO(n60312));
    SB_LUT4 position_2054_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[21] ), .I3(n60310), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_23 (.CI(n60310), .I0(direction_N_3840), 
            .I1(\encoder0_position[21] ), .CO(n60311));
    SB_LUT4 position_2054_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[20] ), .I3(n60309), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_22 (.CI(n60309), .I0(direction_N_3840), 
            .I1(\encoder0_position[20] ), .CO(n60310));
    SB_LUT4 position_2054_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[19] ), .I3(n60308), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_21 (.CI(n60308), .I0(direction_N_3840), 
            .I1(\encoder0_position[19] ), .CO(n60309));
    SB_LUT4 position_2054_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[18] ), .I3(n60307), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_20 (.CI(n60307), .I0(direction_N_3840), 
            .I1(\encoder0_position[18] ), .CO(n60308));
    SB_LUT4 position_2054_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[17] ), .I3(n60306), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_19 (.CI(n60306), .I0(direction_N_3840), 
            .I1(\encoder0_position[17] ), .CO(n60307));
    SB_LUT4 position_2054_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[16] ), .I3(n60305), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_18 (.CI(n60305), .I0(direction_N_3840), 
            .I1(\encoder0_position[16] ), .CO(n60306));
    SB_LUT4 position_2054_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[15] ), .I3(n60304), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_17 (.CI(n60304), .I0(direction_N_3840), 
            .I1(\encoder0_position[15] ), .CO(n60305));
    SB_LUT4 position_2054_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[14] ), .I3(n60303), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_16 (.CI(n60303), .I0(direction_N_3840), 
            .I1(\encoder0_position[14] ), .CO(n60304));
    SB_LUT4 position_2054_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[13] ), .I3(n60302), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_15 (.CI(n60302), .I0(direction_N_3840), 
            .I1(\encoder0_position[13] ), .CO(n60303));
    SB_LUT4 position_2054_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[12] ), .I3(n60301), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_14 (.CI(n60301), .I0(direction_N_3840), 
            .I1(\encoder0_position[12] ), .CO(n60302));
    SB_LUT4 position_2054_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[11] ), .I3(n60300), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_13 (.CI(n60300), .I0(direction_N_3840), 
            .I1(\encoder0_position[11] ), .CO(n60301));
    SB_LUT4 position_2054_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[10] ), .I3(n60299), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_12 (.CI(n60299), .I0(direction_N_3840), 
            .I1(\encoder0_position[10] ), .CO(n60300));
    SB_LUT4 position_2054_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[9] ), .I3(n60298), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_11 (.CI(n60298), .I0(direction_N_3840), 
            .I1(\encoder0_position[9] ), .CO(n60299));
    SB_LUT4 position_2054_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[8] ), .I3(n60297), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_10 (.CI(n60297), .I0(direction_N_3840), 
            .I1(\encoder0_position[8] ), .CO(n60298));
    SB_LUT4 position_2054_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[7] ), .I3(n60296), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_9 (.CI(n60296), .I0(direction_N_3840), 
            .I1(\encoder0_position[7] ), .CO(n60297));
    SB_LUT4 position_2054_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[6] ), .I3(n60295), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_8 (.CI(n60295), .I0(direction_N_3840), 
            .I1(\encoder0_position[6] ), .CO(n60296));
    SB_LUT4 position_2054_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[5] ), .I3(n60294), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_7 (.CI(n60294), .I0(direction_N_3840), 
            .I1(\encoder0_position[5] ), .CO(n60295));
    SB_LUT4 position_2054_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[4] ), .I3(n60293), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_6 (.CI(n60293), .I0(direction_N_3840), 
            .I1(\encoder0_position[4] ), .CO(n60294));
    SB_LUT4 position_2054_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[3] ), .I3(n60292), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_5 (.CI(n60292), .I0(direction_N_3840), 
            .I1(\encoder0_position[3] ), .CO(n60293));
    SB_LUT4 position_2054_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[2] ), .I3(n60291), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_4 (.CI(n60291), .I0(direction_N_3840), 
            .I1(\encoder0_position[2] ), .CO(n60292));
    SB_LUT4 position_2054_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[1] ), .I3(n60290), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_3 (.CI(n60290), .I0(direction_N_3840), 
            .I1(\encoder0_position[1] ), .CO(n60291));
    SB_LUT4 position_2054_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n60290));
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, IntegralLimit, \Kp[4] , n20421, \Kp[5] , 
            PWMLimit, n284, \Kp[2] , \Kp[3] , \Kp[7] , \Kp[6] , 
            \Kp[8] , \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , n258, 
            n356, \Ki[1] , n357, \Ki[0] , n339, \Ki[2] , \Ki[3] , 
            n239, \Kp[13] , \Kp[14] , \Ki[4] , \Ki[5] , \Kp[15] , 
            \Ki[6] , n346, \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , 
            \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , n358, 
            n20422, n299, control_update, duty, clk16MHz, reset, 
            n56, setpoint, \motor_state[9] , n340, VCC_net, \motor_state[8] , 
            n359, \motor_state[7] , \PID_CONTROLLER.integral , n336, 
            \motor_state[6] , \motor_state[5] , n21, n460, n461, n467, 
            n475, n462, n247, n37, n9, n16, n34689, n20, n291, 
            n25, n35, n33, n37_adj_27, n41, n22, n105, n35782, 
            n24, n36147, n36361, \motor_state[4] , n25921, n4, n342, 
            n337, n37307, n37117, n137, n347, n6, \Kp[1] , \Kp[0] , 
            deadband, n8, n25_adj_28, n343, n10, n34, n38, n40, 
            n38_adj_29, n36, n75815, n24_adj_30, n30516, n30515, 
            n30514, n30513, n30512, n30511, n30510, n30509, n30508, 
            n30507, n30505, n30503, n30502, n30501, n30500, n30499, 
            n30498, n30497, n30496, n30495, n30490, n30489, n30481, 
            n29775, n347_adj_31, \control_mode[0] , n53108, \control_mode[1] , 
            n28076, n344, n348, n17, n45282, \motor_state[2] , \motor_state[1] , 
            \motor_state[0] , n349, \motor_state[23] , n38_adj_32, \motor_state[22] , 
            n350, \motor_state[21] , n345, n12, \motor_state[19] , 
            \motor_state[18] , \motor_state[17] , n486, n351, n110, 
            \motor_state[16] , \motor_state[15] , \motor_state[14] , \motor_state[13] , 
            n10_adj_33, n42994, \motor_state[10] , n352, n353, n354, 
            n58586, n322, n20467, n20468, n355, n313) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [23:0]IntegralLimit;
    input \Kp[4] ;
    input n20421;
    input \Kp[5] ;
    input [23:0]PWMLimit;
    output n284;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[7] ;
    input \Kp[6] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    output n258;
    output n356;
    input \Ki[1] ;
    output n357;
    input \Ki[0] ;
    output n339;
    input \Ki[2] ;
    input \Ki[3] ;
    output n239;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Kp[15] ;
    input \Ki[6] ;
    output n346;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    output n358;
    input n20422;
    output n299;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input n56;
    input [23:0]setpoint;
    input \motor_state[9] ;
    output n340;
    input VCC_net;
    input \motor_state[8] ;
    output n359;
    input \motor_state[7] ;
    output [23:0]\PID_CONTROLLER.integral ;
    output n336;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input n21;
    output n460;
    output n461;
    output n467;
    output n475;
    output n462;
    output n247;
    input n37;
    input n9;
    output n16;
    input n34689;
    output n20;
    output n291;
    input n25;
    input n35;
    input n33;
    input n37_adj_27;
    input n41;
    input n22;
    output n105;
    input n35782;
    output n24;
    input n36147;
    input n36361;
    input \motor_state[4] ;
    input n25921;
    input n4;
    output n342;
    output n337;
    input n37307;
    input n37117;
    input n137;
    input n347;
    input n6;
    input \Kp[1] ;
    input \Kp[0] ;
    input [23:0]deadband;
    output n8;
    input n25_adj_28;
    output n343;
    input n10;
    output n34;
    output n38;
    input n40;
    input n38_adj_29;
    input n36;
    input n75815;
    input n24_adj_30;
    input n30516;
    input n30515;
    input n30514;
    input n30513;
    input n30512;
    input n30511;
    input n30510;
    input n30509;
    input n30508;
    input n30507;
    input n30505;
    input n30503;
    input n30502;
    input n30501;
    input n30500;
    input n30499;
    input n30498;
    input n30497;
    input n30496;
    input n30495;
    input n30490;
    input n30489;
    input n30481;
    input n29775;
    input n347_adj_31;
    input \control_mode[0] ;
    input n53108;
    input \control_mode[1] ;
    output n28076;
    output n344;
    output n348;
    input n17;
    output n45282;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input \motor_state[0] ;
    input n349;
    input \motor_state[23] ;
    input n38_adj_32;
    input \motor_state[22] ;
    output n350;
    input \motor_state[21] ;
    output n345;
    input n12;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    output n486;
    output n351;
    input n110;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input n10_adj_33;
    input n42994;
    input \motor_state[10] ;
    output n352;
    output n353;
    output n354;
    output n58586;
    output n322;
    output n20467;
    output n20468;
    output n355;
    output n313;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n59067;
    wire [23:0]n1;
    
    wire n59068, n16_c;
    wire [23:0]n233;
    
    wire n45, n24_c, n43, n25_c, n23, n76006, n75962, n59275;
    wire [4:0]n20418;
    
    wire n417, n59276;
    wire [23:0]n285;
    
    wire n59066, n8_c, n75960, n77553, n77724, n76463, n4_c;
    wire [23:0]n207;
    
    wire n335;
    wire [5:0]n20350;
    
    wire n344_c, n59274, n59065, n58957;
    wire [43:0]n360;
    wire [47:0]n46;
    
    wire n58958, n408, n5076, n75265;
    wire [23:0]n310;
    
    wire n183, n256_adj_5136, n329, n512, n402, n475_c, n585, 
        n658, n548, n731, n804, n75266, n621, n877, n694, n27, 
        n77721, n767, n840, n80, n11_adj_5137, n29, n77722, n153, 
        n226, n33_c, n31, n75992, n75980, n30, n10_c, n35_c, 
        n75976, n78065, n76465, n78219, n37_c, n78220, n39, n78188, 
        n41_c, n78132, n75964, n78042, n950, n1023, n299_c, n372, 
        n1096, n445, n76471, n186, n518, n591, n664, n737, n810, 
        n883, n956, n1029, n1102, n259, n77, n8_adj_5138, n150, 
        n223, n332_adj_5139, n296_adj_5140, n369, n442, n59064, 
        n271, n59273, n78044, n59063, n198, n59272;
    wire [13:0]n61;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n60269, n515, n60268, n79225, counter_31__N_3714, n588, 
        n60267, n125, n59062, n75264;
    wire [23:0]n455;
    
    wire n58956, n661, n60266, n734, n60265;
    wire [12:0]n18700;
    wire [11:0]n19063;
    
    wire n980, n59271, n907, n59270, n58916, n60264, n60263, n59061, 
        n807, n60262, n880, n60261, n60260, n953, n60259, n1026, 
        n834, n59269, n60258, n1099, n761, n59268, n59060, n60257, 
        n59059, n58955, n59058, n688, n59267, n615, n59266, n542, 
        n59265, n59057, n469, n59264, n396, n59263, n59056, n58954, 
        n58917, n59055, n75274, n58915, n323, n59262, n250, n59261, 
        n177, n59260, n74_adj_5146, n5, n147, n220, n59054, n35_adj_5148, 
        n104, n293, n366, n439, n58914, n512_adj_5149, n58953, 
        n585_adj_5151, n58952, n658_adj_5152, n731_adj_5153, n804_adj_5154, 
        n877_adj_5155, n950_adj_5156, n1023_adj_5157, n1096_adj_5158, 
        n481, n58951, n11882, n75285, n4736, n79384, n21_adj_5159, 
        n19_adj_5160, n17_adj_5161, n9_c, n79537, n15_adj_5162, n13_adj_5163, 
        n11_adj_5164, n12_adj_5166, n79501, n79495, n79489, n58950, 
        n79483;
    wire [23:0]n535;
    
    wire n79387, n79477, n79471, n79465, n58949, n58948, n58947, 
        n58913, n45_adj_5167, n39_adj_5168, n41_adj_5169, n58946, 
        n58912, n58945, n76024, n76955, n43_adj_5171, n33_adj_5173, 
        n35_adj_5174, n554, n58944, n27_adj_5175, n76949, n29_adj_5176, 
        n31_adj_5177, n19_adj_5179, n17_adj_5180, n9_adj_5181, n75944, 
        n405, n58943, n15_adj_5182, n13_adj_5183, n11_adj_5184, n75934, 
        n77994, n41_adj_5185, n39_adj_5186, n45_adj_5187, n77407, 
        n12_adj_5188, n29_adj_5189, n31_adj_5190, n43_adj_5191, n37_adj_5192, 
        n10_adj_5193, n30_adj_5194, n17_adj_5195, n19_adj_5196, n21_adj_5198, 
        n23_adj_5200, n25_adj_5201, n75956, n76895, n76889, n9_adj_5203, 
        n25_adj_5204, n23_adj_5205, n77980, n35_adj_5207, n41_adj_5208, 
        n39_adj_5209, n45_adj_5210, n43_adj_5211, n29_adj_5212, n31_adj_5213, 
        n6_c, n77723, n37_adj_5214, n23_adj_5215, n79348, n79351, 
        n25_adj_5216, n35_adj_5217, n9_adj_5218, n17_adj_5219, n19_adj_5220, 
        n21_adj_5221, n33_adj_5222, n43_adj_5223, n77379, n39_adj_5224, 
        n78128, n4_adj_5226, n6_adj_5227, n8_adj_5229, n76188, n78059, 
        n78060, n16_adj_5230, n77951, n79324, n79327, n79321, n79315, 
        n58942, n627, n75259, n31_adj_5233, n700, n478_adj_5234, 
        n6_adj_5235, n77717, n77718, n8_adj_5236, n24_adj_5237, n75900, 
        n75894, n77555, n76473, n4_adj_5238, n77715, n77716, n75923, 
        n75919, n78067, n76475, n78221, n78222, n78186, n75904, 
        n27_adj_5239, n29_adj_5240, n23_adj_5241, n76169, n76158, 
        n551_adj_5245, n28, n30_adj_5246, n26, n34_c, n24_adj_5248, 
        n76154, n78061, n78062, n77947, n77801, n76162, n77978, 
        n76451, n78124, n78125, n11_adj_5252, n13_adj_5253, n15_adj_5254, 
        n27_adj_5255, n37_adj_5256, n15_adj_5257, n13_adj_5258, n19_adj_5259, 
        n17_adj_5260, n7, n11_adj_5261, n5_adj_5262, n75716, n8_adj_5263, 
        n6_adj_5264, n16_adj_5265, n4_adj_5266, n77287, n77288, n75710, 
        n75702, n77874, n76497, n78235, n78236, n41_adj_5268, n29_adj_5269, 
        n31_adj_5270, n33_adj_5271, n39_adj_5272, n27_adj_5273, n75686, 
        n30_adj_5274, n28_adj_5275, n38_c, n79309, n77285, n77286, 
        n58911, n75677, n75675, n77930, n76499, n78183, n78184, 
        n78119, n508, n44726, n25756, n79318, n78046, n76084, 
        n76058, n79303, n12_adj_5277, n79297, n10_adj_5278, n30_adj_5279, 
        n79291, n76116, n77023, n77013, n76481, n78006, n77439, 
        n78136, n16_adj_5280, n79285, n6_adj_5281, n77731, n77732, 
        n79279, n79273, n78048, n8_adj_5282, n79267, n24_adj_5283, 
        n79261, n76032;
    wire [0:0]n12498;
    wire [21:0]n13005;
    
    wire n60586, n60585, n60584, n76026, n77551, n76453, n60583, 
        n60582, n60581, n60580, n4_adj_5284, n77729, n77730, n60579, 
        n76048, n60578, n60577, n75241, n60576, n76044, n78063, 
        n60575, n60574, n60573, n60572, n75254, n76455, n78217, 
        n60571, n60570, n75287, n75288, n78218, n60569, n75255, 
        n75289, n60568, n60567, n75256, n60566, n75291, n75292, 
        n75257, n60565, n75293, n75294;
    wire [20:0]n13970;
    
    wire n60564, n60563, n60562, n60561, n60560, n78190, n76034, 
        n78038;
    wire [0:0]n11922;
    wire [21:0]n12381;
    
    wire n59643, n60559, n59642, n76461;
    wire [2:0]n20492;
    
    wire n4_adj_5288, n277;
    wire [3:0]n20464;
    
    wire n75258, n60558, n60557, n60556, n60555, n490, n71504, 
        n59641, n71508, n78040, n71506, n60554, n131, n71512, 
        n60553, n33_adj_5289, n60552, n11_adj_5290, n4_adj_5291, n68_adj_5292, 
        n71516, n13_adj_5293, n71518, n60551, n79312, n59640, n60550, 
        n60549, n69694, n60548, n60547, n60546, n60545, n15_adj_5295, 
        n60544;
    wire [19:0]n14848;
    
    wire n60543, n60542, n101, n32, n174, n59639, n247_adj_5296, 
        n320, n60541, n393, n27_adj_5297, n21_adj_5298, n59638, 
        n4_adj_5299, n60540, n466_adj_5300, n59637, n539_adj_5301, 
        n60539, n77557, n612, n60538, n685, n19_adj_5305, n23_adj_5306, 
        n60537, n60536, n13_adj_5308, n60535, n60534, n60533, n60532, 
        n758, n59636, n60531, n831, n904, n60530, n60529, n15_adj_5311, 
        n60528, n59635, n977, n1050, n17_adj_5314, n11_adj_5315, 
        n75878, n60527, n60526, n59634, n58941, n59633, n98, n60525, 
        n60524, n58940, n14_adj_5316, n29_adj_5317;
    wire [10:0]n19374;
    wire [9:0]n19637;
    
    wire n60523, n60522, n171, n244_adj_5318, n12_adj_5319, n60521, 
        n59632, n317, n60520, n22_adj_5321, n16_adj_5322, n390_adj_5323, 
        n463_adj_5324, n59631, n536_adj_5326, n59630, n60519, n609, 
        n59629, n682, n59628, n60518, n755, n60517, n59627, n828, 
        n60516, n901, n974, n60515, n1047, n60514, n1120, n122, 
        n53, n41_adj_5328, n110_c, n195;
    wire [18:0]n15644;
    
    wire n60513, n60512, n18_adj_5329, n45309;
    wire [23:0]n1_adj_5701;
    
    wire n60511, n75862, n75857, n78069, n268, n60510, n75864, 
        n77559;
    wire [1:0]n20501;
    
    wire n341, n60509, n414, n1105, n60508, n58939, n487, n78229, 
        n78230, n1032, n60507, n560, n78175, n959, n60506, n886, 
        n60505, n77561, n813, n60504, n41_adj_5335;
    wire [23:0]n48;
    
    wire n23_adj_5336, n740, n60503, n25_adj_5340, n667, n60502, 
        n75263, n79306, n594, n60501, n521, n60500, n448_adj_5342, 
        n60499, n17_adj_5343, n375, n60498, n302_adj_5344, n60497, 
        n75262, n79300, n19_adj_5345, n21_adj_5346, n229, n60496, 
        n7_adj_5347, n156, n60495, n14_adj_5348, n83;
    wire [17:0]n16362;
    
    wire n60494, n60493, n9_adj_5349, n60492, n60491, n11_adj_5350, 
        n1108, n60490, n13_adj_5351, n1035, n60489, n962, n60488, 
        n889, n60487, n816, n60486, n743, n60485, n15_adj_5352, 
        n670, n60484, n597, n60483, n524, n60482, n451_adj_5353, 
        n60481, n378, n60480, n305_adj_5354, n60479, n27_adj_5355, 
        n232, n60478, n439_adj_5356, n59626, n159, n60477, n17_adj_5357, 
        n86;
    wire [8:0]n19856;
    
    wire n770, n60476, n697, n60475, n624, n60474, n35_adj_5358, 
        n551_adj_5359, n60473, n478_adj_5360, n60472, n405_adj_5361, 
        n60471, n29_adj_5362, n332_adj_5363, n60470, n259_adj_5364, 
        n60469, n186_adj_5365, n60468, n44, n113, n75261, n79294, 
        n366_adj_5366, n59625;
    wire [16:0]n17006;
    
    wire n60467, n31_adj_5368, n60466, n60465, n33_adj_5369, n75744, 
        n1111, n60464, n1038, n60463, n293_adj_5370, n59624, n965, 
        n60462, n892, n60461, n819, n60460, n746, n60459, n673, 
        n60458, n600, n60457, n527, n60456, n454, n60455, n381, 
        n60454, n308_adj_5371, n60453, n235_adj_5372, n60452, n162, 
        n60451, n76743, n77299, n77293, n20_adj_5373, n89, n75746, 
        n12_adj_5374, n75139, n4_adj_5375, n77289;
    wire [15:0]n17580;
    
    wire n60450, n77290, n60449, n220_adj_5376, n59623, n1114, n60448, 
        n10_adj_5377, n1041, n60447, n968, n60446, n895, n60445, 
        n30_adj_5378, n822, n60444, n75738, n75735, n77563, n749, 
        n60443, n58938, n676, n60442, n76495, n603, n60441, n147_adj_5379, 
        n59622, n5_adj_5380, n74_adj_5381, n530, n60440, n8_adj_5382, 
        n6_adj_5383, n16_adj_5384, n75760, n77882, n77883, n77706, 
        n77699, n78050, n76493, n78052, n42, n75730, n79794, n44_adj_5387, 
        n77565, n457_adj_5388, n60439;
    wire [9:0]n19778;
    wire [8:0]n19974;
    
    wire n770_adj_5389, n59621, n697_adj_5390, n59620, n384_adj_5391, 
        n60438, n311_adj_5392, n60437, n40_adj_5394, n78071, n624_adj_5395, 
        n59619, n238_adj_5396, n60436, n78072, n47, n77566, n77935, 
        n95, n26_adj_5398, n165, n60435, n23_adj_5399, n92, n75260, 
        n79288, n59618, n168, n59617;
    wire [7:0]n20035;
    
    wire n60434, n79282, n241_adj_5400, n314_adj_5401, n387_adj_5402, 
        n67768, n60433, n460_adj_5404, n533, n606, n75624, n679, 
        n12_adj_5408, n10_adj_5409, n125_adj_5410, n59616, n56_adj_5411, 
        n30_adj_5412, n60432, n752, n75664, n76576, n60431, n59615, 
        n59614, n59613, n825, n76572, n60430, n60429, n898, n198_adj_5413, 
        n77878, n262, n60428, n271_adj_5415, n44_adj_5416, n113_adj_5417, 
        n4_adj_5418, n71550, n189, n60427, n77233, n344_adj_5419, 
        n47_adj_5420, n116;
    wire [2:0]n20470;
    
    wire n4_adj_5421;
    wire [4:0]n20372;
    
    wire n417_adj_5422, n347_adj_5423;
    wire [14:0]n18088;
    
    wire n60426, n6_adj_5424, n67007, n971, n1044, n78099, n1117, 
        n60425, n1117_adj_5425, n16_adj_5426, n71546, n58648, n69342, 
        n62_adj_5427, n6_adj_5428, n77281, n490_adj_5429, n71536, 
        n80190, n71540, n8_adj_5430, n6_adj_5431, n69227, n1044_adj_5432, 
        n60424, n971_adj_5433, n60423, n77282, n75630, n898_adj_5434, 
        n60422, n825_adj_5435, n60421, n752_adj_5436, n60420, n679_adj_5437, 
        n60419, n606_adj_5438, n60418, n533_adj_5439, n60417, n460_adj_5440, 
        n60416, n387_adj_5441, n60415, n314_adj_5442, n60414;
    wire [20:0]n13443;
    
    wire n59590, n59589, n59588, n59587, n59586, n59585, n79249, 
        n8_adj_5443, n59584, n1099_adj_5444, n59583, n1026_adj_5445, 
        n59582, n953_adj_5446, n59581, n24_adj_5447, n75590, n75576, 
        n77569, n76507, n880_adj_5448, n59580, n4_adj_5449, n807_adj_5450, 
        n59579, n734_adj_5451, n59578, n661_adj_5452, n59577, n77277, 
        n588_adj_5453, n59576, n515_adj_5454, n59575, n77278, n442_adj_5455, 
        n59574, n369_adj_5456, n59573, n241_adj_5457, n60413, n296_adj_5458, 
        n59572, n223_adj_5459, n59571, n75613, n75609, n77928, n76509, 
        n150_adj_5460, n59570, n8_adj_5461, n77_adj_5462, n168_adj_5463, 
        n60412;
    wire [19:0]n14367;
    
    wire n59569, n59568, n59567, n910, n59178, n78145, n78146, 
        n78117, n75593, n59566, n837, n59177, n59565, n764, n59176, 
        n59564, n691, n59175, n1102_adj_5464, n59563, n26_adj_5465, 
        n95_adj_5466, n77845, n76515, n78053, n4_adj_5467, n69256, 
        n1029_adj_5468, n59562, n956_adj_5469, n59561;
    wire [13:0]n18534;
    
    wire n1120_adj_5470, n60411, n1047_adj_5471, n60410, n883_adj_5472, 
        n59560, n810_adj_5473, n59559, n618, n59174, n737_adj_5474, 
        n59558, n545_adj_5475, n59173, n664_adj_5476, n59557, n472_adj_5477, 
        n59172, n591_adj_5478, n59556, n399_adj_5479, n59171, n974_adj_5480, 
        n60409, n901_adj_5481, n60408, n518_adj_5482, n59555, n326, 
        n59170, n445_adj_5483, n59554, n253_adj_5484, n59169, n372_adj_5485, 
        n59553, n180, n59168, n299_adj_5486, n59552, n38_adj_5487, 
        n107, n41_adj_5488, n183_adj_5490, n226_adj_5491, n59551, 
        n153_adj_5492, n59550, n11_adj_5493, n80_adj_5494, n828_adj_5495, 
        n60407, n256_adj_5496, n755_adj_5498, n60406, n682_adj_5502, 
        n60405, n329_adj_5504, n92_adj_5506, n23_adj_5507, n165_adj_5508;
    wire [18:0]n15206;
    
    wire n59528, n59527, n59526, n59525, n238_adj_5511, n59524, 
        n1105_adj_5512, n59523, n1032_adj_5513, n59522, n959_adj_5514, 
        n59521, n886_adj_5516, n59520, n813_adj_5517, n59519, n740_adj_5518, 
        n59518, n311_adj_5519, n667_adj_5521, n59517, n594_adj_5522, 
        n59516, n521_adj_5523, n59515, n448_adj_5524, n59514, n609_adj_5525, 
        n60404, n536_adj_5526, n60403, n375_adj_5527, n59513, n384_adj_5528, 
        n457_adj_5529, n302_adj_5530, n59512, n530_adj_5531, n229_adj_5532, 
        n59511, n156_adj_5533, n59510, n14_adj_5535, n83_adj_5536, 
        n463_adj_5537, n60402, n402_adj_5538, n603_adj_5539, n676_adj_5540, 
        n749_adj_5541, n822_adj_5542, n895_adj_5543, n968_adj_5544, 
        n390_adj_5545, n60401, n317_adj_5547, n60400, n1041_adj_5548, 
        n1114_adj_5550, n475_adj_5551, n244_adj_5552, n60399, n119, 
        n50, n171_adj_5554, n60398, n29_adj_5555, n98_adj_5556, n192, 
        n265, n338, n548_adj_5557;
    wire [23:0]n1_adj_5702;
    wire [6:0]n20178;
    
    wire n630, n60397, n557, n60396, n411, n484_adj_5559, n60395, 
        n484_adj_5560, n557_adj_5561, n630_adj_5562, n411_adj_5563, 
        n60394, n621_adj_5564, n338_adj_5567, n60393, n694_adj_5568, 
        n265_adj_5569, n60392, n192_adj_5571, n60391;
    wire [7:0]n20132;
    
    wire n700_adj_5572, n59489, n50_adj_5573, n119_adj_5574;
    wire [12:0]n18922;
    
    wire n1050_adj_5575, n60390, n627_adj_5576, n59488, n977_adj_5577, 
        n60389, n554_adj_5578, n59487, n481_adj_5579, n59486, n767_adj_5582, 
        n904_adj_5583, n60388, n408_adj_5584, n59485, n58937, n335_adj_5587, 
        n59484, n831_adj_5588, n60387, n758_adj_5590, n60386, n262_adj_5591, 
        n59483, n685_adj_5592, n60385, n840_adj_5593, n612_adj_5594, 
        n60384, n89_adj_5595, n189_adj_5596, n59482, n20_adj_5597, 
        n47_adj_5598, n116_adj_5599, n539_adj_5600, n60383, n466_adj_5601, 
        n60382, n393_adj_5602, n60381;
    wire [17:0]n15965;
    
    wire n59481, n59480, n107_adj_5603, n320_adj_5604, n60380, n247_adj_5605, 
        n60379, n174_adj_5606, n60378, n162_adj_5607, n32_adj_5608, 
        n101_adj_5609, n235_adj_5610;
    wire [11:0]n19256;
    
    wire n980_adj_5611, n60377, n308_adj_5612, n907_adj_5614, n60376, 
        n834_adj_5615, n60375, n381_adj_5616, n761_adj_5617, n60374, 
        n59479, n454_adj_5619, n688_adj_5620, n60373, n527_adj_5621, 
        n600_adj_5622, n59478, n673_adj_5623, n58936, n615_adj_5624, 
        n60372, n746_adj_5626, n542_adj_5627, n60371, n819_adj_5628, 
        n892_adj_5630, n1108_adj_5631, n59477, n965_adj_5632, n1035_adj_5633, 
        n59476, n469_adj_5634, n60370, n1038_adj_5635, n1111_adj_5637, 
        n396_adj_5638, n60369, n323_adj_5639, n60368, n250_adj_5640, 
        n60367, n58935, n180_adj_5642, n962_adj_5643, n59475, n889_adj_5644, 
        n59474, n177_adj_5645, n60366, n35_adj_5647, n104_adj_5648, 
        n75323;
    wire [5:0]n20289;
    
    wire n560_adj_5649, n60365, n816_adj_5650, n59473, n253_adj_5652, 
        n743_adj_5653, n59472, n487_adj_5654, n60364, n414_adj_5655, 
        n60363, n670_adj_5656, n59471, n341_adj_5657, n60362, n58910, 
        n326_adj_5660, n268_adj_5662, n60361, n195_adj_5665, n60360, 
        n399_adj_5667, n472_adj_5668, n58934, n597_adj_5669, n59470, 
        n545_adj_5670, n53_adj_5672, n122_adj_5673;
    wire [10:0]n19540;
    
    wire n910_adj_5674, n60359, n837_adj_5675, n60358, n618_adj_5677, 
        n764_adj_5678, n60357, n691_adj_5679, n524_adj_5680, n59469, 
        n451_adj_5681, n59468, n378_adj_5682, n59467, n305_adj_5683, 
        n59466, n232_adj_5684, n59465, n159_adj_5685, n59464, n86_adj_5686, 
        n17_adj_5687, n60356, n60355, n59122, n59121, n60354, n60353, 
        n60352, n59120, n59119, n59118, n59117, n58933, n60351, 
        n59116, n58932, n58909, n58908, n60350, n59115, n79534, 
        n59114, n58931, n60349;
    wire [16:0]n16648;
    
    wire n59444, n59443, n59442, n59113, n59441, n59112, n59440, 
        n59439, n59438, n59111, n59437, n59436, n59110, n59435, 
        n59434, n59433, n59432, n59109, n59431, n58930, n59108, 
        n59430, n59429, n59428, n58929, n60348, n59107, n59106, 
        n59105, n60347, n59104, n59103, n58928, n59102, n60346, 
        n59101, n59100, n60345;
    wire [6:0]n20256;
    
    wire n59409, n59408, n59407, n59406, n58927, n60344, n59405, 
        n59404, n59403, n58926;
    wire [15:0]n17259;
    
    wire n59402, n60343, n59401, n59400, n59099, n59399, n59098, 
        n59398, n59397, n59396, n59395, n59394, n59393, n60342, 
        n58925, n59097, n59392, n59391, n59390, n58924, n59096, 
        n59389, n59095, n59388, n59094, n59093, n59387, n59092, 
        n60341, n59091, n59090, n59089, n59088, n59087, n60340, 
        n60339;
    wire [14:0]n17802;
    
    wire n59369, n60338, n59368, n59367, n59366, n60337, n60336, 
        n60335, n59086, n60334, n59365, n58923, n58922, n59364, 
        n58921, n58920, n59363, n58919, n58918, n59362, n59085, 
        n59361, n59084, n59360, n59359, n59083, n59358, n59357, 
        n59356, n59355, n59082, n59081, n59080, n59079, n59078, 
        n58789, n59338, n59337, n59336, n59077, n59335, n59334, 
        n59333;
    wire [13:0]n18281;
    
    wire n59332, n59331, n59330, n59329, n59328, n58976, n59327, 
        n58975, n59326, n59325, n59324, n59323, n59322, n59321, 
        n59320, n58974, n59319, n58973, n58972, n58971, n58970, 
        n58969, n58968, n59076, n59075, n59303, n59074, n58967, 
        n59073, n59302, n59072, n58966, n59301, n59300, n59071, 
        n59299, n59070, n58965, n59298, n59069, n59297, n58964, 
        n59296, n59295, n59294, n58963, n59293, n59292, n59291, 
        n58962, n58961, n58960, n58959, n79276, n79498, n79492, 
        n79270, n79486, n79480, n79264, n79474, n79258, n79468, 
        n79462, n79246, n58814, n69713, n18_adj_5695, n20_adj_5696, 
        n7_adj_5697, n79222;
    
    SB_CARRY unary_minus_20_add_3_16 (.CI(n59067), .I0(GND_net), .I1(n1[14]), 
            .CO(n59068));
    SB_LUT4 LessThan_17_i24_3_lut (.I0(n16_c), .I1(n233[22]), .I2(n45), 
            .I3(GND_net), .O(n24_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60106_4_lut (.I0(n43), .I1(n25_c), .I2(n23), .I3(n76006), 
            .O(n75962));
    defparam i60106_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6622_6 (.CI(n59275), .I0(n20418[3]), .I1(n417), .CO(n59276));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n59066), .O(n285[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61697_4_lut (.I0(n24_c), .I1(n8_c), .I2(n45), .I3(n75960), 
            .O(n77553));   // verilog/motorControl.v(56[14:36])
    defparam i61697_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60607_3_lut (.I0(n77724), .I1(n233[12]), .I2(n25_c), .I3(GND_net), 
            .O(n76463));   // verilog/motorControl.v(56[14:36])
    defparam i60607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(n233[0]), .I1(n233[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 mult_23_i226_2_lut (.I0(\Kp[4] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6622_5_lut (.I0(GND_net), .I1(n20421), .I2(n344_c), .I3(n59274), 
            .O(n20350[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n59066), .I0(GND_net), .I1(n1[13]), 
            .CO(n59067));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n59065), .O(n285[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_6 (.CI(n58957), .I0(n360[4]), .I1(n46[4]), .CO(n58958));
    SB_LUT4 mult_23_i275_2_lut (.I0(\Kp[5] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59794_2_lut (.I0(PWMLimit[12]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75265));
    defparam i59794_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i21_3_lut (.I0(n233[20]), .I1(n285[20]), .I2(n284), 
            .I3(GND_net), .O(n310[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i124_2_lut (.I0(\Kp[2] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i173_2_lut (.I0(\Kp[3] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_5136));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i222_2_lut (.I0(\Kp[4] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i345_2_lut (.I0(\Kp[7] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i271_2_lut (.I0(\Kp[5] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i320_2_lut (.I0(\Kp[6] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i394_2_lut (.I0(\Kp[8] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i443_2_lut (.I0(\Kp[9] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i369_2_lut (.I0(\Kp[7] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i492_2_lut (.I0(\Kp[10] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i541_2_lut (.I0(\Kp[11] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59780_2_lut (.I0(PWMLimit[13]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75266));
    defparam i59780_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i418_2_lut (.I0(\Kp[8] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i590_2_lut (.I0(\Kp[12] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i467_2_lut (.I0(\Kp[9] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61865_3_lut (.I0(n4_c), .I1(n233[13]), .I2(n27), .I3(GND_net), 
            .O(n77721));   // verilog/motorControl.v(56[14:36])
    defparam i61865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i516_2_lut (.I0(\Kp[10] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i565_2_lut (.I0(\Kp[11] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i4_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n284), .I3(GND_net), 
            .O(n310[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i4_3_lut (.I0(n310[3]), .I1(IntegralLimit[3]), .I2(n258), 
            .I3(GND_net), .O(n356));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i55_2_lut (.I0(\Ki[1] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i8_2_lut (.I0(\Ki[0] ), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n11_adj_5137));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i21_3_lut (.I0(n310[20]), .I1(IntegralLimit[20]), .I2(n258), 
            .I3(GND_net), .O(n339));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61866_3_lut (.I0(n77721), .I1(n233[14]), .I2(n29), .I3(GND_net), 
            .O(n77722));   // verilog/motorControl.v(56[14:36])
    defparam i61866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i104_2_lut (.I0(\Ki[2] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i153_2_lut (.I0(\Ki[3] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60124_4_lut (.I0(n33_c), .I1(n31), .I2(n29), .I3(n75992), 
            .O(n75980));
    defparam i60124_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62209_4_lut (.I0(n30), .I1(n10_c), .I2(n35_c), .I3(n75976), 
            .O(n78065));   // verilog/motorControl.v(56[14:36])
    defparam i62209_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60609_3_lut (.I0(n77722), .I1(n233[15]), .I2(n31), .I3(GND_net), 
            .O(n76465));   // verilog/motorControl.v(56[14:36])
    defparam i60609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62363_4_lut (.I0(n76465), .I1(n78065), .I2(n35_c), .I3(n75980), 
            .O(n78219));   // verilog/motorControl.v(56[14:36])
    defparam i62363_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62364_3_lut (.I0(n78219), .I1(n239), .I2(n37_c), .I3(GND_net), 
            .O(n78220));   // verilog/motorControl.v(56[14:36])
    defparam i62364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62332_3_lut (.I0(n78220), .I1(n233[19]), .I2(n39), .I3(GND_net), 
            .O(n78188));   // verilog/motorControl.v(56[14:36])
    defparam i62332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60108_4_lut (.I0(n43), .I1(n41_c), .I2(n39), .I3(n78132), 
            .O(n75964));
    defparam i60108_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62186_4_lut (.I0(n76463), .I1(n77553), .I2(n45), .I3(n75962), 
            .O(n78042));   // verilog/motorControl.v(56[14:36])
    defparam i62186_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i639_2_lut (.I0(\Kp[13] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i688_2_lut (.I0(\Kp[14] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i202_2_lut (.I0(\Ki[4] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n299_c));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i251_2_lut (.I0(\Ki[5] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i737_2_lut (.I0(\Kp[15] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i300_2_lut (.I0(\Ki[6] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60615_3_lut (.I0(n78188), .I1(n233[20]), .I2(n41_c), .I3(GND_net), 
            .O(n76471));   // verilog/motorControl.v(56[14:36])
    defparam i60615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i126_2_lut (.I0(\Ki[2] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i349_2_lut (.I0(\Ki[7] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i398_2_lut (.I0(\Ki[8] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i447_2_lut (.I0(\Ki[9] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i496_2_lut (.I0(\Ki[10] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i545_2_lut (.I0(\Ki[11] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i594_2_lut (.I0(\Ki[12] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i643_2_lut (.I0(\Ki[13] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i692_2_lut (.I0(\Ki[14] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i741_2_lut (.I0(\Ki[15] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i175_2_lut (.I0(\Ki[3] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i3_3_lut (.I0(n233[2]), .I1(n285[2]), .I2(n284), .I3(GND_net), 
            .O(n310[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i3_3_lut (.I0(n310[2]), .I1(IntegralLimit[2]), .I2(n258), 
            .I3(GND_net), .O(n357));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i53_2_lut (.I0(\Ki[1] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i6_2_lut (.I0(\Ki[0] ), .I1(n357), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_5138));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i102_2_lut (.I0(\Ki[2] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i102_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n59065), .I0(GND_net), .I1(n1[12]), 
            .CO(n59066));
    SB_LUT4 mult_24_i151_2_lut (.I0(\Ki[3] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i224_2_lut (.I0(\Ki[4] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_5139));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i200_2_lut (.I0(\Ki[4] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_5140));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i249_2_lut (.I0(\Ki[5] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i298_2_lut (.I0(\Ki[6] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n59064), .O(n285[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n59064), .I0(GND_net), .I1(n1[11]), 
            .CO(n59065));
    SB_CARRY add_6622_5 (.CI(n59274), .I0(n20421), .I1(n344_c), .CO(n59275));
    SB_LUT4 add_6622_4_lut (.I0(GND_net), .I1(n20422), .I2(n271), .I3(n59273), 
            .O(n20350[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62188_4_lut (.I0(n76471), .I1(n78042), .I2(n45), .I3(n75964), 
            .O(n78044));   // verilog/motorControl.v(56[14:36])
    defparam i62188_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n59063), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6622_4 (.CI(n59273), .I0(n20422), .I1(n271), .CO(n59274));
    SB_LUT4 add_6622_3_lut (.I0(GND_net), .I1(n20418[0]), .I2(n198), .I3(n59272), 
            .O(n20350[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6622_3 (.CI(n59272), .I0(n20418[0]), .I1(n198), .CO(n59273));
    SB_LUT4 counter_2045_2046_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[13]), .I3(n60269), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i347_2_lut (.I0(\Ki[7] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[12]), .I3(n60268), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n79225), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFF control_update_46 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(24[10] 31[6])
    SB_LUT4 mult_24_i396_2_lut (.I0(\Ki[8] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i396_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2045_2046_add_4_14 (.CI(n60268), .I0(GND_net), .I1(counter[12]), 
            .CO(n60269));
    SB_LUT4 counter_2045_2046_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[11]), .I3(n60267), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6622_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20350[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6622_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n59272));
    SB_CARRY counter_2045_2046_add_4_13 (.CI(n60267), .I0(GND_net), .I1(counter[11]), 
            .CO(n60268));
    SB_CARRY unary_minus_20_add_3_12 (.CI(n59063), .I0(GND_net), .I1(n1[10]), 
            .CO(n59064));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n59062), .O(n285[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59620_2_lut (.I0(PWMLimit[11]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75264));
    defparam i59620_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(n360[3]), .I2(n46[3]), .I3(n58956), 
            .O(n455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i445_2_lut (.I0(\Ki[9] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[10]), .I3(n60266), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_12 (.CI(n60266), .I0(GND_net), .I1(counter[10]), 
            .CO(n60267));
    SB_LUT4 mult_24_i494_2_lut (.I0(\Ki[10] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[9]), .I3(n60265), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_14_lut (.I0(GND_net), .I1(n19063[11]), .I2(n980), 
            .I3(n59271), .O(n18700[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_13_lut (.I0(GND_net), .I1(n19063[10]), .I2(n907), 
            .I3(n59270), .O(n18700[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n58916), .O(n207[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_11 (.CI(n60265), .I0(GND_net), .I1(counter[9]), 
            .CO(n60266));
    SB_LUT4 counter_2045_2046_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[8]), .I3(n60264), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_10 (.CI(n60264), .I0(GND_net), .I1(counter[8]), 
            .CO(n60265));
    SB_LUT4 counter_2045_2046_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n60263), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n59062), .I0(GND_net), .I1(n1[9]), 
            .CO(n59063));
    SB_LUT4 i62189_3_lut (.I0(n78044), .I1(IntegralLimit[23]), .I2(n233[23]), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(56[14:36])
    defparam i62189_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY counter_2045_2046_add_4_9 (.CI(n60263), .I0(GND_net), .I1(counter[7]), 
            .CO(n60264));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n59061), .O(n285[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_13 (.CI(n59270), .I0(n19063[10]), .I1(n907), .CO(n59271));
    SB_LUT4 mult_24_i543_2_lut (.I0(\Ki[11] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n60262), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i592_2_lut (.I0(\Ki[12] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i20_3_lut (.I0(n233[19]), .I1(n285[19]), .I2(n284), 
            .I3(GND_net), .O(n310[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i20_3_lut (.I0(n310[19]), .I1(IntegralLimit[19]), .I2(n258), 
            .I3(GND_net), .O(n340));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_2045_2046_add_4_8 (.CI(n60262), .I0(GND_net), .I1(counter[6]), 
            .CO(n60263));
    SB_LUT4 counter_2045_2046_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n60261), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_7 (.CI(n60261), .I0(GND_net), .I1(counter[5]), 
            .CO(n60262));
    SB_LUT4 counter_2045_2046_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n60260), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i641_2_lut (.I0(\Ki[13] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i641_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2045_2046_add_4_6 (.CI(n60260), .I0(GND_net), .I1(counter[4]), 
            .CO(n60261));
    SB_LUT4 counter_2045_2046_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n60259), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i690_2_lut (.I0(\Ki[14] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i690_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2045_2046_add_4_5 (.CI(n60259), .I0(GND_net), .I1(counter[3]), 
            .CO(n60260));
    SB_LUT4 add_6481_12_lut (.I0(GND_net), .I1(n19063[9]), .I2(n834), 
            .I3(n59269), .O(n18700[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_12 (.CI(n59269), .I0(n19063[9]), .I1(n834), .CO(n59270));
    SB_LUT4 counter_2045_2046_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n60258), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i739_2_lut (.I0(\Ki[15] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i739_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2045_2046_add_4_4 (.CI(n60258), .I0(GND_net), .I1(counter[2]), 
            .CO(n60259));
    SB_LUT4 LessThan_17_i37_2_lut (.I0(IntegralLimit[18]), .I1(n239), .I2(GND_net), 
            .I3(GND_net), .O(n37_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6481_11_lut (.I0(GND_net), .I1(n19063[8]), .I2(n761), 
            .I3(n59268), .O(n18700[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n59061), .I0(GND_net), .I1(n1[8]), 
            .CO(n59062));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n59060), .O(n285[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n59060), .I0(GND_net), .I1(n1[7]), 
            .CO(n59061));
    SB_LUT4 counter_2045_2046_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n60257), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_3 (.CI(n60257), .I0(GND_net), .I1(counter[1]), 
            .CO(n60258));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n59059), .O(n285[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_5 (.CI(n58956), .I0(n360[3]), .I1(n46[3]), .CO(n58957));
    SB_LUT4 counter_2045_2046_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(n360[2]), .I2(n46[2]), .I3(n58955), 
            .O(n455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n60257));
    SB_CARRY add_6481_11 (.CI(n59268), .I0(n19063[8]), .I1(n761), .CO(n59269));
    SB_CARRY unary_minus_20_add_3_8 (.CI(n59059), .I0(GND_net), .I1(n1[6]), 
            .CO(n59060));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n59058), .O(n285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_10_lut (.I0(GND_net), .I1(n19063[7]), .I2(n688), 
            .I3(n59267), .O(n18700[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_10 (.CI(n59267), .I0(n19063[7]), .I1(n688), .CO(n59268));
    SB_LUT4 add_6481_9_lut (.I0(GND_net), .I1(n19063[6]), .I2(n615), .I3(n59266), 
            .O(n18700[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_9 (.CI(n59266), .I0(n19063[6]), .I1(n615), .CO(n59267));
    SB_LUT4 add_6481_8_lut (.I0(GND_net), .I1(n19063[5]), .I2(n542), .I3(n59265), 
            .O(n18700[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n59058), .I0(GND_net), .I1(n1[5]), 
            .CO(n59059));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n59057), .O(n285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_8 (.CI(n59265), .I0(n19063[5]), .I1(n542), .CO(n59266));
    SB_LUT4 add_6481_7_lut (.I0(GND_net), .I1(n19063[4]), .I2(n469), .I3(n59264), 
            .O(n18700[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n59057), .I0(GND_net), .I1(n1[4]), 
            .CO(n59058));
    SB_CARRY add_6481_7 (.CI(n59264), .I0(n19063[4]), .I1(n469), .CO(n59265));
    SB_CARRY add_25_4 (.CI(n58955), .I0(n360[2]), .I1(n46[2]), .CO(n58956));
    SB_LUT4 add_6481_6_lut (.I0(GND_net), .I1(n19063[3]), .I2(n396), .I3(n59263), 
            .O(n18700[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n59056), .O(n285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_6 (.CI(n59263), .I0(n19063[3]), .I1(n396), .CO(n59264));
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(n360[1]), .I2(n46[1]), .I3(n58954), 
            .O(n455[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_11 (.CI(n58916), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n58917));
    SB_CARRY unary_minus_20_add_3_5 (.CI(n59056), .I0(GND_net), .I1(n1[3]), 
            .CO(n59057));
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n59055), .O(n285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_3 (.CI(n58954), .I0(n360[1]), .I1(n46[1]), .CO(n58955));
    SB_LUT4 i59765_2_lut (.I0(PWMLimit[14]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75274));
    defparam i59765_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n58915), .O(n207[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_5_lut (.I0(GND_net), .I1(n19063[2]), .I2(n323), .I3(n59262), 
            .O(n18700[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n59055), .I0(GND_net), .I1(n1[2]), 
            .CO(n59056));
    SB_CARRY add_6481_5 (.CI(n59262), .I0(n19063[2]), .I1(n323), .CO(n59263));
    SB_LUT4 add_6481_4_lut (.I0(GND_net), .I1(n19063[1]), .I2(n250), .I3(n59261), 
            .O(n18700[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(n360[0]), .I2(n46[0]), .I3(GND_net), 
            .O(n455[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_4 (.CI(n59261), .I0(n19063[1]), .I1(n250), .CO(n59262));
    SB_LUT4 add_6481_3_lut (.I0(GND_net), .I1(n19063[0]), .I2(n177), .I3(n59260), 
            .O(n18700[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_21_i2_3_lut (.I0(n233[1]), .I1(n285[1]), .I2(n284), .I3(GND_net), 
            .O(n310[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i2_3_lut (.I0(n310[1]), .I1(IntegralLimit[1]), .I2(n258), 
            .I3(GND_net), .O(n358));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i51_2_lut (.I0(\Ki[1] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_5146));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i4_2_lut (.I0(\Ki[0] ), .I1(n358), .I2(GND_net), .I3(GND_net), 
            .O(n5));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i100_2_lut (.I0(\Ki[2] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i45_2_lut (.I0(IntegralLimit[22]), .I1(n233[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i149_2_lut (.I0(\Ki[3] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6481_3 (.CI(n59260), .I0(n19063[0]), .I1(n177), .CO(n59261));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n59054), .O(n285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_2_lut (.I0(GND_net), .I1(n35_adj_5148), .I2(n104), 
            .I3(GND_net), .O(n18700[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_2 (.CI(GND_net), .I0(n360[0]), .I1(n46[0]), .CO(n58954));
    SB_LUT4 LessThan_17_i41_2_lut (.I0(IntegralLimit[20]), .I1(n233[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_15_add_2_10 (.CI(n58915), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n58916));
    SB_LUT4 mult_24_i198_2_lut (.I0(\Ki[4] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i198_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6481_2 (.CI(GND_net), .I0(n35_adj_5148), .I1(n104), .CO(n59260));
    SB_LUT4 mult_24_i247_2_lut (.I0(\Ki[5] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i43_2_lut (.I0(IntegralLimit[21]), .I1(n233[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i296_2_lut (.I0(\Ki[6] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n58914), .O(n207[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n59054), .I0(GND_net), .I1(n1[1]), 
            .CO(n59055));
    SB_LUT4 LessThan_17_i35_2_lut (.I0(IntegralLimit[17]), .I1(n233[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i31_2_lut (.I0(IntegralLimit[15]), .I1(n233[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i345_2_lut (.I0(\Ki[7] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_5149));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n207[23]), .I3(n58953), .O(n233[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i394_2_lut (.I0(\Ki[8] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_5151));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n59054));
    SB_LUT4 add_16_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n207[23]), .I3(n58952), .O(n233[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_24 (.CI(n58952), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n207[23]), .CO(n58953));
    SB_LUT4 mult_24_i443_2_lut (.I0(\Ki[9] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_5152));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i492_2_lut (.I0(\Ki[10] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_5153));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i541_2_lut (.I0(\Ki[11] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_5154));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i590_2_lut (.I0(\Ki[12] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_5155));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i639_2_lut (.I0(\Ki[13] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_5156));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i33_2_lut (.I0(IntegralLimit[16]), .I1(n233[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i688_2_lut (.I0(\Ki[14] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_5157));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i737_2_lut (.I0(\Ki[15] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_5158));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i324_2_lut (.I0(\Kp[6] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i39_2_lut (.I0(IntegralLimit[19]), .I1(n233[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_16_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n207[23]), .I3(n58951), .O(n233[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11882_bdd_4_lut_63541 (.I0(n11882), .I1(n75285), .I2(setpoint[15]), 
            .I3(n4736), .O(n79384));
    defparam n11882_bdd_4_lut_63541.LUT_INIT = 16'he4aa;
    SB_CARRY add_16_23 (.CI(n58951), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n207[23]), .CO(n58952));
    SB_LUT4 mux_21_i24_3_lut (.I0(n233[23]), .I1(n285[23]), .I2(n284), 
            .I3(GND_net), .O(n310[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i24_3_lut (.I0(n310[23]), .I1(IntegralLimit[23]), .I2(n258), 
            .I3(GND_net), .O(n336));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i29_2_lut (.I0(IntegralLimit[14]), .I1(n233[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60150_4_lut (.I0(n21_adj_5159), .I1(n19_adj_5160), .I2(n17_adj_5161), 
            .I3(n9_c), .O(n76006));
    defparam i60150_4_lut.LUT_INIT = 16'haaab;
    SB_DFFER result_i0_i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n79537), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i60136_4_lut (.I0(n27), .I1(n15_adj_5162), .I2(n13_adj_5163), 
            .I3(n11_adj_5164), .O(n75992));
    defparam i60136_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n233[7]), .I1(n233[16]), .I2(n33_c), 
            .I3(GND_net), .O(n12_adj_5166));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n79501), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n79495), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n79489), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_16_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n207[23]), .I3(n58950), .O(n233[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_22_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n79483), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 n79384_bdd_4_lut (.I0(n79384), .I1(n535[15]), .I2(n455[15]), 
            .I3(n4736), .O(n79387));
    defparam n79384_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_16_22 (.CI(n58950), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n207[23]), .CO(n58951));
    SB_DFFER result_i0_i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n79477), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n233[5]), .I1(n233[6]), .I2(n13_adj_5163), 
            .I3(GND_net), .O(n10_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i30_3_lut (.I0(n12_adj_5166), .I1(n233[17]), .I2(n35_c), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n79471), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n79465), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_16_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n207[23]), .I3(n58949), .O(n233[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_21 (.CI(n58949), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n207[23]), .CO(n58950));
    SB_LUT4 add_16_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n207[22]), .I3(n58948), .O(n239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_9 (.CI(n58914), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n58915));
    SB_CARRY add_16_20 (.CI(n58948), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n207[22]), .CO(n58949));
    SB_LUT4 add_16_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n207[21]), .I3(n58947), .O(n233[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n58913), .O(n207[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_19 (.CI(n58947), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n207[21]), .CO(n58948));
    SB_LUT4 LessThan_19_i45_2_lut (.I0(n233[22]), .I1(n285[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5167));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(n233[19]), .I1(n285[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5168));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(n233[20]), .I1(n285[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5169));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_16_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n207[20]), .I3(n58946), .O(n233[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_8 (.CI(n58913), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n58914));
    SB_LUT4 sub_15_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n58912), .O(n207[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_18 (.CI(n58946), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n207[20]), .CO(n58947));
    SB_LUT4 add_16_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n207[19]), .I3(n58945), .O(n233[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_17 (.CI(n58945), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n207[19]), .CO(n58946));
    SB_LUT4 i61099_4_lut (.I0(n13_adj_5163), .I1(n11_adj_5164), .I2(n9_c), 
            .I3(n76024), .O(n76955));
    defparam i61099_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(n233[21]), .I1(n285[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5171));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(n233[16]), .I1(n285[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5173));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(n233[17]), .I1(n285[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5174));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i373_2_lut (.I0(\Kp[7] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n207[18]), .I3(n58944), .O(n233[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(n233[13]), .I1(n285[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5175));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i61093_4_lut (.I0(n19_adj_5160), .I1(n17_adj_5161), .I2(n15_adj_5162), 
            .I3(n76955), .O(n76949));
    defparam i61093_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(n233[14]), .I1(n285[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5176));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_15_add_2_7 (.CI(n58912), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n58913));
    SB_CARRY add_16_16 (.CI(n58944), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n207[18]), .CO(n58945));
    SB_LUT4 LessThan_19_i31_2_lut (.I0(n233[15]), .I1(n285[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5177));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60088_4_lut (.I0(n21), .I1(n19_adj_5179), .I2(n17_adj_5180), 
            .I3(n9_adj_5181), .O(n75944));
    defparam i60088_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i273_2_lut (.I0(\Ki[5] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n207[17]), .I3(n58943), .O(n233[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60078_4_lut (.I0(n27_adj_5175), .I1(n15_adj_5182), .I2(n13_adj_5183), 
            .I3(n11_adj_5184), .O(n75934));
    defparam i60078_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62138_4_lut (.I0(n25_c), .I1(n23), .I2(n21_adj_5159), .I3(n76949), 
            .O(n77994));
    defparam i62138_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_32_i41_2_lut (.I0(n455[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5185));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i39_2_lut (.I0(n460), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5186));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i45_2_lut (.I0(n455[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5187));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i61551_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n77994), 
            .O(n77407));
    defparam i61551_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n285[7]), .I1(n285[16]), .I2(n33_adj_5173), 
            .I3(GND_net), .O(n12_adj_5188));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i29_2_lut (.I0(n455[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5189));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i31_2_lut (.I0(n455[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5190));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i43_2_lut (.I0(n455[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5191));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i37_2_lut (.I0(n461), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5192));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n285[5]), .I1(n285[6]), .I2(n13_adj_5183), 
            .I3(GND_net), .O(n10_adj_5193));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62276_4_lut (.I0(n37_c), .I1(n35_c), .I2(n33_c), .I3(n77407), 
            .O(n78132));
    defparam i62276_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_5188), .I1(n285[17]), .I2(n35_adj_5174), 
            .I3(GND_net), .O(n30_adj_5194));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i17_2_lut (.I0(n455[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5195));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i19_2_lut (.I0(n455[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5196));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i21_2_lut (.I0(n455[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5198));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i23_2_lut (.I0(n455[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5200));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i25_2_lut (.I0(n467), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5201));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i61039_4_lut (.I0(n13_adj_5183), .I1(n11_adj_5184), .I2(n9_adj_5181), 
            .I3(n75956), .O(n76895));
    defparam i61039_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n233[9]), .I1(n233[21]), .I2(n43), 
            .I3(GND_net), .O(n16_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61033_4_lut (.I0(n19_adj_5179), .I1(n17_adj_5180), .I2(n15_adj_5182), 
            .I3(n76895), .O(n76889));
    defparam i61033_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_32_i9_2_lut (.I0(n475), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5203));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62124_4_lut (.I0(n25_adj_5204), .I1(n23_adj_5205), .I2(n21), 
            .I3(n76889), .O(n77980));
    defparam i62124_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_32_i35_2_lut (.I0(n462), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5207));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(setpoint[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5208));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(setpoint[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5209));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i45_2_lut (.I0(setpoint[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5210));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5211));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(setpoint[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5212));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i31_2_lut (.I0(setpoint[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5213));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i61867_3_lut (.I0(n6_c), .I1(n247), .I2(n21_adj_5159), .I3(GND_net), 
            .O(n77723));   // verilog/motorControl.v(56[14:36])
    defparam i61867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(setpoint[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5214));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(setpoint[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5215));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n11882_bdd_4_lut_63476 (.I0(n11882), .I1(n75274), .I2(setpoint[14]), 
            .I3(n4736), .O(n79348));
    defparam n11882_bdd_4_lut_63476.LUT_INIT = 16'he4aa;
    SB_LUT4 n79348_bdd_4_lut (.I0(n79348), .I1(n535[14]), .I2(n455[14]), 
            .I3(n4736), .O(n79351));
    defparam n79348_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFER result_i0_i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n79387), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_11_i25_2_lut (.I0(setpoint[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5216));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i61868_3_lut (.I0(n77723), .I1(n233[11]), .I2(n23), .I3(GND_net), 
            .O(n77724));   // verilog/motorControl.v(56[14:36])
    defparam i61868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(setpoint[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5217));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(setpoint[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5218));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(setpoint[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5219));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(setpoint[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5220));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(setpoint[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5221));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5222));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i43_2_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5223));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i61523_4_lut (.I0(n31_adj_5177), .I1(n29_adj_5176), .I2(n27_adj_5175), 
            .I3(n77980), .O(n77379));
    defparam i61523_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n233[4]), .I1(n233[8]), .I2(n17_adj_5161), 
            .I3(GND_net), .O(n8_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i39_2_lut (.I0(PWMLimit[19]), .I1(setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5224));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62272_4_lut (.I0(n37), .I1(n35_adj_5174), .I2(n33_adj_5173), 
            .I3(n77379), .O(n78128));
    defparam i62272_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_9_i4_4_lut (.I0(PWMLimit[0]), .I1(setpoint[1]), .I2(PWMLimit[1]), 
            .I3(setpoint[0]), .O(n4_adj_5226));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_9_i8_3_lut (.I0(n6_adj_5227), .I1(setpoint[4]), .I2(n9), 
            .I3(GND_net), .O(n8_adj_5229));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62203_4_lut (.I0(n8_adj_5229), .I1(n4_adj_5226), .I2(n9), 
            .I3(n76188), .O(n78059));   // verilog/motorControl.v(45[16:33])
    defparam i62203_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62204_3_lut (.I0(n78059), .I1(setpoint[5]), .I2(PWMLimit[5]), 
            .I3(GND_net), .O(n78060));   // verilog/motorControl.v(45[16:33])
    defparam i62204_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n285[9]), .I1(n285[21]), .I2(n43_adj_5171), 
            .I3(GND_net), .O(n16_adj_5230));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62095_3_lut (.I0(n78060), .I1(setpoint[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n77951));   // verilog/motorControl.v(45[16:33])
    defparam i62095_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60591_3_lut (.I0(n77951), .I1(setpoint[7]), .I2(PWMLimit[7]), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(45[16:33])
    defparam i60591_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFER result_i0_i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n79351), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 n11882_bdd_4_lut_63447 (.I0(n11882), .I1(n75266), .I2(setpoint[13]), 
            .I3(n4736), .O(n79324));
    defparam n11882_bdd_4_lut_63447.LUT_INIT = 16'he4aa;
    SB_DFFER result_i0_i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n79327), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n79321), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n79315), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_9_i20_3_lut (.I0(n34689), .I1(setpoint[9]), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_16_15 (.CI(n58943), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n207[17]), .CO(n58944));
    SB_LUT4 add_16_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n207[16]), .I3(n58942), .O(n233[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i422_2_lut (.I0(\Kp[8] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59797_2_lut (.I0(PWMLimit[6]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75259));
    defparam i59797_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i31_2_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5233));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i471_2_lut (.I0(\Kp[9] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i322_2_lut (.I0(\Ki[6] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_5234));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61861_3_lut (.I0(n6_adj_5235), .I1(n299), .I2(n21), .I3(GND_net), 
            .O(n77717));   // verilog/motorControl.v(58[23:46])
    defparam i61861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61862_3_lut (.I0(n77717), .I1(n285[11]), .I2(n23_adj_5205), 
            .I3(GND_net), .O(n77718));   // verilog/motorControl.v(58[23:46])
    defparam i61862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n285[4]), .I1(n285[8]), .I2(n17_adj_5180), 
            .I3(GND_net), .O(n8_adj_5236));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_5230), .I1(n285[22]), .I2(n45_adj_5167), 
            .I3(GND_net), .O(n24_adj_5237));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60044_4_lut (.I0(n43_adj_5171), .I1(n25_adj_5204), .I2(n23_adj_5205), 
            .I3(n75944), .O(n75900));
    defparam i60044_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61699_4_lut (.I0(n24_adj_5237), .I1(n8_adj_5236), .I2(n45_adj_5167), 
            .I3(n75894), .O(n77555));   // verilog/motorControl.v(58[23:46])
    defparam i61699_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60617_3_lut (.I0(n77718), .I1(n285[12]), .I2(n25_adj_5204), 
            .I3(GND_net), .O(n76473));   // verilog/motorControl.v(58[23:46])
    defparam i60617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(n233[0]), .I1(n285[1]), .I2(n233[1]), 
            .I3(n285[0]), .O(n4_adj_5238));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61859_3_lut (.I0(n4_adj_5238), .I1(n285[13]), .I2(n27_adj_5175), 
            .I3(GND_net), .O(n77715));   // verilog/motorControl.v(58[23:46])
    defparam i61859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61860_3_lut (.I0(n77715), .I1(n285[14]), .I2(n29_adj_5176), 
            .I3(GND_net), .O(n77716));   // verilog/motorControl.v(58[23:46])
    defparam i61860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60067_4_lut (.I0(n33_adj_5173), .I1(n31_adj_5177), .I2(n29_adj_5176), 
            .I3(n75934), .O(n75923));
    defparam i60067_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62211_4_lut (.I0(n30_adj_5194), .I1(n10_adj_5193), .I2(n35_adj_5174), 
            .I3(n75919), .O(n78067));   // verilog/motorControl.v(58[23:46])
    defparam i62211_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60619_3_lut (.I0(n77716), .I1(n285[15]), .I2(n31_adj_5177), 
            .I3(GND_net), .O(n76475));   // verilog/motorControl.v(58[23:46])
    defparam i60619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62365_4_lut (.I0(n76475), .I1(n78067), .I2(n35_adj_5174), 
            .I3(n75923), .O(n78221));   // verilog/motorControl.v(58[23:46])
    defparam i62365_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62366_3_lut (.I0(n78221), .I1(n291), .I2(n37), .I3(GND_net), 
            .O(n78222));   // verilog/motorControl.v(58[23:46])
    defparam i62366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62330_3_lut (.I0(n78222), .I1(n285[19]), .I2(n39_adj_5168), 
            .I3(GND_net), .O(n78186));   // verilog/motorControl.v(58[23:46])
    defparam i62330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60048_4_lut (.I0(n43_adj_5171), .I1(n41_adj_5169), .I2(n39_adj_5168), 
            .I3(n78128), .O(n75904));
    defparam i60048_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_9_i27_2_lut (.I0(PWMLimit[13]), .I1(setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5239));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i29_2_lut (.I0(PWMLimit[14]), .I1(setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5240));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i23_2_lut (.I0(PWMLimit[11]), .I1(setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5241));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60313_4_lut (.I0(n29_adj_5240), .I1(n27_adj_5239), .I2(n25), 
            .I3(n23_adj_5241), .O(n76169));
    defparam i60313_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60302_4_lut (.I0(n35), .I1(n33), .I2(n31_adj_5233), .I3(n76169), 
            .O(n76158));
    defparam i60302_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i371_2_lut (.I0(\Ki[7] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_5245));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i30_3_lut (.I0(n28), .I1(setpoint[16]), .I2(n33), 
            .I3(GND_net), .O(n30_adj_5246));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i34_3_lut (.I0(n26), .I1(setpoint[18]), .I2(n37_adj_27), 
            .I3(GND_net), .O(n34_c));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62205_4_lut (.I0(n34_c), .I1(n24_adj_5248), .I2(n37_adj_27), 
            .I3(n76154), .O(n78061));   // verilog/motorControl.v(45[16:33])
    defparam i62205_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62206_3_lut (.I0(n78061), .I1(setpoint[19]), .I2(n39_adj_5224), 
            .I3(GND_net), .O(n78062));   // verilog/motorControl.v(45[16:33])
    defparam i62206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62091_3_lut (.I0(n78062), .I1(setpoint[20]), .I2(n41), .I3(GND_net), 
            .O(n77947));   // verilog/motorControl.v(45[16:33])
    defparam i62091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61945_4_lut (.I0(n41), .I1(n39_adj_5224), .I2(n37_adj_27), 
            .I3(n76158), .O(n77801));
    defparam i61945_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62122_4_lut (.I0(n30_adj_5246), .I1(n22), .I2(n33), .I3(n76162), 
            .O(n77978));   // verilog/motorControl.v(45[16:33])
    defparam i62122_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 n79324_bdd_4_lut (.I0(n79324), .I1(n535[13]), .I2(n455[13]), 
            .I3(n4736), .O(n79327));
    defparam n79324_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i60595_3_lut (.I0(n77947), .I1(setpoint[21]), .I2(n43_adj_5223), 
            .I3(GND_net), .O(n76451));   // verilog/motorControl.v(45[16:33])
    defparam i60595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62268_4_lut (.I0(n76451), .I1(n77978), .I2(n43_adj_5223), 
            .I3(n77801), .O(n78124));   // verilog/motorControl.v(45[16:33])
    defparam i62268_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62269_3_lut (.I0(n78124), .I1(setpoint[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n78125));   // verilog/motorControl.v(45[16:33])
    defparam i62269_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61986_3_lut (.I0(n78125), .I1(PWMLimit[23]), .I2(setpoint[23]), 
            .I3(GND_net), .O(n105));   // verilog/motorControl.v(45[16:33])
    defparam i61986_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(setpoint[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5252));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(setpoint[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5253));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(setpoint[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5254));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(setpoint[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5255));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i37_2_lut (.I0(PWMLimit[18]), .I1(n461), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5256));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i15_2_lut (.I0(PWMLimit[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5257));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i13_2_lut (.I0(PWMLimit[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5258));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i19_2_lut (.I0(PWMLimit[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5259));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i17_2_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5260));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i7_2_lut (.I0(PWMLimit[3]), .I1(n455[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i11_2_lut (.I0(PWMLimit[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5261));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i5_2_lut (.I0(PWMLimit[2]), .I1(n455[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5262));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59860_4_lut (.I0(n11_adj_5261), .I1(n35782), .I2(n7), .I3(n5_adj_5262), 
            .O(n75716));
    defparam i59860_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_30_i8_3_lut (.I0(n475), .I1(n455[8]), .I2(n17_adj_5260), 
            .I3(GND_net), .O(n8_adj_5263));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i6_3_lut (.I0(n455[2]), .I1(n455[3]), .I2(n7), 
            .I3(GND_net), .O(n6_adj_5264));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i16_3_lut (.I0(n8_adj_5263), .I1(n455[9]), .I2(n19_adj_5259), 
            .I3(GND_net), .O(n16_adj_5265));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i4_4_lut (.I0(n455[0]), .I1(n455[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_5266));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i61431_3_lut (.I0(n4_adj_5266), .I1(n455[5]), .I2(n11_adj_5261), 
            .I3(GND_net), .O(n77287));   // verilog/motorControl.v(63[16:31])
    defparam i61431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61432_3_lut (.I0(n77287), .I1(n455[6]), .I2(n13_adj_5258), 
            .I3(GND_net), .O(n77288));   // verilog/motorControl.v(63[16:31])
    defparam i61432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59854_4_lut (.I0(n17_adj_5260), .I1(n15_adj_5257), .I2(n13_adj_5258), 
            .I3(n75716), .O(n75710));
    defparam i59854_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62018_4_lut (.I0(n16_adj_5265), .I1(n6_adj_5264), .I2(n19_adj_5259), 
            .I3(n75702), .O(n77874));   // verilog/motorControl.v(63[16:31])
    defparam i62018_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60641_3_lut (.I0(n77288), .I1(n455[7]), .I2(n15_adj_5257), 
            .I3(GND_net), .O(n76497));   // verilog/motorControl.v(63[16:31])
    defparam i60641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62379_4_lut (.I0(n76497), .I1(n77874), .I2(n19_adj_5259), 
            .I3(n75710), .O(n78235));   // verilog/motorControl.v(63[16:31])
    defparam i62379_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62380_3_lut (.I0(n78235), .I1(n455[10]), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n78236));   // verilog/motorControl.v(63[16:31])
    defparam i62380_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62302_3_lut (.I0(n78236), .I1(n455[11]), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(63[16:31])
    defparam i62302_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_30_i41_2_lut (.I0(PWMLimit[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5268));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i29_2_lut (.I0(PWMLimit[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5269));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i31_2_lut (.I0(PWMLimit[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5270));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i33_2_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5271));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i39_2_lut (.I0(PWMLimit[19]), .I1(n460), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5272));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i27_2_lut (.I0(PWMLimit[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5273));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59830_4_lut (.I0(n33_adj_5271), .I1(n31_adj_5270), .I2(n29_adj_5269), 
            .I3(n27_adj_5273), .O(n75686));
    defparam i59830_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_30_i30_3_lut (.I0(n455[15]), .I1(n460), .I2(n39_adj_5272), 
            .I3(GND_net), .O(n30_adj_5274));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i28_3_lut (.I0(n455[13]), .I1(n455[14]), .I2(n29_adj_5269), 
            .I3(GND_net), .O(n28_adj_5275));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i38_3_lut (.I0(n30_adj_5274), .I1(n455[20]), .I2(n41_adj_5268), 
            .I3(GND_net), .O(n38_c));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n79309), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i61429_3_lut (.I0(n36147), .I1(n455[16]), .I2(n33_adj_5271), 
            .I3(GND_net), .O(n77285));   // verilog/motorControl.v(63[16:31])
    defparam i61429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61430_3_lut (.I0(n77285), .I1(n462), .I2(n36361), .I3(GND_net), 
            .O(n77286));   // verilog/motorControl.v(63[16:31])
    defparam i61430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_15_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n58911), .O(n207[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59821_4_lut (.I0(n39_adj_5272), .I1(n37_adj_5256), .I2(n36361), 
            .I3(n75686), .O(n75677));
    defparam i59821_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62074_4_lut (.I0(n38_c), .I1(n28_adj_5275), .I2(n41_adj_5268), 
            .I3(n75675), .O(n77930));   // verilog/motorControl.v(63[16:31])
    defparam i62074_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60643_3_lut (.I0(n77286), .I1(n461), .I2(n37_adj_5256), .I3(GND_net), 
            .O(n76499));   // verilog/motorControl.v(63[16:31])
    defparam i60643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62327_4_lut (.I0(n76499), .I1(n77930), .I2(n41_adj_5268), 
            .I3(n75677), .O(n78183));   // verilog/motorControl.v(63[16:31])
    defparam i62327_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62328_3_lut (.I0(n78183), .I1(n455[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n78184));   // verilog/motorControl.v(63[16:31])
    defparam i62328_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62263_3_lut (.I0(n78184), .I1(n455[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n78119));   // verilog/motorControl.v(63[16:31])
    defparam i62263_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60649_3_lut (.I0(n78119), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(GND_net), .O(n508));   // verilog/motorControl.v(63[16:31])
    defparam i60649_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut (.I0(n44726), .I1(n25921), .I2(GND_net), .I3(GND_net), 
            .O(n25756));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 n11882_bdd_4_lut_63428 (.I0(n11882), .I1(n75265), .I2(setpoint[12]), 
            .I3(n4736), .O(n79318));
    defparam n11882_bdd_4_lut_63428.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_4_lut (.I0(control_update), .I1(n25756), .I2(n4), .I3(n508), 
            .O(n5076));
    defparam i2_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 i62190_4_lut (.I0(n76473), .I1(n77555), .I2(n45_adj_5167), 
            .I3(n75900), .O(n78046));   // verilog/motorControl.v(58[23:46])
    defparam i62190_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60228_4_lut (.I0(n21_adj_5221), .I1(n19_adj_5220), .I2(n17_adj_5219), 
            .I3(n9_adj_5218), .O(n76084));
    defparam i60228_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60202_4_lut (.I0(n27_adj_5255), .I1(n15_adj_5254), .I2(n13_adj_5253), 
            .I3(n11_adj_5252), .O(n76058));
    defparam i60202_4_lut.LUT_INIT = 16'haaab;
    SB_DFFER result_i0_i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n79303), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_5222), 
            .I3(GND_net), .O(n12_adj_5277));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n79297), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 n79318_bdd_4_lut (.I0(n79318), .I1(n535[12]), .I2(n467), .I3(n4736), 
            .O(n79321));
    defparam n79318_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_5253), 
            .I3(GND_net), .O(n10_adj_5278));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_5277), .I1(n535[17]), .I2(n35_adj_5217), 
            .I3(GND_net), .O(n30_adj_5279));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n79291), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i61167_4_lut (.I0(n13_adj_5253), .I1(n11_adj_5252), .I2(n9_adj_5218), 
            .I3(n76116), .O(n77023));
    defparam i61167_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61157_4_lut (.I0(n19_adj_5220), .I1(n17_adj_5219), .I2(n15_adj_5254), 
            .I3(n77023), .O(n77013));
    defparam i61157_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60625_3_lut (.I0(n78186), .I1(n285[20]), .I2(n41_adj_5169), 
            .I3(GND_net), .O(n76481));   // verilog/motorControl.v(58[23:46])
    defparam i60625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62150_4_lut (.I0(n25_adj_5216), .I1(n23_adj_5215), .I2(n21_adj_5221), 
            .I3(n77013), .O(n78006));
    defparam i62150_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61583_4_lut (.I0(n31_adj_5213), .I1(n29_adj_5212), .I2(n27_adj_5255), 
            .I3(n78006), .O(n77439));
    defparam i61583_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i62280_4_lut (.I0(n37_adj_5214), .I1(n35_adj_5217), .I2(n33_adj_5222), 
            .I3(n77439), .O(n78136));
    defparam i62280_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_5211), 
            .I3(GND_net), .O(n16_adj_5280));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n79285), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i61875_3_lut (.I0(n6_adj_5281), .I1(n535[10]), .I2(n21_adj_5221), 
            .I3(GND_net), .O(n77731));   // verilog/motorControl.v(47[25:43])
    defparam i61875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(IntegralLimit[4]), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(IntegralLimit[5]), .I1(n233[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5164));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(IntegralLimit[6]), .I1(n233[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5163));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i61876_3_lut (.I0(n77731), .I1(n535[11]), .I2(n23_adj_5215), 
            .I3(GND_net), .O(n77732));   // verilog/motorControl.v(47[25:43])
    defparam i61876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(IntegralLimit[7]), .I1(n233[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5162));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_DFFER result_i0_i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n79279), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_17_i21_2_lut (.I0(IntegralLimit[10]), .I1(n247), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5159));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_DFFER result_i0_i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n79273), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i62192_4_lut (.I0(n76481), .I1(n78046), .I2(n45_adj_5167), 
            .I3(n75904), .O(n78048));   // verilog/motorControl.v(58[23:46])
    defparam i62192_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(IntegralLimit[9]), .I1(n233[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5160));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(IntegralLimit[8]), .I1(n233[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5161));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(IntegralLimit[11]), .I1(n233[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i25_2_lut (.I0(IntegralLimit[12]), .I1(n233[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i27_2_lut (.I0(IntegralLimit[13]), .I1(n233[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(n233[4]), .I1(n285[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5181));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(n233[5]), .I1(n285[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5184));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(n233[6]), .I1(n285[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5183));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(n233[7]), .I1(n285[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5182));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(n233[9]), .I1(n285[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5179));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(n233[8]), .I1(n285[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5180));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(n233[11]), .I1(n285[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5205));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(n233[12]), .I1(n285[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5204));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_5219), 
            .I3(GND_net), .O(n8_adj_5282));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n79267), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16_adj_5280), .I1(n535[22]), .I2(n45_adj_5210), 
            .I3(GND_net), .O(n24_adj_5283));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0_i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n79261), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i60176_4_lut (.I0(n43_adj_5211), .I1(n25_adj_5216), .I2(n23_adj_5215), 
            .I3(n76084), .O(n76032));
    defparam i60176_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62193_3_lut (.I0(n78048), .I1(n233[23]), .I2(n285[23]), .I3(GND_net), 
            .O(n284));   // verilog/motorControl.v(58[23:46])
    defparam i62193_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_add_1225_24_lut (.I0(n336), .I1(n13005[21]), .I2(GND_net), 
            .I3(n60586), .O(n12498[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_add_1225_23_lut (.I0(GND_net), .I1(n13005[20]), .I2(GND_net), 
            .I3(n60585), .O(n46[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_23 (.CI(n60585), .I0(n13005[20]), .I1(GND_net), 
            .CO(n60586));
    SB_LUT4 mult_24_add_1225_22_lut (.I0(GND_net), .I1(n13005[19]), .I2(GND_net), 
            .I3(n60584), .O(n46[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61695_4_lut (.I0(n24_adj_5283), .I1(n8_adj_5282), .I2(n45_adj_5210), 
            .I3(n76026), .O(n77551));   // verilog/motorControl.v(47[25:43])
    defparam i61695_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60597_3_lut (.I0(n77732), .I1(n535[12]), .I2(n25_adj_5216), 
            .I3(GND_net), .O(n76453));   // verilog/motorControl.v(47[25:43])
    defparam i60597_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_22 (.CI(n60584), .I0(n13005[19]), .I1(GND_net), 
            .CO(n60585));
    SB_LUT4 mult_24_add_1225_21_lut (.I0(GND_net), .I1(n13005[18]), .I2(GND_net), 
            .I3(n60583), .O(n46[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_21 (.CI(n60583), .I0(n13005[18]), .I1(GND_net), 
            .CO(n60584));
    SB_LUT4 mult_24_add_1225_20_lut (.I0(GND_net), .I1(n13005[17]), .I2(GND_net), 
            .I3(n60582), .O(n46[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_20 (.CI(n60582), .I0(n13005[17]), .I1(GND_net), 
            .CO(n60583));
    SB_LUT4 mult_24_add_1225_19_lut (.I0(GND_net), .I1(n13005[16]), .I2(GND_net), 
            .I3(n60581), .O(n46[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_19 (.CI(n60581), .I0(n13005[16]), .I1(GND_net), 
            .CO(n60582));
    SB_LUT4 mult_24_add_1225_18_lut (.I0(GND_net), .I1(n13005[15]), .I2(GND_net), 
            .I3(n60580), .O(n46[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_18 (.CI(n60580), .I0(n13005[15]), .I1(GND_net), 
            .CO(n60581));
    SB_LUT4 LessThan_11_i4_4_lut (.I0(setpoint[0]), .I1(n535[1]), .I2(setpoint[1]), 
            .I3(n535[0]), .O(n4_adj_5284));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61873_3_lut (.I0(n4_adj_5284), .I1(n535[13]), .I2(n27_adj_5255), 
            .I3(GND_net), .O(n77729));   // verilog/motorControl.v(47[25:43])
    defparam i61873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61874_3_lut (.I0(n77729), .I1(n535[14]), .I2(n29_adj_5212), 
            .I3(GND_net), .O(n77730));   // verilog/motorControl.v(47[25:43])
    defparam i61874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_17_lut (.I0(GND_net), .I1(n13005[14]), .I2(GND_net), 
            .I3(n60579), .O(n46[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60192_4_lut (.I0(n33_adj_5222), .I1(n31_adj_5213), .I2(n29_adj_5212), 
            .I3(n76058), .O(n76048));
    defparam i60192_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mult_24_add_1225_17 (.CI(n60579), .I0(n13005[14]), .I1(GND_net), 
            .CO(n60580));
    SB_LUT4 mult_24_add_1225_16_lut (.I0(GND_net), .I1(n13005[13]), .I2(n1096_adj_5158), 
            .I3(n60578), .O(n46[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_16 (.CI(n60578), .I0(n13005[13]), .I1(n1096_adj_5158), 
            .CO(n60579));
    SB_LUT4 mult_24_add_1225_15_lut (.I0(GND_net), .I1(n13005[12]), .I2(n1023_adj_5157), 
            .I3(n60577), .O(n46[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59550_2_lut (.I0(PWMLimit[0]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75241));
    defparam i59550_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_15 (.CI(n60577), .I0(n13005[12]), .I1(n1023_adj_5157), 
            .CO(n60578));
    SB_LUT4 mult_24_add_1225_14_lut (.I0(GND_net), .I1(n13005[11]), .I2(n950_adj_5156), 
            .I3(n60576), .O(n46[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62207_4_lut (.I0(n30_adj_5279), .I1(n10_adj_5278), .I2(n35_adj_5217), 
            .I3(n76044), .O(n78063));   // verilog/motorControl.v(47[25:43])
    defparam i62207_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY mult_24_add_1225_14 (.CI(n60576), .I0(n13005[11]), .I1(n950_adj_5156), 
            .CO(n60577));
    SB_LUT4 mult_24_add_1225_13_lut (.I0(GND_net), .I1(n13005[10]), .I2(n877_adj_5155), 
            .I3(n60575), .O(n46[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_13 (.CI(n60575), .I0(n13005[10]), .I1(n877_adj_5155), 
            .CO(n60576));
    SB_LUT4 mult_24_add_1225_12_lut (.I0(GND_net), .I1(n13005[9]), .I2(n804_adj_5154), 
            .I3(n60574), .O(n46[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_12 (.CI(n60574), .I0(n13005[9]), .I1(n804_adj_5154), 
            .CO(n60575));
    SB_LUT4 mult_24_add_1225_11_lut (.I0(GND_net), .I1(n13005[8]), .I2(n731_adj_5153), 
            .I3(n60573), .O(n46[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_11 (.CI(n60573), .I0(n13005[8]), .I1(n731_adj_5153), 
            .CO(n60574));
    SB_LUT4 mult_24_add_1225_10_lut (.I0(GND_net), .I1(n13005[7]), .I2(n658_adj_5152), 
            .I3(n60572), .O(n46[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_10 (.CI(n60572), .I0(n13005[7]), .I1(n658_adj_5152), 
            .CO(n60573));
    SB_LUT4 i59862_2_lut (.I0(PWMLimit[1]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75254));
    defparam i59862_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60599_3_lut (.I0(n77730), .I1(n535[15]), .I2(n31_adj_5213), 
            .I3(GND_net), .O(n76455));   // verilog/motorControl.v(47[25:43])
    defparam i60599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62361_4_lut (.I0(n76455), .I1(n78063), .I2(n35_adj_5217), 
            .I3(n76048), .O(n78217));   // verilog/motorControl.v(47[25:43])
    defparam i62361_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_add_1225_9_lut (.I0(GND_net), .I1(n13005[6]), .I2(n585_adj_5151), 
            .I3(n60571), .O(n46[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_9 (.CI(n60571), .I0(n13005[6]), .I1(n585_adj_5151), 
            .CO(n60572));
    SB_LUT4 mult_24_add_1225_8_lut (.I0(GND_net), .I1(n13005[5]), .I2(n512_adj_5149), 
            .I3(n60570), .O(n46[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_8 (.CI(n60570), .I0(n13005[5]), .I1(n512_adj_5149), 
            .CO(n60571));
    SB_LUT4 i59748_2_lut (.I0(PWMLimit[16]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75287));
    defparam i59748_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59648_2_lut (.I0(PWMLimit[17]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75288));
    defparam i59648_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i62362_3_lut (.I0(n78217), .I1(n535[18]), .I2(n37_adj_5214), 
            .I3(GND_net), .O(n78218));   // verilog/motorControl.v(47[25:43])
    defparam i62362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_7_lut (.I0(GND_net), .I1(n13005[4]), .I2(n439), 
            .I3(n60569), .O(n46[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_7 (.CI(n60569), .I0(n13005[4]), .I1(n439), 
            .CO(n60570));
    SB_LUT4 i59799_2_lut (.I0(PWMLimit[2]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75255));
    defparam i59799_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59790_2_lut (.I0(PWMLimit[18]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75289));
    defparam i59790_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_6_lut (.I0(GND_net), .I1(n13005[3]), .I2(n366), 
            .I3(n60568), .O(n46[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_6 (.CI(n60568), .I0(n13005[3]), .I1(n366), 
            .CO(n60569));
    SB_LUT4 mult_24_add_1225_5_lut (.I0(GND_net), .I1(n13005[2]), .I2(n293), 
            .I3(n60567), .O(n46[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59635_2_lut (.I0(PWMLimit[3]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75256));
    defparam i59635_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_5 (.CI(n60567), .I0(n13005[2]), .I1(n293), 
            .CO(n60568));
    SB_LUT4 mult_24_add_1225_4_lut (.I0(GND_net), .I1(n13005[1]), .I2(n220), 
            .I3(n60566), .O(n46[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_4 (.CI(n60566), .I0(n13005[1]), .I1(n220), 
            .CO(n60567));
    SB_LUT4 i59710_2_lut (.I0(PWMLimit[19]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75291));
    defparam i59710_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59789_2_lut (.I0(PWMLimit[20]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75292));
    defparam i59789_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59798_2_lut (.I0(PWMLimit[4]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75257));
    defparam i59798_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_3_lut (.I0(GND_net), .I1(n13005[0]), .I2(n147), 
            .I3(n60565), .O(n46[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_3 (.CI(n60565), .I0(n13005[0]), .I1(n147), 
            .CO(n60566));
    SB_LUT4 i59782_2_lut (.I0(PWMLimit[21]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75293));
    defparam i59782_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74_adj_5146), 
            .I3(GND_net), .O(n46[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74_adj_5146), 
            .CO(n60565));
    SB_LUT4 i59788_2_lut (.I0(PWMLimit[22]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75294));
    defparam i59788_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6189_23_lut (.I0(GND_net), .I1(n13970[20]), .I2(GND_net), 
            .I3(n60564), .O(n13005[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6189_22_lut (.I0(GND_net), .I1(n13970[19]), .I2(GND_net), 
            .I3(n60563), .O(n13005[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_22 (.CI(n60563), .I0(n13970[19]), .I1(GND_net), 
            .CO(n60564));
    SB_LUT4 add_6189_21_lut (.I0(GND_net), .I1(n13970[18]), .I2(GND_net), 
            .I3(n60562), .O(n13005[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_21 (.CI(n60562), .I0(n13970[18]), .I1(GND_net), 
            .CO(n60563));
    SB_LUT4 add_6189_20_lut (.I0(GND_net), .I1(n13970[17]), .I2(GND_net), 
            .I3(n60561), .O(n13005[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_20 (.CI(n60561), .I0(n13970[17]), .I1(GND_net), 
            .CO(n60562));
    SB_LUT4 add_6189_19_lut (.I0(GND_net), .I1(n13970[16]), .I2(GND_net), 
            .I3(n60560), .O(n13005[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62334_3_lut (.I0(n78218), .I1(n535[19]), .I2(n39_adj_5209), 
            .I3(GND_net), .O(n78190));   // verilog/motorControl.v(47[25:43])
    defparam i62334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60178_4_lut (.I0(n43_adj_5211), .I1(n41_adj_5208), .I2(n39_adj_5209), 
            .I3(n78136), .O(n76034));
    defparam i60178_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62182_4_lut (.I0(n76453), .I1(n77551), .I2(n45_adj_5210), 
            .I3(n76032), .O(n78038));   // verilog/motorControl.v(47[25:43])
    defparam i62182_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_add_1221_24_lut (.I0(n207[23]), .I1(n12381[21]), .I2(GND_net), 
            .I3(n59643), .O(n11922[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6189_19 (.CI(n60560), .I0(n13970[16]), .I1(GND_net), 
            .CO(n60561));
    SB_LUT4 add_6189_18_lut (.I0(GND_net), .I1(n13970[15]), .I2(GND_net), 
            .I3(n60559), .O(n13005[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_23_lut (.I0(GND_net), .I1(n12381[20]), .I2(GND_net), 
            .I3(n59642), .O(n360[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_23 (.CI(n59642), .I0(n12381[20]), .I1(GND_net), 
            .CO(n59643));
    SB_LUT4 i60605_3_lut (.I0(n78190), .I1(n535[20]), .I2(n41_adj_5208), 
            .I3(GND_net), .O(n76461));   // verilog/motorControl.v(47[25:43])
    defparam i60605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n20492[1]), .I1(n4_adj_5288), .I2(n277), .I3(GND_net), 
            .O(n20464[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mult_24_i281_2_lut (.I0(\Ki[5] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59636_2_lut (.I0(PWMLimit[5]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75258));
    defparam i59636_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6189_18 (.CI(n60559), .I0(n13970[15]), .I1(GND_net), 
            .CO(n60560));
    SB_LUT4 add_6189_17_lut (.I0(GND_net), .I1(n13970[14]), .I2(GND_net), 
            .I3(n60558), .O(n13005[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_17 (.CI(n60558), .I0(n13970[14]), .I1(GND_net), 
            .CO(n60559));
    SB_LUT4 add_6189_16_lut (.I0(GND_net), .I1(n13970[13]), .I2(n1099), 
            .I3(n60557), .O(n13005[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_16 (.CI(n60557), .I0(n13970[13]), .I1(n1099), .CO(n60558));
    SB_LUT4 add_6189_15_lut (.I0(GND_net), .I1(n13970[12]), .I2(n1026), 
            .I3(n60556), .O(n13005[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_15 (.CI(n60556), .I0(n13970[12]), .I1(n1026), .CO(n60557));
    SB_LUT4 add_6189_14_lut (.I0(GND_net), .I1(n13970[11]), .I2(n953), 
            .I3(n60555), .O(n13005[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_14 (.CI(n60555), .I0(n13970[11]), .I1(n953), .CO(n60556));
    SB_LUT4 mult_24_i330_2_lut (.I0(\Ki[6] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(n337), .I3(n336), 
            .O(n71504));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut.LUT_INIT = 16'h93a0;
    SB_LUT4 mult_23_add_1221_22_lut (.I0(GND_net), .I1(n12381[19]), .I2(GND_net), 
            .I3(n59641), .O(n360[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n37307), .I1(\Ki[4] ), .I2(\Ki[5] ), 
            .I3(n340), .O(n71508));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'h6ca0;
    SB_LUT4 i62184_4_lut (.I0(n76461), .I1(n78038), .I2(n45_adj_5210), 
            .I3(n76034), .O(n78040));   // verilog/motorControl.v(47[25:43])
    defparam i62184_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(\Ki[3] ), .I1(n37117), .I2(n339), .I3(\Ki[2] ), 
            .O(n71506));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'h6ca0;
    SB_CARRY mult_23_add_1221_22 (.CI(n59641), .I0(n12381[19]), .I1(GND_net), 
            .CO(n59642));
    SB_LUT4 add_6189_13_lut (.I0(GND_net), .I1(n13970[10]), .I2(n880), 
            .I3(n60554), .O(n13005[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62185_3_lut (.I0(n78040), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(47[25:43])
    defparam i62185_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_6189_13 (.CI(n60554), .I0(n13970[10]), .I1(n880), .CO(n60555));
    SB_LUT4 i1_3_lut_adj_1787 (.I0(n71506), .I1(n71508), .I2(n71504), 
            .I3(GND_net), .O(n71512));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_adj_1787.LUT_INIT = 16'h9696;
    SB_LUT4 add_6189_12_lut (.I0(GND_net), .I1(n13970[9]), .I2(n807), 
            .I3(n60553), .O(n13005[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_12 (.CI(n60553), .I0(n13970[9]), .I1(n807), .CO(n60554));
    SB_LUT4 LessThan_32_i33_2_lut (.I0(n455[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5289));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6189_11_lut (.I0(GND_net), .I1(n13970[8]), .I2(n734), 
            .I3(n60552), .O(n13005[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i11_2_lut (.I0(n455[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5290));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6189_11 (.CI(n60552), .I0(n13970[8]), .I1(n734), .CO(n60553));
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n4_adj_5291), .I1(n71512), .I2(n68_adj_5292), 
            .I3(n137), .O(n71516));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'h9666;
    SB_LUT4 LessThan_32_i13_2_lut (.I0(n455[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5293));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n20492[1]), .I1(n71516), .I2(n277), 
            .I3(n4_adj_5288), .O(n71518));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'h366c;
    SB_LUT4 add_6189_10_lut (.I0(GND_net), .I1(n13970[7]), .I2(n661), 
            .I3(n60551), .O(n13005[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11882_bdd_4_lut_63423 (.I0(n11882), .I1(n75264), .I2(setpoint[11]), 
            .I3(n4736), .O(n79312));
    defparam n11882_bdd_4_lut_63423.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_add_1221_21_lut (.I0(GND_net), .I1(n12381[18]), .I2(GND_net), 
            .I3(n59640), .O(n360[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_10 (.CI(n60551), .I0(n13970[7]), .I1(n661), .CO(n60552));
    SB_LUT4 add_6189_9_lut (.I0(GND_net), .I1(n13970[6]), .I2(n588), .I3(n60550), 
            .O(n13005[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_9 (.CI(n60550), .I0(n13970[6]), .I1(n588), .CO(n60551));
    SB_LUT4 add_6189_8_lut (.I0(GND_net), .I1(n13970[5]), .I2(n515), .I3(n60549), 
            .O(n13005[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_8 (.CI(n60549), .I0(n13970[5]), .I1(n515), .CO(n60550));
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n71518), .I1(n20464[2]), .I2(n347), 
            .I3(n6), .O(n69694));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'h566a;
    SB_LUT4 i1_3_lut_adj_1791 (.I0(n20464[2]), .I1(n6), .I2(n347), .I3(GND_net), 
            .O(n20418[3]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_adj_1791.LUT_INIT = 16'h9696;
    SB_LUT4 add_6189_7_lut (.I0(GND_net), .I1(n13970[4]), .I2(n442), .I3(n60548), 
            .O(n13005[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_7 (.CI(n60548), .I0(n13970[4]), .I1(n442), .CO(n60549));
    SB_LUT4 add_6189_6_lut (.I0(GND_net), .I1(n13970[3]), .I2(n369), .I3(n60547), 
            .O(n13005[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_6 (.CI(n60547), .I0(n13970[3]), .I1(n369), .CO(n60548));
    SB_LUT4 add_6189_5_lut (.I0(GND_net), .I1(n13970[2]), .I2(n296_adj_5140), 
            .I3(n60546), .O(n13005[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_5 (.CI(n60546), .I0(n13970[2]), .I1(n296_adj_5140), 
            .CO(n60547));
    SB_LUT4 add_6189_4_lut (.I0(GND_net), .I1(n13970[1]), .I2(n223), .I3(n60545), 
            .O(n13005[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i15_2_lut (.I0(n455[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5295));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6189_4 (.CI(n60545), .I0(n13970[1]), .I1(n223), .CO(n60546));
    SB_LUT4 add_6189_3_lut (.I0(GND_net), .I1(n13970[0]), .I2(n150), .I3(n60544), 
            .O(n13005[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_3 (.CI(n60544), .I0(n13970[0]), .I1(n150), .CO(n60545));
    SB_LUT4 add_6189_2_lut (.I0(GND_net), .I1(n8_adj_5138), .I2(n77), 
            .I3(GND_net), .O(n13005[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_21 (.CI(n59640), .I0(n12381[18]), .I1(GND_net), 
            .CO(n59641));
    SB_CARRY add_6189_2 (.CI(GND_net), .I0(n8_adj_5138), .I1(n77), .CO(n60544));
    SB_LUT4 add_6232_22_lut (.I0(GND_net), .I1(n14848[19]), .I2(GND_net), 
            .I3(n60543), .O(n13970[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6232_21_lut (.I0(GND_net), .I1(n14848[18]), .I2(GND_net), 
            .I3(n60542), .O(n13970[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i69_2_lut (.I0(\Kp[1] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i22_2_lut (.I0(\Kp[0] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i118_2_lut (.I0(\Kp[2] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_20_lut (.I0(GND_net), .I1(n12381[17]), .I2(GND_net), 
            .I3(n59639), .O(n360[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i167_2_lut (.I0(\Kp[3] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_5296));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i216_2_lut (.I0(\Kp[4] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6232_21 (.CI(n60542), .I0(n14848[18]), .I1(GND_net), 
            .CO(n60543));
    SB_LUT4 add_6232_20_lut (.I0(GND_net), .I1(n14848[17]), .I2(GND_net), 
            .I3(n60541), .O(n13970[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i265_2_lut (.I0(\Kp[5] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i27_2_lut (.I0(n455[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5297));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i21_2_lut (.I0(deadband[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5298));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_23_add_1221_20 (.CI(n59639), .I0(n12381[17]), .I1(GND_net), 
            .CO(n59640));
    SB_LUT4 mult_23_add_1221_19_lut (.I0(GND_net), .I1(n12381[16]), .I2(GND_net), 
            .I3(n59638), .O(n360[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_20 (.CI(n60541), .I0(n14848[17]), .I1(GND_net), 
            .CO(n60542));
    SB_LUT4 LessThan_26_i4_4_lut (.I0(deadband[0]), .I1(n455[1]), .I2(deadband[1]), 
            .I3(n455[0]), .O(n4_adj_5299));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_16_14 (.CI(n58942), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n207[16]), .CO(n58943));
    SB_LUT4 add_6232_19_lut (.I0(GND_net), .I1(n14848[16]), .I2(GND_net), 
            .I3(n60540), .O(n13970[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_19 (.CI(n60540), .I0(n14848[16]), .I1(GND_net), 
            .CO(n60541));
    SB_CARRY mult_23_add_1221_19 (.CI(n59638), .I0(n12381[16]), .I1(GND_net), 
            .CO(n59639));
    SB_LUT4 mult_23_i314_2_lut (.I0(\Kp[6] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_5300));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_18_lut (.I0(GND_net), .I1(n12381[15]), .I2(GND_net), 
            .I3(n59637), .O(n360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i363_2_lut (.I0(\Kp[7] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_5301));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_18 (.CI(n59637), .I0(n12381[15]), .I1(GND_net), 
            .CO(n59638));
    SB_LUT4 add_6232_18_lut (.I0(GND_net), .I1(n14848[15]), .I2(GND_net), 
            .I3(n60539), .O(n13970[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61701_3_lut (.I0(n4_adj_5299), .I1(n455[2]), .I2(deadband[2]), 
            .I3(GND_net), .O(n77557));   // verilog/motorControl.v(62[14:31])
    defparam i61701_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i412_2_lut (.I0(\Kp[8] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61702_3_lut (.I0(n77557), .I1(n455[3]), .I2(deadband[3]), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(62[14:31])
    defparam i61702_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6232_18 (.CI(n60539), .I0(n14848[15]), .I1(GND_net), 
            .CO(n60540));
    SB_LUT4 add_6232_17_lut (.I0(GND_net), .I1(n14848[14]), .I2(GND_net), 
            .I3(n60538), .O(n13970[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i461_2_lut (.I0(\Kp[9] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6232_17 (.CI(n60538), .I0(n14848[14]), .I1(GND_net), 
            .CO(n60539));
    SB_LUT4 LessThan_26_i19_2_lut (.I0(deadband[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5305));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(deadband[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5306));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6232_16_lut (.I0(GND_net), .I1(n14848[13]), .I2(n1102), 
            .I3(n60537), .O(n13970[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6232_16 (.CI(n60537), .I0(n14848[13]), .I1(n1102), .CO(n60538));
    SB_LUT4 add_6232_15_lut (.I0(GND_net), .I1(n14848[12]), .I2(n1029), 
            .I3(n60536), .O(n13970[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(deadband[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5308));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6232_15 (.CI(n60536), .I0(n14848[12]), .I1(n1029), .CO(n60537));
    SB_LUT4 add_6232_14_lut (.I0(GND_net), .I1(n14848[11]), .I2(n956), 
            .I3(n60535), .O(n13970[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_14 (.CI(n60535), .I0(n14848[11]), .I1(n956), .CO(n60536));
    SB_LUT4 add_6232_13_lut (.I0(GND_net), .I1(n14848[10]), .I2(n883), 
            .I3(n60534), .O(n13970[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_13 (.CI(n60534), .I0(n14848[10]), .I1(n883), .CO(n60535));
    SB_LUT4 add_6232_12_lut (.I0(GND_net), .I1(n14848[9]), .I2(n810), 
            .I3(n60533), .O(n13970[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_12 (.CI(n60533), .I0(n14848[9]), .I1(n810), .CO(n60534));
    SB_LUT4 add_6232_11_lut (.I0(GND_net), .I1(n14848[8]), .I2(n737), 
            .I3(n60532), .O(n13970[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i510_2_lut (.I0(\Kp[10] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_17_lut (.I0(GND_net), .I1(n12381[14]), .I2(GND_net), 
            .I3(n59636), .O(n360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_11 (.CI(n60532), .I0(n14848[8]), .I1(n737), .CO(n60533));
    SB_CARRY mult_23_add_1221_17 (.CI(n59636), .I0(n12381[14]), .I1(GND_net), 
            .CO(n59637));
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6232_10_lut (.I0(GND_net), .I1(n14848[7]), .I2(n664), 
            .I3(n60531), .O(n13970[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i559_2_lut (.I0(\Kp[11] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6232_10 (.CI(n60531), .I0(n14848[7]), .I1(n664), .CO(n60532));
    SB_LUT4 mult_23_i608_2_lut (.I0(\Kp[12] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6232_9_lut (.I0(GND_net), .I1(n14848[6]), .I2(n591), .I3(n60530), 
            .O(n13970[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_9 (.CI(n60530), .I0(n14848[6]), .I1(n591), .CO(n60531));
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6232_8_lut (.I0(GND_net), .I1(n14848[5]), .I2(n518), .I3(n60529), 
            .O(n13970[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_8 (.CI(n60529), .I0(n14848[5]), .I1(n518), .CO(n60530));
    SB_LUT4 LessThan_26_i15_2_lut (.I0(deadband[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5311));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6232_7_lut (.I0(GND_net), .I1(n14848[4]), .I2(n445), .I3(n60528), 
            .O(n13970[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_16_lut (.I0(GND_net), .I1(n12381[13]), .I2(n1096), 
            .I3(n59635), .O(n360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i657_2_lut (.I0(\Kp[13] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_23_add_1221_16 (.CI(n59635), .I0(n12381[13]), .I1(n1096), 
            .CO(n59636));
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i706_2_lut (.I0(\Kp[14] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(deadband[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5314));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i11_2_lut (.I0(deadband[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5315));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i60022_4_lut (.I0(n17_adj_5314), .I1(n15_adj_5311), .I2(n13_adj_5308), 
            .I3(n11_adj_5315), .O(n75878));
    defparam i60022_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6232_7 (.CI(n60528), .I0(n14848[4]), .I1(n445), .CO(n60529));
    SB_LUT4 add_6232_6_lut (.I0(GND_net), .I1(n14848[3]), .I2(n372), .I3(n60527), 
            .O(n13970[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_6 (.CI(n60527), .I0(n14848[3]), .I1(n372), .CO(n60528));
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6232_5_lut (.I0(GND_net), .I1(n14848[2]), .I2(n299_c), 
            .I3(n60526), .O(n13970[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_15_lut (.I0(GND_net), .I1(n12381[12]), .I2(n1023), 
            .I3(n59634), .O(n360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_15 (.CI(n59634), .I0(n12381[12]), .I1(n1023), 
            .CO(n59635));
    SB_LUT4 add_16_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n207[15]), .I3(n58941), .O(n233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_14_lut (.I0(GND_net), .I1(n12381[11]), .I2(n950), 
            .I3(n59633), .O(n360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i67_2_lut (.I0(\Kp[1] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6232_5 (.CI(n60526), .I0(n14848[2]), .I1(n299_c), .CO(n60527));
    SB_LUT4 add_6232_4_lut (.I0(GND_net), .I1(n14848[1]), .I2(n226), .I3(n60525), 
            .O(n13970[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_4 (.CI(n60525), .I0(n14848[1]), .I1(n226), .CO(n60526));
    SB_CARRY mult_23_add_1221_14 (.CI(n59633), .I0(n12381[11]), .I1(n950), 
            .CO(n59634));
    SB_CARRY add_16_13 (.CI(n58941), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n207[15]), .CO(n58942));
    SB_LUT4 add_6232_3_lut (.I0(GND_net), .I1(n14848[0]), .I2(n153), .I3(n60524), 
            .O(n13970[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n207[14]), .I3(n58940), .O(n247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i14_3_lut (.I0(n455[7]), .I1(n455[11]), .I2(n23_adj_5306), 
            .I3(GND_net), .O(n14_adj_5316));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6232_3 (.CI(n60524), .I0(n14848[0]), .I1(n153), .CO(n60525));
    SB_LUT4 mult_23_i20_2_lut (.I0(\Kp[0] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5317));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6232_2_lut (.I0(GND_net), .I1(n11_adj_5137), .I2(n80), 
            .I3(GND_net), .O(n13970[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_2 (.CI(GND_net), .I0(n11_adj_5137), .I1(n80), .CO(n60524));
    SB_LUT4 add_6529_12_lut (.I0(GND_net), .I1(n19637[9]), .I2(n840), 
            .I3(n60523), .O(n19374[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6529_11_lut (.I0(GND_net), .I1(n19637[8]), .I2(n767), 
            .I3(n60522), .O(n19374[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i116_2_lut (.I0(\Kp[2] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6529_11 (.CI(n60522), .I0(n19637[8]), .I1(n767), .CO(n60523));
    SB_LUT4 mult_23_i165_2_lut (.I0(\Kp[3] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_5318));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_5308), 
            .I3(GND_net), .O(n12_adj_5319));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6529_10_lut (.I0(GND_net), .I1(n19637[7]), .I2(n694), 
            .I3(n60521), .O(n19374[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_13_lut (.I0(GND_net), .I1(n12381[10]), .I2(n877), 
            .I3(n59632), .O(n360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_10 (.CI(n60521), .I0(n19637[7]), .I1(n694), .CO(n60522));
    SB_LUT4 mult_23_i214_2_lut (.I0(\Kp[4] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6529_9_lut (.I0(GND_net), .I1(n19637[6]), .I2(n621), .I3(n60520), 
            .O(n19374[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i22_3_lut (.I0(n14_adj_5316), .I1(n467), .I2(n25_adj_28), 
            .I3(GND_net), .O(n22_adj_5321));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i16_3_lut (.I0(n455[8]), .I1(n455[9]), .I2(n19_adj_5305), 
            .I3(GND_net), .O(n16_adj_5322));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i263_2_lut (.I0(\Kp[5] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_5323));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i312_2_lut (.I0(\Kp[6] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_5324));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_13 (.CI(n59632), .I0(n12381[10]), .I1(n877), 
            .CO(n59633));
    SB_LUT4 mult_23_add_1221_12_lut (.I0(GND_net), .I1(n12381[9]), .I2(n804), 
            .I3(n59631), .O(n360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i361_2_lut (.I0(\Kp[7] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_5326));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6529_9 (.CI(n60520), .I0(n19637[6]), .I1(n621), .CO(n60521));
    SB_CARRY add_16_12 (.CI(n58940), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n207[14]), .CO(n58941));
    SB_CARRY mult_23_add_1221_12 (.CI(n59631), .I0(n12381[9]), .I1(n804), 
            .CO(n59632));
    SB_LUT4 mult_23_add_1221_11_lut (.I0(GND_net), .I1(n12381[8]), .I2(n731), 
            .I3(n59630), .O(n360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6529_8_lut (.I0(GND_net), .I1(n19637[5]), .I2(n548), .I3(n60519), 
            .O(n19374[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i410_2_lut (.I0(\Kp[8] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i410_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6529_8 (.CI(n60519), .I0(n19637[5]), .I1(n548), .CO(n60520));
    SB_CARRY mult_23_add_1221_11 (.CI(n59630), .I0(n12381[8]), .I1(n731), 
            .CO(n59631));
    SB_LUT4 mult_23_add_1221_10_lut (.I0(GND_net), .I1(n12381[7]), .I2(n658), 
            .I3(n59629), .O(n360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i459_2_lut (.I0(\Kp[9] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_10 (.CI(n59629), .I0(n12381[7]), .I1(n658), 
            .CO(n59630));
    SB_LUT4 mult_23_add_1221_9_lut (.I0(GND_net), .I1(n12381[6]), .I2(n585), 
            .I3(n59628), .O(n360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6529_7_lut (.I0(GND_net), .I1(n19637[4]), .I2(n475_c), 
            .I3(n60518), .O(n19374[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_7 (.CI(n60518), .I0(n19637[4]), .I1(n475_c), .CO(n60519));
    SB_LUT4 mult_23_i508_2_lut (.I0(\Kp[10] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6529_6_lut (.I0(GND_net), .I1(n19637[3]), .I2(n402), .I3(n60517), 
            .O(n19374[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_9 (.CI(n59628), .I0(n12381[6]), .I1(n585), 
            .CO(n59629));
    SB_LUT4 mult_23_add_1221_8_lut (.I0(GND_net), .I1(n12381[5]), .I2(n512), 
            .I3(n59627), .O(n360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i557_2_lut (.I0(\Kp[11] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6529_6 (.CI(n60517), .I0(n19637[3]), .I1(n402), .CO(n60518));
    SB_LUT4 add_6529_5_lut (.I0(GND_net), .I1(n19637[2]), .I2(n329), .I3(n60516), 
            .O(n19374[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_5 (.CI(n60516), .I0(n19637[2]), .I1(n329), .CO(n60517));
    SB_LUT4 mult_23_i606_2_lut (.I0(\Kp[12] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i655_2_lut (.I0(\Kp[13] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6529_4_lut (.I0(GND_net), .I1(n19637[1]), .I2(n256_adj_5136), 
            .I3(n60515), .O(n19374[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_8 (.CI(n59627), .I0(n12381[5]), .I1(n512), 
            .CO(n59628));
    SB_LUT4 mult_23_i704_2_lut (.I0(\Kp[14] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i704_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6529_4 (.CI(n60515), .I0(n19637[1]), .I1(n256_adj_5136), 
            .CO(n60516));
    SB_LUT4 add_6529_3_lut (.I0(GND_net), .I1(n19637[0]), .I2(n183), .I3(n60514), 
            .O(n19374[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_3 (.CI(n60514), .I0(n19637[0]), .I1(n183), .CO(n60515));
    SB_LUT4 mult_23_i753_2_lut (.I0(\Kp[15] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i83_2_lut (.I0(\Ki[1] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n79312_bdd_4_lut (.I0(n79312), .I1(n535[11]), .I2(n455[11]), 
            .I3(n4736), .O(n79315));
    defparam n79312_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i36_2_lut (.I0(\Ki[0] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6529_2_lut (.I0(GND_net), .I1(n41_adj_5328), .I2(n110_c), 
            .I3(GND_net), .O(n19374[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_2 (.CI(GND_net), .I0(n41_adj_5328), .I1(n110_c), 
            .CO(n60514));
    SB_LUT4 mult_24_i132_2_lut (.I0(\Ki[2] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_21_lut (.I0(GND_net), .I1(n15644[18]), .I2(GND_net), 
            .I3(n60513), .O(n14848[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6272_20_lut (.I0(GND_net), .I1(n15644[17]), .I2(GND_net), 
            .I3(n60512), .O(n14848[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_20 (.CI(n60512), .I0(n15644[17]), .I1(GND_net), 
            .CO(n60513));
    SB_LUT4 LessThan_26_i18_3_lut (.I0(n16_adj_5322), .I1(n455[10]), .I2(n21_adj_5298), 
            .I3(GND_net), .O(n18_adj_5329));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31217_1_lut (.I0(n455[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45309));   // verilog/motorControl.v(61[20:40])
    defparam i31217_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[0]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6272_19_lut (.I0(GND_net), .I1(n15644[16]), .I2(GND_net), 
            .I3(n60511), .O(n14848[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_19 (.CI(n60511), .I0(n15644[16]), .I1(GND_net), 
            .CO(n60512));
    SB_LUT4 i60006_4_lut (.I0(n23_adj_5306), .I1(n21_adj_5298), .I2(n19_adj_5305), 
            .I3(n75878), .O(n75862));
    defparam i60006_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62213_4_lut (.I0(n22_adj_5321), .I1(n12_adj_5319), .I2(n25_adj_28), 
            .I3(n75857), .O(n78069));   // verilog/motorControl.v(62[14:31])
    defparam i62213_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i181_2_lut (.I0(\Ki[3] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_18_lut (.I0(GND_net), .I1(n15644[15]), .I2(GND_net), 
            .I3(n60510), .O(n14848[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_18 (.CI(n60510), .I0(n15644[15]), .I1(GND_net), 
            .CO(n60511));
    SB_LUT4 i61703_4_lut (.I0(n18_adj_5329), .I1(n10), .I2(n21_adj_5298), 
            .I3(n75864), .O(n77559));   // verilog/motorControl.v(62[14:31])
    defparam i61703_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i44661_2_lut_4_lut (.I0(\Ki[0] ), .I1(n337), .I2(n37117), 
            .I3(\Ki[1] ), .O(n20501[0]));   // verilog/motorControl.v(61[29:40])
    defparam i44661_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_24_i230_2_lut (.I0(\Ki[4] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[1]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6272_17_lut (.I0(GND_net), .I1(n15644[14]), .I2(GND_net), 
            .I3(n60509), .O(n14848[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i279_2_lut (.I0(\Ki[5] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i279_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_17 (.CI(n60509), .I0(n15644[14]), .I1(GND_net), 
            .CO(n60510));
    SB_LUT4 add_6272_16_lut (.I0(GND_net), .I1(n15644[13]), .I2(n1105), 
            .I3(n60508), .O(n14848[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_16 (.CI(n60508), .I0(n15644[13]), .I1(n1105), .CO(n60509));
    SB_LUT4 add_16_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n207[13]), .I3(n58939), .O(n233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i328_2_lut (.I0(\Ki[6] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i62373_4_lut (.I0(n77559), .I1(n78069), .I2(n25_adj_28), .I3(n75862), 
            .O(n78229));   // verilog/motorControl.v(62[14:31])
    defparam i62373_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62374_3_lut (.I0(n78229), .I1(n455[13]), .I2(deadband[13]), 
            .I3(GND_net), .O(n78230));   // verilog/motorControl.v(62[14:31])
    defparam i62374_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6272_15_lut (.I0(GND_net), .I1(n15644[12]), .I2(n1032), 
            .I3(n60507), .O(n14848[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i377_2_lut (.I0(\Ki[7] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_15 (.CI(n60507), .I0(n15644[12]), .I1(n1032), .CO(n60508));
    SB_LUT4 unary_minus_27_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[2]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62319_3_lut (.I0(n78230), .I1(n455[14]), .I2(deadband[14]), 
            .I3(GND_net), .O(n78175));   // verilog/motorControl.v(62[14:31])
    defparam i62319_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6272_14_lut (.I0(GND_net), .I1(n15644[11]), .I2(n959), 
            .I3(n60506), .O(n14848[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_14 (.CI(n60506), .I0(n15644[11]), .I1(n959), .CO(n60507));
    SB_LUT4 add_6272_13_lut (.I0(GND_net), .I1(n15644[10]), .I2(n886), 
            .I3(n60505), .O(n14848[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61705_3_lut (.I0(n78175), .I1(n455[15]), .I2(deadband[15]), 
            .I3(GND_net), .O(n77561));   // verilog/motorControl.v(62[14:31])
    defparam i61705_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_6272_13 (.CI(n60505), .I0(n15644[10]), .I1(n886), .CO(n60506));
    SB_LUT4 i61706_3_lut (.I0(n77561), .I1(n455[16]), .I2(deadband[16]), 
            .I3(GND_net), .O(n34));   // verilog/motorControl.v(62[14:31])
    defparam i61706_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6272_12_lut (.I0(GND_net), .I1(n15644[9]), .I2(n813), 
            .I3(n60504), .O(n14848[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i41_2_lut (.I0(deadband[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5335));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i23_2_lut (.I0(n455[11]), .I1(n48[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5336));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6272_12 (.CI(n60504), .I0(n15644[9]), .I1(n813), .CO(n60505));
    SB_LUT4 add_6272_11_lut (.I0(GND_net), .I1(n15644[8]), .I2(n740), 
            .I3(n60503), .O(n14848[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[3]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6272_11 (.CI(n60503), .I0(n15644[8]), .I1(n740), .CO(n60504));
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[4]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[5]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_28_i25_2_lut (.I0(n467), .I1(n48[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5340));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[6]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6272_10_lut (.I0(GND_net), .I1(n15644[7]), .I2(n667), 
            .I3(n60502), .O(n14848[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11882_bdd_4_lut_63418 (.I0(n11882), .I1(n75263), .I2(setpoint[10]), 
            .I3(n4736), .O(n79306));
    defparam n11882_bdd_4_lut_63418.LUT_INIT = 16'he4aa;
    SB_CARRY add_6272_10 (.CI(n60502), .I0(n15644[7]), .I1(n667), .CO(n60503));
    SB_LUT4 add_6272_9_lut (.I0(GND_net), .I1(n15644[6]), .I2(n594), .I3(n60501), 
            .O(n14848[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_9 (.CI(n60501), .I0(n15644[6]), .I1(n594), .CO(n60502));
    SB_LUT4 add_6272_8_lut (.I0(GND_net), .I1(n15644[5]), .I2(n521), .I3(n60500), 
            .O(n14848[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_8 (.CI(n60500), .I0(n15644[5]), .I1(n521), .CO(n60501));
    SB_LUT4 add_6272_7_lut (.I0(GND_net), .I1(n15644[4]), .I2(n448_adj_5342), 
            .I3(n60499), .O(n14848[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n79306_bdd_4_lut (.I0(n79306), .I1(n535[10]), .I2(n455[10]), 
            .I3(n4736), .O(n79309));
    defparam n79306_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_28_i17_2_lut (.I0(n455[8]), .I1(n48[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5343));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6272_7 (.CI(n60499), .I0(n15644[4]), .I1(n448_adj_5342), 
            .CO(n60500));
    SB_LUT4 add_6272_6_lut (.I0(GND_net), .I1(n15644[3]), .I2(n375), .I3(n60498), 
            .O(n14848[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_6 (.CI(n60498), .I0(n15644[3]), .I1(n375), .CO(n60499));
    SB_LUT4 add_6272_5_lut (.I0(GND_net), .I1(n15644[2]), .I2(n302_adj_5344), 
            .I3(n60497), .O(n14848[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11882_bdd_4_lut_63413 (.I0(n11882), .I1(n75262), .I2(setpoint[9]), 
            .I3(n4736), .O(n79300));
    defparam n11882_bdd_4_lut_63413.LUT_INIT = 16'he4aa;
    SB_LUT4 n79300_bdd_4_lut (.I0(n79300), .I1(n535[9]), .I2(n455[9]), 
            .I3(n4736), .O(n79303));
    defparam n79300_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_28_i19_2_lut (.I0(n455[9]), .I1(n48[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5345));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i21_2_lut (.I0(n455[10]), .I1(n48[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5346));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6272_5 (.CI(n60497), .I0(n15644[2]), .I1(n302_adj_5344), 
            .CO(n60498));
    SB_LUT4 add_6272_4_lut (.I0(GND_net), .I1(n15644[1]), .I2(n229), .I3(n60496), 
            .O(n14848[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_4 (.CI(n60496), .I0(n15644[1]), .I1(n229), .CO(n60497));
    SB_LUT4 LessThan_28_i7_2_lut (.I0(n455[3]), .I1(n48[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5347));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6272_3_lut (.I0(GND_net), .I1(n15644[0]), .I2(n156), .I3(n60495), 
            .O(n14848[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_3 (.CI(n60495), .I0(n15644[0]), .I1(n156), .CO(n60496));
    SB_LUT4 add_6272_2_lut (.I0(GND_net), .I1(n14_adj_5348), .I2(n83), 
            .I3(GND_net), .O(n14848[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_2 (.CI(GND_net), .I0(n14_adj_5348), .I1(n83), .CO(n60495));
    SB_LUT4 add_6310_20_lut (.I0(GND_net), .I1(n16362[17]), .I2(GND_net), 
            .I3(n60494), .O(n15644[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6310_19_lut (.I0(GND_net), .I1(n16362[16]), .I2(GND_net), 
            .I3(n60493), .O(n15644[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i9_2_lut (.I0(n475), .I1(n48[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5349));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6310_19 (.CI(n60493), .I0(n16362[16]), .I1(GND_net), 
            .CO(n60494));
    SB_LUT4 add_6310_18_lut (.I0(GND_net), .I1(n16362[15]), .I2(GND_net), 
            .I3(n60492), .O(n15644[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_18 (.CI(n60492), .I0(n16362[15]), .I1(GND_net), 
            .CO(n60493));
    SB_LUT4 add_6310_17_lut (.I0(GND_net), .I1(n16362[14]), .I2(GND_net), 
            .I3(n60491), .O(n15644[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_17 (.CI(n60491), .I0(n16362[14]), .I1(GND_net), 
            .CO(n60492));
    SB_LUT4 LessThan_28_i11_2_lut (.I0(n455[5]), .I1(n48[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5350));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6310_16_lut (.I0(GND_net), .I1(n16362[13]), .I2(n1108), 
            .I3(n60490), .O(n15644[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_16 (.CI(n60490), .I0(n16362[13]), .I1(n1108), .CO(n60491));
    SB_LUT4 LessThan_28_i13_2_lut (.I0(n455[6]), .I1(n48[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5351));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6310_15_lut (.I0(GND_net), .I1(n16362[12]), .I2(n1035), 
            .I3(n60489), .O(n15644[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_15 (.CI(n60489), .I0(n16362[12]), .I1(n1035), .CO(n60490));
    SB_LUT4 add_6310_14_lut (.I0(GND_net), .I1(n16362[11]), .I2(n962), 
            .I3(n60488), .O(n15644[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_14 (.CI(n60488), .I0(n16362[11]), .I1(n962), .CO(n60489));
    SB_LUT4 add_6310_13_lut (.I0(GND_net), .I1(n16362[10]), .I2(n889), 
            .I3(n60487), .O(n15644[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_13 (.CI(n60487), .I0(n16362[10]), .I1(n889), .CO(n60488));
    SB_LUT4 add_6310_12_lut (.I0(GND_net), .I1(n16362[9]), .I2(n816), 
            .I3(n60486), .O(n15644[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_12 (.CI(n60486), .I0(n16362[9]), .I1(n816), .CO(n60487));
    SB_LUT4 add_6310_11_lut (.I0(GND_net), .I1(n16362[8]), .I2(n743), 
            .I3(n60485), .O(n15644[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i15_2_lut (.I0(n455[7]), .I1(n48[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5352));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6310_11 (.CI(n60485), .I0(n16362[8]), .I1(n743), .CO(n60486));
    SB_LUT4 add_6310_10_lut (.I0(GND_net), .I1(n16362[7]), .I2(n670), 
            .I3(n60484), .O(n15644[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_10 (.CI(n60484), .I0(n16362[7]), .I1(n670), .CO(n60485));
    SB_LUT4 add_6310_9_lut (.I0(GND_net), .I1(n16362[6]), .I2(n597), .I3(n60483), 
            .O(n15644[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_9 (.CI(n60483), .I0(n16362[6]), .I1(n597), .CO(n60484));
    SB_LUT4 add_6310_8_lut (.I0(GND_net), .I1(n16362[5]), .I2(n524), .I3(n60482), 
            .O(n15644[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_8 (.CI(n60482), .I0(n16362[5]), .I1(n524), .CO(n60483));
    SB_LUT4 add_6310_7_lut (.I0(GND_net), .I1(n16362[4]), .I2(n451_adj_5353), 
            .I3(n60481), .O(n15644[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_7 (.CI(n60481), .I0(n16362[4]), .I1(n451_adj_5353), 
            .CO(n60482));
    SB_LUT4 add_6310_6_lut (.I0(GND_net), .I1(n16362[3]), .I2(n378), .I3(n60480), 
            .O(n15644[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_6 (.CI(n60480), .I0(n16362[3]), .I1(n378), .CO(n60481));
    SB_LUT4 add_6310_5_lut (.I0(GND_net), .I1(n16362[2]), .I2(n305_adj_5354), 
            .I3(n60479), .O(n15644[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_5 (.CI(n60479), .I0(n16362[2]), .I1(n305_adj_5354), 
            .CO(n60480));
    SB_LUT4 LessThan_28_i27_2_lut (.I0(n455[13]), .I1(n48[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5355));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6310_4_lut (.I0(GND_net), .I1(n16362[1]), .I2(n232), .I3(n60478), 
            .O(n15644[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_7_lut (.I0(GND_net), .I1(n12381[4]), .I2(n439_adj_5356), 
            .I3(n59626), .O(n360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_4 (.CI(n60478), .I0(n16362[1]), .I1(n232), .CO(n60479));
    SB_CARRY mult_23_add_1221_7 (.CI(n59626), .I0(n12381[4]), .I1(n439_adj_5356), 
            .CO(n59627));
    SB_LUT4 add_6310_3_lut (.I0(GND_net), .I1(n16362[0]), .I2(n159), .I3(n60477), 
            .O(n15644[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_3 (.CI(n60477), .I0(n16362[0]), .I1(n159), .CO(n60478));
    SB_LUT4 add_6310_2_lut (.I0(GND_net), .I1(n17_adj_5357), .I2(n86), 
            .I3(GND_net), .O(n15644[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_2 (.CI(GND_net), .I0(n17_adj_5357), .I1(n86), .CO(n60477));
    SB_LUT4 add_6550_11_lut (.I0(GND_net), .I1(n19856[8]), .I2(n770), 
            .I3(n60476), .O(n19637[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_11 (.CI(n58939), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n207[13]), .CO(n58940));
    SB_LUT4 add_6550_10_lut (.I0(GND_net), .I1(n19856[7]), .I2(n697), 
            .I3(n60475), .O(n19637[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_10 (.CI(n60475), .I0(n19856[7]), .I1(n697), .CO(n60476));
    SB_LUT4 add_6550_9_lut (.I0(GND_net), .I1(n19856[6]), .I2(n624), .I3(n60474), 
            .O(n19637[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_9 (.CI(n60474), .I0(n19856[6]), .I1(n624), .CO(n60475));
    SB_LUT4 LessThan_28_i35_2_lut (.I0(n462), .I1(n48[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5358));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6550_8_lut (.I0(GND_net), .I1(n19856[5]), .I2(n551_adj_5359), 
            .I3(n60473), .O(n19637[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_8 (.CI(n60473), .I0(n19856[5]), .I1(n551_adj_5359), 
            .CO(n60474));
    SB_LUT4 add_6550_7_lut (.I0(GND_net), .I1(n19856[4]), .I2(n478_adj_5360), 
            .I3(n60472), .O(n19637[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_7 (.CI(n60472), .I0(n19856[4]), .I1(n478_adj_5360), 
            .CO(n60473));
    SB_LUT4 add_6550_6_lut (.I0(GND_net), .I1(n19856[3]), .I2(n405_adj_5361), 
            .I3(n60471), .O(n19637[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i29_2_lut (.I0(n455[14]), .I1(n48[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5362));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6550_6 (.CI(n60471), .I0(n19856[3]), .I1(n405_adj_5361), 
            .CO(n60472));
    SB_LUT4 add_6550_5_lut (.I0(GND_net), .I1(n19856[2]), .I2(n332_adj_5363), 
            .I3(n60470), .O(n19637[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_5 (.CI(n60470), .I0(n19856[2]), .I1(n332_adj_5363), 
            .CO(n60471));
    SB_LUT4 add_6550_4_lut (.I0(GND_net), .I1(n19856[1]), .I2(n259_adj_5364), 
            .I3(n60469), .O(n19637[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_4 (.CI(n60469), .I0(n19856[1]), .I1(n259_adj_5364), 
            .CO(n60470));
    SB_LUT4 add_6550_3_lut (.I0(GND_net), .I1(n19856[0]), .I2(n186_adj_5365), 
            .I3(n60468), .O(n19637[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_3 (.CI(n60468), .I0(n19856[0]), .I1(n186_adj_5365), 
            .CO(n60469));
    SB_LUT4 add_6550_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19637[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11882_bdd_4_lut_63408 (.I0(n11882), .I1(n75261), .I2(setpoint[8]), 
            .I3(n4736), .O(n79294));
    defparam n11882_bdd_4_lut_63408.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_add_1221_6_lut (.I0(GND_net), .I1(n12381[3]), .I2(n366_adj_5366), 
            .I3(n59625), .O(n360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n60468));
    SB_LUT4 add_6346_19_lut (.I0(GND_net), .I1(n17006[16]), .I2(GND_net), 
            .I3(n60467), .O(n16362[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i31_2_lut (.I0(n455[15]), .I1(n48[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5368));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6346_18_lut (.I0(GND_net), .I1(n17006[15]), .I2(GND_net), 
            .I3(n60466), .O(n16362[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_18 (.CI(n60466), .I0(n17006[15]), .I1(GND_net), 
            .CO(n60467));
    SB_LUT4 add_6346_17_lut (.I0(GND_net), .I1(n17006[14]), .I2(GND_net), 
            .I3(n60465), .O(n16362[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i33_2_lut (.I0(n455[16]), .I1(n48[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5369));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6346_17 (.CI(n60465), .I0(n17006[14]), .I1(GND_net), 
            .CO(n60466));
    SB_LUT4 i59888_4_lut (.I0(n27_adj_5355), .I1(n15_adj_5352), .I2(n13_adj_5351), 
            .I3(n11_adj_5350), .O(n75744));
    defparam i59888_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6346_16_lut (.I0(GND_net), .I1(n17006[13]), .I2(n1111), 
            .I3(n60464), .O(n16362[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_16 (.CI(n60464), .I0(n17006[13]), .I1(n1111), .CO(n60465));
    SB_LUT4 add_6346_15_lut (.I0(GND_net), .I1(n17006[12]), .I2(n1038), 
            .I3(n60463), .O(n16362[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_6 (.CI(n59625), .I0(n12381[3]), .I1(n366_adj_5366), 
            .CO(n59626));
    SB_LUT4 mult_23_add_1221_5_lut (.I0(GND_net), .I1(n12381[2]), .I2(n293_adj_5370), 
            .I3(n59624), .O(n360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_15 (.CI(n60463), .I0(n17006[12]), .I1(n1038), .CO(n60464));
    SB_LUT4 add_6346_14_lut (.I0(GND_net), .I1(n17006[11]), .I2(n965), 
            .I3(n60462), .O(n16362[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_14 (.CI(n60462), .I0(n17006[11]), .I1(n965), .CO(n60463));
    SB_LUT4 add_6346_13_lut (.I0(GND_net), .I1(n17006[10]), .I2(n892), 
            .I3(n60461), .O(n16362[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_13 (.CI(n60461), .I0(n17006[10]), .I1(n892), .CO(n60462));
    SB_LUT4 add_6346_12_lut (.I0(GND_net), .I1(n17006[9]), .I2(n819), 
            .I3(n60460), .O(n16362[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_12 (.CI(n60460), .I0(n17006[9]), .I1(n819), .CO(n60461));
    SB_LUT4 add_6346_11_lut (.I0(GND_net), .I1(n17006[8]), .I2(n746), 
            .I3(n60459), .O(n16362[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_11 (.CI(n60459), .I0(n17006[8]), .I1(n746), .CO(n60460));
    SB_LUT4 add_6346_10_lut (.I0(GND_net), .I1(n17006[7]), .I2(n673), 
            .I3(n60458), .O(n16362[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_10 (.CI(n60458), .I0(n17006[7]), .I1(n673), .CO(n60459));
    SB_LUT4 add_6346_9_lut (.I0(GND_net), .I1(n17006[6]), .I2(n600), .I3(n60457), 
            .O(n16362[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_9 (.CI(n60457), .I0(n17006[6]), .I1(n600), .CO(n60458));
    SB_LUT4 add_6346_8_lut (.I0(GND_net), .I1(n17006[5]), .I2(n527), .I3(n60456), 
            .O(n16362[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_8 (.CI(n60456), .I0(n17006[5]), .I1(n527), .CO(n60457));
    SB_LUT4 add_6346_7_lut (.I0(GND_net), .I1(n17006[4]), .I2(n454), .I3(n60455), 
            .O(n16362[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_7 (.CI(n60455), .I0(n17006[4]), .I1(n454), .CO(n60456));
    SB_LUT4 add_6346_6_lut (.I0(GND_net), .I1(n17006[3]), .I2(n381), .I3(n60454), 
            .O(n16362[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_6 (.CI(n60454), .I0(n17006[3]), .I1(n381), .CO(n60455));
    SB_LUT4 add_6346_5_lut (.I0(GND_net), .I1(n17006[2]), .I2(n308_adj_5371), 
            .I3(n60453), .O(n16362[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_5 (.CI(n60453), .I0(n17006[2]), .I1(n308_adj_5371), 
            .CO(n60454));
    SB_LUT4 add_6346_4_lut (.I0(GND_net), .I1(n17006[1]), .I2(n235_adj_5372), 
            .I3(n60452), .O(n16362[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_4 (.CI(n60452), .I0(n17006[1]), .I1(n235_adj_5372), 
            .CO(n60453));
    SB_LUT4 add_6346_3_lut (.I0(GND_net), .I1(n17006[0]), .I2(n162), .I3(n60451), 
            .O(n16362[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60887_4_lut (.I0(n9_adj_5349), .I1(n7_adj_5347), .I2(n455[2]), 
            .I3(n48[2]), .O(n76743));
    defparam i60887_4_lut.LUT_INIT = 16'heffe;
    SB_CARRY add_6346_3 (.CI(n60451), .I0(n17006[0]), .I1(n162), .CO(n60452));
    SB_DFFSR counter_2045_2046__i1 (.Q(counter[0]), .C(clk16MHz), .D(n61[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 i61443_4_lut (.I0(n15_adj_5352), .I1(n13_adj_5351), .I2(n11_adj_5350), 
            .I3(n76743), .O(n77299));
    defparam i61443_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61437_4_lut (.I0(n21_adj_5346), .I1(n19_adj_5345), .I2(n17_adj_5343), 
            .I3(n77299), .O(n77293));
    defparam i61437_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_6346_2_lut (.I0(GND_net), .I1(n20_adj_5373), .I2(n89), 
            .I3(GND_net), .O(n16362[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_2045_2046__i14 (.Q(counter[13]), .C(clk16MHz), .D(n61[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i13 (.Q(counter[12]), .C(clk16MHz), .D(n61[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i12 (.Q(counter[11]), .C(clk16MHz), .D(n61[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i11 (.Q(counter[10]), .C(clk16MHz), .D(n61[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i10 (.Q(counter[9]), .C(clk16MHz), .D(n61[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i9 (.Q(counter[8]), .C(clk16MHz), .D(n61[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i8 (.Q(counter[7]), .C(clk16MHz), .D(n61[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i7 (.Q(counter[6]), .C(clk16MHz), .D(n61[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i6 (.Q(counter[5]), .C(clk16MHz), .D(n61[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i5 (.Q(counter[4]), .C(clk16MHz), .D(n61[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i4 (.Q(counter[3]), .C(clk16MHz), .D(n61[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i3 (.Q(counter[2]), .C(clk16MHz), .D(n61[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i2 (.Q(counter[1]), .C(clk16MHz), .D(n61[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 i59890_4_lut (.I0(n27_adj_5355), .I1(n25_adj_5340), .I2(n23_adj_5336), 
            .I3(n77293), .O(n75746));
    defparam i59890_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_28_i12_3_lut (.I0(n48[7]), .I1(n48[16]), .I2(n33_adj_5369), 
            .I3(GND_net), .O(n12_adj_5374));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6346_2 (.CI(GND_net), .I0(n20_adj_5373), .I1(n89), .CO(n60451));
    SB_LUT4 LessThan_28_i4_3_lut (.I0(n75139), .I1(n48[1]), .I2(n455[1]), 
            .I3(GND_net), .O(n4_adj_5375));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY mult_23_add_1221_5 (.CI(n59624), .I0(n12381[2]), .I1(n293_adj_5370), 
            .CO(n59625));
    SB_LUT4 i61433_3_lut (.I0(n4_adj_5375), .I1(n48[13]), .I2(n27_adj_5355), 
            .I3(GND_net), .O(n77289));   // verilog/motorControl.v(62[35:55])
    defparam i61433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6380_18_lut (.I0(GND_net), .I1(n17580[15]), .I2(GND_net), 
            .I3(n60450), .O(n17006[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61434_3_lut (.I0(n77289), .I1(n48[14]), .I2(n29_adj_5362), 
            .I3(GND_net), .O(n77290));   // verilog/motorControl.v(62[35:55])
    defparam i61434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6380_17_lut (.I0(GND_net), .I1(n17580[14]), .I2(GND_net), 
            .I3(n60449), .O(n17006[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_4_lut (.I0(GND_net), .I1(n12381[1]), .I2(n220_adj_5376), 
            .I3(n59623), .O(n360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_17 (.CI(n60449), .I0(n17580[14]), .I1(GND_net), 
            .CO(n60450));
    SB_LUT4 add_6380_16_lut (.I0(GND_net), .I1(n17580[13]), .I2(n1114), 
            .I3(n60448), .O(n17006[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_16 (.CI(n60448), .I0(n17580[13]), .I1(n1114), .CO(n60449));
    SB_LUT4 LessThan_28_i10_3_lut (.I0(n48[5]), .I1(n48[6]), .I2(n13_adj_5351), 
            .I3(GND_net), .O(n10_adj_5377));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6380_15_lut (.I0(GND_net), .I1(n17580[12]), .I2(n1041), 
            .I3(n60447), .O(n17006[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_15 (.CI(n60447), .I0(n17580[12]), .I1(n1041), .CO(n60448));
    SB_LUT4 add_6380_14_lut (.I0(GND_net), .I1(n17580[11]), .I2(n968), 
            .I3(n60446), .O(n17006[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_14 (.CI(n60446), .I0(n17580[11]), .I1(n968), .CO(n60447));
    SB_LUT4 add_6380_13_lut (.I0(GND_net), .I1(n17580[10]), .I2(n895), 
            .I3(n60445), .O(n17006[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i30_3_lut (.I0(n12_adj_5374), .I1(n48[17]), .I2(n35_adj_5358), 
            .I3(GND_net), .O(n30_adj_5378));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6380_13 (.CI(n60445), .I0(n17580[10]), .I1(n895), .CO(n60446));
    SB_LUT4 add_6380_12_lut (.I0(GND_net), .I1(n17580[9]), .I2(n822), 
            .I3(n60444), .O(n17006[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_12 (.CI(n60444), .I0(n17580[9]), .I1(n822), .CO(n60445));
    SB_CARRY mult_23_add_1221_4 (.CI(n59623), .I0(n12381[1]), .I1(n220_adj_5376), 
            .CO(n59624));
    SB_LUT4 i59882_4_lut (.I0(n33_adj_5369), .I1(n31_adj_5368), .I2(n29_adj_5362), 
            .I3(n75744), .O(n75738));
    defparam i59882_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61707_4_lut (.I0(n30_adj_5378), .I1(n10_adj_5377), .I2(n35_adj_5358), 
            .I3(n75735), .O(n77563));   // verilog/motorControl.v(62[35:55])
    defparam i61707_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_6380_11_lut (.I0(GND_net), .I1(n17580[8]), .I2(n749), 
            .I3(n60443), .O(n17006[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n207[12]), .I3(n58938), .O(n233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_11 (.CI(n60443), .I0(n17580[8]), .I1(n749), .CO(n60444));
    SB_LUT4 add_6380_10_lut (.I0(GND_net), .I1(n17580[7]), .I2(n676), 
            .I3(n60442), .O(n17006[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_10 (.CI(n60442), .I0(n17580[7]), .I1(n676), .CO(n60443));
    SB_LUT4 i60639_3_lut (.I0(n77290), .I1(n48[15]), .I2(n31_adj_5368), 
            .I3(GND_net), .O(n76495));   // verilog/motorControl.v(62[35:55])
    defparam i60639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6380_9_lut (.I0(GND_net), .I1(n17580[6]), .I2(n603), .I3(n60441), 
            .O(n17006[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_9 (.CI(n60441), .I0(n17580[6]), .I1(n603), .CO(n60442));
    SB_LUT4 mult_23_add_1221_3_lut (.I0(GND_net), .I1(n12381[0]), .I2(n147_adj_5379), 
            .I3(n59622), .O(n360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_3 (.CI(n59622), .I0(n12381[0]), .I1(n147_adj_5379), 
            .CO(n59623));
    SB_LUT4 mult_23_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_5380), .I2(n74_adj_5381), 
            .I3(GND_net), .O(n360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6380_8_lut (.I0(GND_net), .I1(n17580[5]), .I2(n530), .I3(n60440), 
            .O(n17006[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i8_3_lut (.I0(n48[4]), .I1(n48[8]), .I2(n17_adj_5343), 
            .I3(GND_net), .O(n8_adj_5382));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i6_3_lut (.I0(n48[2]), .I1(n48[3]), .I2(n7_adj_5347), 
            .I3(GND_net), .O(n6_adj_5383));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i16_3_lut (.I0(n8_adj_5382), .I1(n48[9]), .I2(n19_adj_5345), 
            .I3(GND_net), .O(n16_adj_5384));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62026_4_lut (.I0(n16_adj_5384), .I1(n6_adj_5383), .I2(n19_adj_5345), 
            .I3(n75760), .O(n77882));   // verilog/motorControl.v(62[35:55])
    defparam i62026_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62027_3_lut (.I0(n77882), .I1(n48[10]), .I2(n21_adj_5346), 
            .I3(GND_net), .O(n77883));   // verilog/motorControl.v(62[35:55])
    defparam i62027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61850_3_lut (.I0(n77883), .I1(n48[11]), .I2(n23_adj_5336), 
            .I3(GND_net), .O(n77706));   // verilog/motorControl.v(62[35:55])
    defparam i61850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61843_4_lut (.I0(n33_adj_5369), .I1(n31_adj_5368), .I2(n29_adj_5362), 
            .I3(n75746), .O(n77699));
    defparam i61843_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62194_4_lut (.I0(n76495), .I1(n77563), .I2(n35_adj_5358), 
            .I3(n75738), .O(n78050));   // verilog/motorControl.v(62[35:55])
    defparam i62194_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60637_3_lut (.I0(n77706), .I1(n48[12]), .I2(n25_adj_5340), 
            .I3(GND_net), .O(n76493));   // verilog/motorControl.v(62[35:55])
    defparam i60637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62196_4_lut (.I0(n76493), .I1(n78050), .I2(n35_adj_5358), 
            .I3(n77699), .O(n78052));   // verilog/motorControl.v(62[35:55])
    defparam i62196_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_28_i38_3_lut (.I0(n78052), .I1(n48[18]), .I2(n461), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_6380_8 (.CI(n60440), .I0(n17580[5]), .I1(n530), .CO(n60441));
    SB_LUT4 LessThan_28_i42_3_lut (.I0(n48[20]), .I1(n48[21]), .I2(n455[21]), 
            .I3(GND_net), .O(n42));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59874_4_lut (.I0(n455[21]), .I1(n455[20]), .I2(n48[21]), 
            .I3(n48[20]), .O(n75730));
    defparam i59874_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_28_i45_rep_153_2_lut (.I0(n455[22]), .I1(n48[22]), 
            .I2(GND_net), .I3(GND_net), .O(n79794));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i45_rep_153_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_23_add_1221_2 (.CI(GND_net), .I0(n5_adj_5380), .I1(n74_adj_5381), 
            .CO(n59622));
    SB_LUT4 LessThan_28_i44_3_lut (.I0(n42), .I1(n48[22]), .I2(n455[22]), 
            .I3(GND_net), .O(n44_adj_5387));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i44_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61709_4_lut (.I0(n44_adj_5387), .I1(n40), .I2(n79794), .I3(n75730), 
            .O(n77565));   // verilog/motorControl.v(62[35:55])
    defparam i61709_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_6380_7_lut (.I0(GND_net), .I1(n17580[4]), .I2(n457_adj_5388), 
            .I3(n60439), .O(n17006[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6562_11_lut (.I0(GND_net), .I1(n19974[8]), .I2(n770_adj_5389), 
            .I3(n59621), .O(n19778[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_7 (.CI(n60439), .I0(n17580[4]), .I1(n457_adj_5388), 
            .CO(n60440));
    SB_LUT4 add_6562_10_lut (.I0(GND_net), .I1(n19974[7]), .I2(n697_adj_5390), 
            .I3(n59620), .O(n19778[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6380_6_lut (.I0(GND_net), .I1(n17580[3]), .I2(n384_adj_5391), 
            .I3(n60438), .O(n17006[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_6 (.CI(n60438), .I0(n17580[3]), .I1(n384_adj_5391), 
            .CO(n60439));
    SB_LUT4 add_6380_5_lut (.I0(GND_net), .I1(n17580[2]), .I2(n311_adj_5392), 
            .I3(n60437), .O(n17006[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_10 (.CI(n59620), .I0(n19974[7]), .I1(n697_adj_5390), 
            .CO(n59621));
    SB_LUT4 LessThan_26_i40_3_lut (.I0(n38_adj_29), .I1(n455[20]), .I2(n41_adj_5335), 
            .I3(GND_net), .O(n40_adj_5394));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62215_4_lut (.I0(n40_adj_5394), .I1(n36), .I2(n41_adj_5335), 
            .I3(n75815), .O(n78071));   // verilog/motorControl.v(62[14:31])
    defparam i62215_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_6562_9_lut (.I0(GND_net), .I1(n19974[6]), .I2(n624_adj_5395), 
            .I3(n59619), .O(n19778[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_5 (.CI(n60437), .I0(n17580[2]), .I1(n311_adj_5392), 
            .CO(n60438));
    SB_LUT4 add_6380_4_lut (.I0(GND_net), .I1(n17580[1]), .I2(n238_adj_5396), 
            .I3(n60436), .O(n17006[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62216_3_lut (.I0(n78071), .I1(n455[21]), .I2(deadband[21]), 
            .I3(GND_net), .O(n78072));   // verilog/motorControl.v(62[14:31])
    defparam i62216_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_6380_4 (.CI(n60436), .I0(n17580[1]), .I1(n238_adj_5396), 
            .CO(n60437));
    SB_LUT4 i61710_3_lut (.I0(n77565), .I1(n455[23]), .I2(n47), .I3(GND_net), 
            .O(n77566));   // verilog/motorControl.v(62[35:55])
    defparam i61710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62079_3_lut (.I0(n78072), .I1(n455[22]), .I2(deadband[22]), 
            .I3(GND_net), .O(n77935));   // verilog/motorControl.v(62[14:31])
    defparam i62079_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30637_4_lut (.I0(n77935), .I1(n77566), .I2(deadband[23]), 
            .I3(n455[23]), .O(n44726));
    defparam i30637_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 mult_23_i65_2_lut (.I0(\Kp[1] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i18_2_lut (.I0(\Kp[0] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_5398));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6562_9 (.CI(n59619), .I0(n19974[6]), .I1(n624_adj_5395), 
            .CO(n59620));
    SB_LUT4 add_6380_3_lut (.I0(GND_net), .I1(n17580[0]), .I2(n165), .I3(n60435), 
            .O(n17006[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_3 (.CI(n60435), .I0(n17580[0]), .I1(n165), .CO(n60436));
    SB_LUT4 n79294_bdd_4_lut (.I0(n79294), .I1(n535[8]), .I2(n455[8]), 
            .I3(n4736), .O(n79297));
    defparam n79294_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_6380_2_lut (.I0(GND_net), .I1(n23_adj_5399), .I2(n92), 
            .I3(GND_net), .O(n17006[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11882_bdd_4_lut_63403 (.I0(n11882), .I1(n75260), .I2(setpoint[7]), 
            .I3(n4736), .O(n79288));
    defparam n11882_bdd_4_lut_63403.LUT_INIT = 16'he4aa;
    SB_LUT4 n79288_bdd_4_lut (.I0(n79288), .I1(n535[7]), .I2(n455[7]), 
            .I3(n4736), .O(n79291));
    defparam n79288_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_6562_8_lut (.I0(GND_net), .I1(n19974[5]), .I2(n551_adj_5245), 
            .I3(n59618), .O(n19778[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_8 (.CI(n59618), .I0(n19974[5]), .I1(n551_adj_5245), 
            .CO(n59619));
    SB_LUT4 mult_23_i114_2_lut (.I0(\Kp[2] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6562_7_lut (.I0(GND_net), .I1(n19974[4]), .I2(n478_adj_5234), 
            .I3(n59617), .O(n19778[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_2 (.CI(GND_net), .I0(n23_adj_5399), .I1(n92), .CO(n60435));
    SB_LUT4 add_6569_10_lut (.I0(GND_net), .I1(n20035[7]), .I2(n700), 
            .I3(n60434), .O(n19856[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11882_bdd_4_lut_63398 (.I0(n11882), .I1(n75259), .I2(setpoint[6]), 
            .I3(n4736), .O(n79282));
    defparam n11882_bdd_4_lut_63398.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i163_2_lut (.I0(\Kp[3] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_5400));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i212_2_lut (.I0(\Kp[4] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_5401));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i261_2_lut (.I0(\Kp[5] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_5402));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[7]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51961_2_lut (.I0(n25921), .I1(n44726), .I2(GND_net), .I3(GND_net), 
            .O(n67768));
    defparam i51961_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_6569_9_lut (.I0(GND_net), .I1(n20035[6]), .I2(n627), .I3(n60433), 
            .O(n19856[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_7 (.CI(n59617), .I0(n19974[4]), .I1(n478_adj_5234), 
            .CO(n59618));
    SB_LUT4 mult_23_i310_2_lut (.I0(\Kp[6] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_5404));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i359_2_lut (.I0(\Kp[7] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[8]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i408_2_lut (.I0(\Kp[8] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(n131), .I1(n5076), .I2(n67768), .I3(n24_adj_30), 
            .O(n4736));
    defparam i3_4_lut.LUT_INIT = 16'hcfdf;
    SB_CARRY add_6569_9 (.CI(n60433), .I0(n20035[6]), .I1(n627), .CO(n60434));
    SB_LUT4 i59836_2_lut (.I0(PWMLimit[15]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75285));
    defparam i59836_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[9]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i59768_4_lut (.I0(n27_adj_5297), .I1(n15_adj_5295), .I2(n13_adj_5293), 
            .I3(n11_adj_5290), .O(n75624));
    defparam i59768_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i457_2_lut (.I0(\Kp[9] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_5289), 
            .I3(GND_net), .O(n12_adj_5408));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_5293), 
            .I3(GND_net), .O(n10_adj_5409));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i85_2_lut (.I0(\Kp[1] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_5410));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6562_6_lut (.I0(GND_net), .I1(n19974[3]), .I2(n405), .I3(n59616), 
            .O(n19778[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i38_2_lut (.I0(\Kp[0] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_5411));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i30_3_lut (.I0(n12_adj_5408), .I1(n535[17]), .I2(n35_adj_5207), 
            .I3(GND_net), .O(n30_adj_5412));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6569_8_lut (.I0(GND_net), .I1(n20035[5]), .I2(n554), .I3(n60432), 
            .O(n19856[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_8 (.CI(n60432), .I0(n20035[5]), .I1(n554), .CO(n60433));
    SB_LUT4 mult_23_i506_2_lut (.I0(\Kp[10] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6562_6 (.CI(n59616), .I0(n19974[3]), .I1(n405), .CO(n59617));
    SB_LUT4 i60720_4_lut (.I0(n13_adj_5293), .I1(n11_adj_5290), .I2(n9_adj_5203), 
            .I3(n75664), .O(n76576));
    defparam i60720_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_6569_7_lut (.I0(GND_net), .I1(n20035[4]), .I2(n481), .I3(n60431), 
            .O(n19856[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6562_5_lut (.I0(GND_net), .I1(n19974[2]), .I2(n332_adj_5139), 
            .I3(n59615), .O(n19778[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_5 (.CI(n59615), .I0(n19974[2]), .I1(n332_adj_5139), 
            .CO(n59616));
    SB_LUT4 add_6562_4_lut (.I0(GND_net), .I1(n19974[1]), .I2(n259), .I3(n59614), 
            .O(n19778[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_4 (.CI(n59614), .I0(n19974[1]), .I1(n259), .CO(n59615));
    SB_LUT4 add_6562_3_lut (.I0(GND_net), .I1(n19974[0]), .I2(n186), .I3(n59613), 
            .O(n19778[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_3 (.CI(n59613), .I0(n19974[0]), .I1(n186), .CO(n59614));
    SB_LUT4 mult_23_i555_2_lut (.I0(\Kp[11] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60716_4_lut (.I0(n19_adj_5196), .I1(n17_adj_5195), .I2(n15_adj_5295), 
            .I3(n76576), .O(n76572));
    defparam i60716_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_6569_7 (.CI(n60431), .I0(n20035[4]), .I1(n481), .CO(n60432));
    SB_LUT4 add_6569_6_lut (.I0(GND_net), .I1(n20035[3]), .I2(n408), .I3(n60430), 
            .O(n19856[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_6 (.CI(n60430), .I0(n20035[3]), .I1(n408), .CO(n60431));
    SB_LUT4 add_6569_5_lut (.I0(GND_net), .I1(n20035[2]), .I2(n335), .I3(n60429), 
            .O(n19856[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i604_2_lut (.I0(\Kp[12] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6569_5 (.CI(n60429), .I0(n20035[2]), .I1(n335), .CO(n60430));
    SB_LUT4 mult_23_i134_2_lut (.I0(\Kp[2] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_5413));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i62022_4_lut (.I0(n25_adj_5201), .I1(n23_adj_5200), .I2(n21_adj_5198), 
            .I3(n76572), .O(n77878));
    defparam i62022_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[10]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6569_4_lut (.I0(GND_net), .I1(n20035[1]), .I2(n262), .I3(n60428), 
            .O(n19856[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i183_2_lut (.I0(\Kp[3] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_5415));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6562_2_lut (.I0(GND_net), .I1(n44_adj_5416), .I2(n113_adj_5417), 
            .I3(GND_net), .O(n19778[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_2 (.CI(GND_net), .I0(n44_adj_5416), .I1(n113_adj_5417), 
            .CO(n59613));
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n30516), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n30515), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n30514), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n30513), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n30512), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n30511), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n30510), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_6569_4 (.CI(n60428), .I0(n20035[1]), .I1(n262), .CO(n60429));
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n30509), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n30508), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n207[23]), .I1(\Kp[2] ), .I2(n4_adj_5418), 
            .I3(n207[22]), .O(n71550));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'h6ca0;
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n30507), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n30505), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n30503), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n30502), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n30501), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n30500), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n30499), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6569_3_lut (.I0(GND_net), .I1(n20035[0]), .I2(n189), .I3(n60427), 
            .O(n19856[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n30498), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n30497), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n30496), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i61377_4_lut (.I0(n31_adj_5190), .I1(n29_adj_5189), .I2(n27_adj_5297), 
            .I3(n77878), .O(n77233));
    defparam i61377_4_lut.LUT_INIT = 16'hfeff;
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n30495), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n30490), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_6569_3 (.CI(n60427), .I0(n20035[0]), .I1(n189), .CO(n60428));
    SB_LUT4 mult_23_i232_2_lut (.I0(\Kp[4] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_5419));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i232_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n30489), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6569_2_lut (.I0(GND_net), .I1(n47_adj_5420), .I2(n116), 
            .I3(GND_net), .O(n19856[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n30481), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n207[22]), .I1(n20470[1]), .I2(n4_adj_5421), 
            .I3(\Kp[3] ), .O(n20372[2]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hc66c;
    SB_LUT4 mult_23_i281_2_lut (.I0(\Kp[5] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_5422));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i234_2_lut (.I0(\Kp[4] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347_adj_5423));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i234_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6569_2 (.CI(GND_net), .I0(n47_adj_5420), .I1(n116), .CO(n60427));
    SB_LUT4 add_6412_17_lut (.I0(GND_net), .I1(n18088[14]), .I2(GND_net), 
            .I3(n60426), .O(n17580[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1794 (.I0(n20470[1]), .I1(n6_adj_5424), .I2(n347_adj_5423), 
            .I3(n67007), .O(n20372[3]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_i653_2_lut (.I0(\Kp[13] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i702_2_lut (.I0(\Kp[14] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i62243_4_lut (.I0(n37_adj_5192), .I1(n35_adj_5207), .I2(n33_adj_5289), 
            .I3(n77233), .O(n78099));
    defparam i62243_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_6412_16_lut (.I0(GND_net), .I1(n18088[13]), .I2(n1117), 
            .I3(n60425), .O(n17580[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i751_2_lut (.I0(\Kp[15] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_5425));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_5191), 
            .I3(GND_net), .O(n16_adj_5426));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1795 (.I0(n71546), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5421));   // verilog/motorControl.v(61[20:26])
    defparam i1_2_lut_adj_1795.LUT_INIT = 16'h8888;
    SB_LUT4 i44643_4_lut (.I0(n20470[1]), .I1(\Kp[3] ), .I2(n4_adj_5421), 
            .I3(n207[22]), .O(n6_adj_5424));   // verilog/motorControl.v(61[20:26])
    defparam i44643_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_3_lut_adj_1796 (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n71546));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_adj_1796.LUT_INIT = 16'hc8c8;
    SB_LUT4 i56250_3_lut (.I0(n207[23]), .I1(n71546), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n67007));   // verilog/motorControl.v(61[20:26])
    defparam i56250_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i44774_3_lut (.I0(n207[23]), .I1(n58648), .I2(n69342), .I3(GND_net), 
            .O(n20470[1]));   // verilog/motorControl.v(61[20:26])
    defparam i44774_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_23_i40_2_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_5427));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1797 (.I0(\Kp[1] ), .I1(\Kp[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5418));
    defparam i1_2_lut_adj_1797.LUT_INIT = 16'h6666;
    SB_LUT4 i61425_3_lut (.I0(n6_adj_5428), .I1(n535[10]), .I2(n21_adj_5198), 
            .I3(GND_net), .O(n77281));   // verilog/motorControl.v(65[25:41])
    defparam i61425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i330_2_lut (.I0(\Kp[6] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_5429));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(n207[23]), .I1(\Kp[5] ), .I2(n69342), 
            .I3(n207[22]), .O(n71536));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hc60a;
    SB_LUT4 i1_rep_549_2_lut (.I0(n20470[1]), .I1(n67007), .I2(GND_net), 
            .I3(GND_net), .O(n80190));   // verilog/motorControl.v(61[20:26])
    defparam i1_rep_549_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n58648), .I1(n71536), .I2(\Kp[4] ), 
            .I3(n207[23]), .O(n71540));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'h9666;
    SB_LUT4 i44651_4_lut (.I0(n80190), .I1(\Kp[4] ), .I2(n6_adj_5424), 
            .I3(n207[22]), .O(n8_adj_5430));   // verilog/motorControl.v(61[20:26])
    defparam i44651_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i44604_4_lut (.I0(n20470[1]), .I1(\Kp[3] ), .I2(n71546), .I3(n207[23]), 
            .O(n6_adj_5431));   // verilog/motorControl.v(61[20:26])
    defparam i44604_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n6_adj_5431), .I1(n8_adj_5430), .I2(n71540), 
            .I3(n67007), .O(n69227));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'h6996;
    SB_CARRY add_6412_16 (.CI(n60425), .I0(n18088[13]), .I1(n1117), .CO(n60426));
    SB_LUT4 add_6412_15_lut (.I0(GND_net), .I1(n18088[12]), .I2(n1044_adj_5432), 
            .I3(n60424), .O(n17580[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_15 (.CI(n60424), .I0(n18088[12]), .I1(n1044_adj_5432), 
            .CO(n60425));
    SB_LUT4 add_6412_14_lut (.I0(GND_net), .I1(n18088[11]), .I2(n971_adj_5433), 
            .I3(n60423), .O(n17580[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_14 (.CI(n60423), .I0(n18088[11]), .I1(n971_adj_5433), 
            .CO(n60424));
    SB_LUT4 i61426_3_lut (.I0(n77281), .I1(n535[11]), .I2(n23_adj_5200), 
            .I3(GND_net), .O(n77282));   // verilog/motorControl.v(65[25:41])
    defparam i61426_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_16_10 (.CI(n58938), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n207[12]), .CO(n58939));
    SB_LUT4 i59774_4_lut (.I0(n21_adj_5198), .I1(n19_adj_5196), .I2(n17_adj_5195), 
            .I3(n9_adj_5203), .O(n75630));
    defparam i59774_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6412_13_lut (.I0(GND_net), .I1(n18088[10]), .I2(n898_adj_5434), 
            .I3(n60422), .O(n17580[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_13 (.CI(n60422), .I0(n18088[10]), .I1(n898_adj_5434), 
            .CO(n60423));
    SB_LUT4 add_6412_12_lut (.I0(GND_net), .I1(n18088[9]), .I2(n825_adj_5435), 
            .I3(n60421), .O(n17580[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_12 (.CI(n60421), .I0(n18088[9]), .I1(n825_adj_5435), 
            .CO(n60422));
    SB_LUT4 add_6412_11_lut (.I0(GND_net), .I1(n18088[8]), .I2(n752_adj_5436), 
            .I3(n60420), .O(n17580[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_11 (.CI(n60420), .I0(n18088[8]), .I1(n752_adj_5436), 
            .CO(n60421));
    SB_LUT4 add_6412_10_lut (.I0(GND_net), .I1(n18088[7]), .I2(n679_adj_5437), 
            .I3(n60419), .O(n17580[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_10 (.CI(n60419), .I0(n18088[7]), .I1(n679_adj_5437), 
            .CO(n60420));
    SB_LUT4 add_6412_9_lut (.I0(GND_net), .I1(n18088[6]), .I2(n606_adj_5438), 
            .I3(n60418), .O(n17580[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_9 (.CI(n60418), .I0(n18088[6]), .I1(n606_adj_5438), 
            .CO(n60419));
    SB_LUT4 add_6412_8_lut (.I0(GND_net), .I1(n18088[5]), .I2(n533_adj_5439), 
            .I3(n60417), .O(n17580[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_8 (.CI(n60417), .I0(n18088[5]), .I1(n533_adj_5439), 
            .CO(n60418));
    SB_LUT4 add_6412_7_lut (.I0(GND_net), .I1(n18088[4]), .I2(n460_adj_5440), 
            .I3(n60416), .O(n17580[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_7 (.CI(n60416), .I0(n18088[4]), .I1(n460_adj_5440), 
            .CO(n60417));
    SB_LUT4 add_6412_6_lut (.I0(GND_net), .I1(n18088[3]), .I2(n387_adj_5441), 
            .I3(n60415), .O(n17580[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_6 (.CI(n60415), .I0(n18088[3]), .I1(n387_adj_5441), 
            .CO(n60416));
    SB_LUT4 add_6412_5_lut (.I0(GND_net), .I1(n18088[2]), .I2(n314_adj_5442), 
            .I3(n60414), .O(n17580[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_5 (.CI(n60414), .I0(n18088[2]), .I1(n314_adj_5442), 
            .CO(n60415));
    SB_LUT4 add_6139_23_lut (.I0(GND_net), .I1(n13443[20]), .I2(GND_net), 
            .I3(n59590), .O(n12381[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6139_22_lut (.I0(GND_net), .I1(n13443[19]), .I2(GND_net), 
            .I3(n59589), .O(n12381[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_22 (.CI(n59589), .I0(n13443[19]), .I1(GND_net), 
            .CO(n59590));
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29775), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6139_21_lut (.I0(GND_net), .I1(n13443[18]), .I2(GND_net), 
            .I3(n59588), .O(n12381[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_21 (.CI(n59588), .I0(n13443[18]), .I1(GND_net), 
            .CO(n59589));
    SB_LUT4 add_6139_20_lut (.I0(GND_net), .I1(n13443[17]), .I2(GND_net), 
            .I3(n59587), .O(n12381[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_20 (.CI(n59587), .I0(n13443[17]), .I1(GND_net), 
            .CO(n59588));
    SB_LUT4 add_6139_19_lut (.I0(GND_net), .I1(n13443[16]), .I2(GND_net), 
            .I3(n59586), .O(n12381[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_19 (.CI(n59586), .I0(n13443[16]), .I1(GND_net), 
            .CO(n59587));
    SB_LUT4 add_6139_18_lut (.I0(GND_net), .I1(n13443[15]), .I2(GND_net), 
            .I3(n59585), .O(n12381[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n79249), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_32_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_5195), 
            .I3(GND_net), .O(n8_adj_5443));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6139_18 (.CI(n59585), .I0(n13443[15]), .I1(GND_net), 
            .CO(n59586));
    SB_LUT4 add_6139_17_lut (.I0(GND_net), .I1(n13443[14]), .I2(GND_net), 
            .I3(n59584), .O(n12381[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_17 (.CI(n59584), .I0(n13443[14]), .I1(GND_net), 
            .CO(n59585));
    SB_LUT4 add_6139_16_lut (.I0(GND_net), .I1(n13443[13]), .I2(n1099_adj_5444), 
            .I3(n59583), .O(n12381[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_16 (.CI(n59583), .I0(n13443[13]), .I1(n1099_adj_5444), 
            .CO(n59584));
    SB_LUT4 add_6139_15_lut (.I0(GND_net), .I1(n13443[12]), .I2(n1026_adj_5445), 
            .I3(n59582), .O(n12381[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_15 (.CI(n59582), .I0(n13443[12]), .I1(n1026_adj_5445), 
            .CO(n59583));
    SB_LUT4 add_6139_14_lut (.I0(GND_net), .I1(n13443[11]), .I2(n953_adj_5446), 
            .I3(n59581), .O(n12381[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_14 (.CI(n59581), .I0(n13443[11]), .I1(n953_adj_5446), 
            .CO(n59582));
    SB_LUT4 LessThan_32_i24_3_lut (.I0(n16_adj_5426), .I1(n535[22]), .I2(n45_adj_5187), 
            .I3(GND_net), .O(n24_adj_5447));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59734_4_lut (.I0(n43_adj_5191), .I1(n25_adj_5201), .I2(n23_adj_5200), 
            .I3(n75630), .O(n75590));
    defparam i59734_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61713_4_lut (.I0(n24_adj_5447), .I1(n8_adj_5443), .I2(n45_adj_5187), 
            .I3(n75576), .O(n77569));   // verilog/motorControl.v(65[25:41])
    defparam i61713_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60651_3_lut (.I0(n77282), .I1(n535[12]), .I2(n25_adj_5201), 
            .I3(GND_net), .O(n76507));   // verilog/motorControl.v(65[25:41])
    defparam i60651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6139_13_lut (.I0(GND_net), .I1(n13443[10]), .I2(n880_adj_5448), 
            .I3(n59580), .O(n12381[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i4_4_lut (.I0(n455[0]), .I1(n535[1]), .I2(n455[1]), 
            .I3(n535[0]), .O(n4_adj_5449));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_6139_13 (.CI(n59580), .I0(n13443[10]), .I1(n880_adj_5448), 
            .CO(n59581));
    SB_LUT4 add_6139_12_lut (.I0(GND_net), .I1(n13443[9]), .I2(n807_adj_5450), 
            .I3(n59579), .O(n12381[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_12 (.CI(n59579), .I0(n13443[9]), .I1(n807_adj_5450), 
            .CO(n59580));
    SB_LUT4 add_6139_11_lut (.I0(GND_net), .I1(n13443[8]), .I2(n734_adj_5451), 
            .I3(n59578), .O(n12381[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_11 (.CI(n59578), .I0(n13443[8]), .I1(n734_adj_5451), 
            .CO(n59579));
    SB_LUT4 add_6139_10_lut (.I0(GND_net), .I1(n13443[7]), .I2(n661_adj_5452), 
            .I3(n59577), .O(n12381[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_10 (.CI(n59577), .I0(n13443[7]), .I1(n661_adj_5452), 
            .CO(n59578));
    SB_LUT4 i61421_3_lut (.I0(n4_adj_5449), .I1(n535[13]), .I2(n27_adj_5297), 
            .I3(GND_net), .O(n77277));   // verilog/motorControl.v(65[25:41])
    defparam i61421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6139_9_lut (.I0(GND_net), .I1(n13443[6]), .I2(n588_adj_5453), 
            .I3(n59576), .O(n12381[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_9 (.CI(n59576), .I0(n13443[6]), .I1(n588_adj_5453), 
            .CO(n59577));
    SB_LUT4 add_6139_8_lut (.I0(GND_net), .I1(n13443[5]), .I2(n515_adj_5454), 
            .I3(n59575), .O(n12381[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61422_3_lut (.I0(n77277), .I1(n535[14]), .I2(n29_adj_5189), 
            .I3(GND_net), .O(n77278));   // verilog/motorControl.v(65[25:41])
    defparam i61422_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6139_8 (.CI(n59575), .I0(n13443[5]), .I1(n515_adj_5454), 
            .CO(n59576));
    SB_LUT4 add_6139_7_lut (.I0(GND_net), .I1(n13443[4]), .I2(n442_adj_5455), 
            .I3(n59574), .O(n12381[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_7 (.CI(n59574), .I0(n13443[4]), .I1(n442_adj_5455), 
            .CO(n59575));
    SB_LUT4 add_6139_6_lut (.I0(GND_net), .I1(n13443[3]), .I2(n369_adj_5456), 
            .I3(n59573), .O(n12381[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_6 (.CI(n59573), .I0(n13443[3]), .I1(n369_adj_5456), 
            .CO(n59574));
    SB_LUT4 add_6412_4_lut (.I0(GND_net), .I1(n18088[1]), .I2(n241_adj_5457), 
            .I3(n60413), .O(n17580[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6139_5_lut (.I0(GND_net), .I1(n13443[2]), .I2(n296_adj_5458), 
            .I3(n59572), .O(n12381[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_5 (.CI(n59572), .I0(n13443[2]), .I1(n296_adj_5458), 
            .CO(n59573));
    SB_LUT4 add_6139_4_lut (.I0(GND_net), .I1(n13443[1]), .I2(n223_adj_5459), 
            .I3(n59571), .O(n12381[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_4 (.CI(n60413), .I0(n18088[1]), .I1(n241_adj_5457), 
            .CO(n60414));
    SB_LUT4 i59757_4_lut (.I0(n33_adj_5289), .I1(n31_adj_5190), .I2(n29_adj_5189), 
            .I3(n75624), .O(n75613));
    defparam i59757_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62072_4_lut (.I0(n30_adj_5412), .I1(n10_adj_5409), .I2(n35_adj_5207), 
            .I3(n75609), .O(n77928));   // verilog/motorControl.v(65[25:41])
    defparam i62072_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60653_3_lut (.I0(n77278), .I1(n535[15]), .I2(n31_adj_5190), 
            .I3(GND_net), .O(n76509));   // verilog/motorControl.v(65[25:41])
    defparam i60653_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6139_4 (.CI(n59571), .I0(n13443[1]), .I1(n223_adj_5459), 
            .CO(n59572));
    SB_LUT4 add_6139_3_lut (.I0(GND_net), .I1(n13443[0]), .I2(n150_adj_5460), 
            .I3(n59570), .O(n12381[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_3 (.CI(n59570), .I0(n13443[0]), .I1(n150_adj_5460), 
            .CO(n59571));
    SB_LUT4 add_6139_2_lut (.I0(GND_net), .I1(n8_adj_5461), .I2(n77_adj_5462), 
            .I3(GND_net), .O(n12381[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6412_3_lut (.I0(GND_net), .I1(n18088[0]), .I2(n168_adj_5463), 
            .I3(n60412), .O(n17580[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_2 (.CI(GND_net), .I0(n8_adj_5461), .I1(n77_adj_5462), 
            .CO(n59570));
    SB_LUT4 add_6208_22_lut (.I0(GND_net), .I1(n14367[19]), .I2(GND_net), 
            .I3(n59569), .O(n13443[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_21_lut (.I0(GND_net), .I1(n14367[18]), .I2(GND_net), 
            .I3(n59568), .O(n13443[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_21 (.CI(n59568), .I0(n14367[18]), .I1(GND_net), 
            .CO(n59569));
    SB_CARRY add_6412_3 (.CI(n60412), .I0(n18088[0]), .I1(n168_adj_5463), 
            .CO(n60413));
    SB_LUT4 add_6208_20_lut (.I0(GND_net), .I1(n14367[17]), .I2(GND_net), 
            .I3(n59567), .O(n13443[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6506_13_lut (.I0(GND_net), .I1(n19374[10]), .I2(n910), 
            .I3(n59178), .O(n19063[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62289_4_lut (.I0(n76509), .I1(n77928), .I2(n35_adj_5207), 
            .I3(n75613), .O(n78145));   // verilog/motorControl.v(65[25:41])
    defparam i62289_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62290_3_lut (.I0(n78145), .I1(n535[18]), .I2(n37_adj_5192), 
            .I3(GND_net), .O(n78146));   // verilog/motorControl.v(65[25:41])
    defparam i62290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62261_3_lut (.I0(n78146), .I1(n535[19]), .I2(n39_adj_5186), 
            .I3(GND_net), .O(n78117));   // verilog/motorControl.v(65[25:41])
    defparam i62261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59737_4_lut (.I0(n43_adj_5191), .I1(n41_adj_5185), .I2(n39_adj_5186), 
            .I3(n78099), .O(n75593));
    defparam i59737_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6208_20 (.CI(n59567), .I0(n14367[17]), .I1(GND_net), 
            .CO(n59568));
    SB_LUT4 add_6208_19_lut (.I0(GND_net), .I1(n14367[16]), .I2(GND_net), 
            .I3(n59566), .O(n13443[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6506_12_lut (.I0(GND_net), .I1(n19374[9]), .I2(n837), 
            .I3(n59177), .O(n19063[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_12 (.CI(n59177), .I0(n19374[9]), .I1(n837), .CO(n59178));
    SB_CARRY add_6208_19 (.CI(n59566), .I0(n14367[16]), .I1(GND_net), 
            .CO(n59567));
    SB_LUT4 add_6208_18_lut (.I0(GND_net), .I1(n14367[15]), .I2(GND_net), 
            .I3(n59565), .O(n13443[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6506_11_lut (.I0(GND_net), .I1(n19374[8]), .I2(n764), 
            .I3(n59176), .O(n19063[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_11 (.CI(n59176), .I0(n19374[8]), .I1(n764), .CO(n59177));
    SB_CARRY add_6208_18 (.CI(n59565), .I0(n14367[15]), .I1(GND_net), 
            .CO(n59566));
    SB_LUT4 add_6208_17_lut (.I0(GND_net), .I1(n14367[14]), .I2(GND_net), 
            .I3(n59564), .O(n13443[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6506_10_lut (.I0(GND_net), .I1(n19374[7]), .I2(n691), 
            .I3(n59175), .O(n19063[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_10 (.CI(n59175), .I0(n19374[7]), .I1(n691), .CO(n59176));
    SB_CARRY add_6208_17 (.CI(n59564), .I0(n14367[14]), .I1(GND_net), 
            .CO(n59565));
    SB_LUT4 add_6208_16_lut (.I0(GND_net), .I1(n14367[13]), .I2(n1102_adj_5464), 
            .I3(n59563), .O(n13443[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6412_2_lut (.I0(GND_net), .I1(n26_adj_5465), .I2(n95_adj_5466), 
            .I3(GND_net), .O(n17580[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_16 (.CI(n59563), .I0(n14367[13]), .I1(n1102_adj_5464), 
            .CO(n59564));
    SB_LUT4 i61989_4_lut (.I0(n76507), .I1(n77569), .I2(n45_adj_5187), 
            .I3(n75590), .O(n77845));   // verilog/motorControl.v(65[25:41])
    defparam i61989_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60659_3_lut (.I0(n78117), .I1(n535[20]), .I2(n41_adj_5185), 
            .I3(GND_net), .O(n76515));   // verilog/motorControl.v(65[25:41])
    defparam i60659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62197_4_lut (.I0(n76515), .I1(n77845), .I2(n45_adj_5187), 
            .I3(n75593), .O(n78053));   // verilog/motorControl.v(65[25:41])
    defparam i62197_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2_4_lut_adj_1801 (.I0(n78053), .I1(n4_adj_5467), .I2(n455[23]), 
            .I3(n535[23]), .O(n69256));
    defparam i2_4_lut_adj_1801.LUT_INIT = 16'hdfcd;
    SB_LUT4 i6058_4_lut (.I0(n131), .I1(n4736), .I2(n24_adj_30), .I3(n69256), 
            .O(n11882));
    defparam i6058_4_lut.LUT_INIT = 16'h0737;
    SB_CARRY add_6412_2 (.CI(GND_net), .I0(n26_adj_5465), .I1(n95_adj_5466), 
            .CO(n60412));
    SB_LUT4 add_6208_15_lut (.I0(GND_net), .I1(n14367[12]), .I2(n1029_adj_5468), 
            .I3(n59562), .O(n13443[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_15 (.CI(n59562), .I0(n14367[12]), .I1(n1029_adj_5468), 
            .CO(n59563));
    SB_LUT4 add_6208_14_lut (.I0(GND_net), .I1(n14367[11]), .I2(n956_adj_5469), 
            .I3(n59561), .O(n13443[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6442_16_lut (.I0(GND_net), .I1(n18534[13]), .I2(n1120_adj_5470), 
            .I3(n60411), .O(n18088[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_14 (.CI(n59561), .I0(n14367[11]), .I1(n956_adj_5469), 
            .CO(n59562));
    SB_LUT4 add_6442_15_lut (.I0(GND_net), .I1(n18534[12]), .I2(n1047_adj_5471), 
            .I3(n60410), .O(n18088[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_13_lut (.I0(GND_net), .I1(n14367[10]), .I2(n883_adj_5472), 
            .I3(n59560), .O(n13443[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_13 (.CI(n59560), .I0(n14367[10]), .I1(n883_adj_5472), 
            .CO(n59561));
    SB_LUT4 add_6208_12_lut (.I0(GND_net), .I1(n14367[9]), .I2(n810_adj_5473), 
            .I3(n59559), .O(n13443[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6506_9_lut (.I0(GND_net), .I1(n19374[6]), .I2(n618), .I3(n59174), 
            .O(n19063[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_12 (.CI(n59559), .I0(n14367[9]), .I1(n810_adj_5473), 
            .CO(n59560));
    SB_LUT4 add_6208_11_lut (.I0(GND_net), .I1(n14367[8]), .I2(n737_adj_5474), 
            .I3(n59558), .O(n13443[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_9 (.CI(n59174), .I0(n19374[6]), .I1(n618), .CO(n59175));
    SB_LUT4 add_6506_8_lut (.I0(GND_net), .I1(n19374[5]), .I2(n545_adj_5475), 
            .I3(n59173), .O(n19063[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_11 (.CI(n59558), .I0(n14367[8]), .I1(n737_adj_5474), 
            .CO(n59559));
    SB_LUT4 add_6208_10_lut (.I0(GND_net), .I1(n14367[7]), .I2(n664_adj_5476), 
            .I3(n59557), .O(n13443[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_8 (.CI(n59173), .I0(n19374[5]), .I1(n545_adj_5475), 
            .CO(n59174));
    SB_LUT4 add_6506_7_lut (.I0(GND_net), .I1(n19374[4]), .I2(n472_adj_5477), 
            .I3(n59172), .O(n19063[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_10 (.CI(n59557), .I0(n14367[7]), .I1(n664_adj_5476), 
            .CO(n59558));
    SB_LUT4 add_6208_9_lut (.I0(GND_net), .I1(n14367[6]), .I2(n591_adj_5478), 
            .I3(n59556), .O(n13443[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_7 (.CI(n59172), .I0(n19374[4]), .I1(n472_adj_5477), 
            .CO(n59173));
    SB_LUT4 add_6506_6_lut (.I0(GND_net), .I1(n19374[3]), .I2(n399_adj_5479), 
            .I3(n59171), .O(n19063[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_9 (.CI(n59556), .I0(n14367[6]), .I1(n591_adj_5478), 
            .CO(n59557));
    SB_CARRY add_6442_15 (.CI(n60410), .I0(n18534[12]), .I1(n1047_adj_5471), 
            .CO(n60411));
    SB_LUT4 add_6442_14_lut (.I0(GND_net), .I1(n18534[11]), .I2(n974_adj_5480), 
            .I3(n60409), .O(n18088[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_14 (.CI(n60409), .I0(n18534[11]), .I1(n974_adj_5480), 
            .CO(n60410));
    SB_LUT4 add_6442_13_lut (.I0(GND_net), .I1(n18534[10]), .I2(n901_adj_5481), 
            .I3(n60408), .O(n18088[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_8_lut (.I0(GND_net), .I1(n14367[5]), .I2(n518_adj_5482), 
            .I3(n59555), .O(n13443[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_6 (.CI(n59171), .I0(n19374[3]), .I1(n399_adj_5479), 
            .CO(n59172));
    SB_LUT4 add_6506_5_lut (.I0(GND_net), .I1(n19374[2]), .I2(n326), .I3(n59170), 
            .O(n19063[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_8 (.CI(n59555), .I0(n14367[5]), .I1(n518_adj_5482), 
            .CO(n59556));
    SB_LUT4 add_6208_7_lut (.I0(GND_net), .I1(n14367[4]), .I2(n445_adj_5483), 
            .I3(n59554), .O(n13443[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_5 (.CI(n59170), .I0(n19374[2]), .I1(n326), .CO(n59171));
    SB_LUT4 add_6506_4_lut (.I0(GND_net), .I1(n19374[1]), .I2(n253_adj_5484), 
            .I3(n59169), .O(n19063[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_7 (.CI(n59554), .I0(n14367[4]), .I1(n445_adj_5483), 
            .CO(n59555));
    SB_LUT4 add_6208_6_lut (.I0(GND_net), .I1(n14367[3]), .I2(n372_adj_5485), 
            .I3(n59553), .O(n13443[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_4 (.CI(n59169), .I0(n19374[1]), .I1(n253_adj_5484), 
            .CO(n59170));
    SB_LUT4 add_6506_3_lut (.I0(GND_net), .I1(n19374[0]), .I2(n180), .I3(n59168), 
            .O(n19063[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_6 (.CI(n59553), .I0(n14367[3]), .I1(n372_adj_5485), 
            .CO(n59554));
    SB_LUT4 add_6208_5_lut (.I0(GND_net), .I1(n14367[2]), .I2(n299_adj_5486), 
            .I3(n59552), .O(n13443[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_3 (.CI(n59168), .I0(n19374[0]), .I1(n180), .CO(n59169));
    SB_LUT4 add_6506_2_lut (.I0(GND_net), .I1(n38_adj_5487), .I2(n107), 
            .I3(GND_net), .O(n19063[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_5 (.CI(n59552), .I0(n14367[2]), .I1(n299_adj_5486), 
            .CO(n59553));
    SB_LUT4 mult_24_i28_2_lut (.I0(\Ki[0] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5488));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i124_2_lut (.I0(\Ki[2] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_5490));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6208_4_lut (.I0(GND_net), .I1(n14367[1]), .I2(n226_adj_5491), 
            .I3(n59551), .O(n13443[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_4 (.CI(n59551), .I0(n14367[1]), .I1(n226_adj_5491), 
            .CO(n59552));
    SB_LUT4 add_6208_3_lut (.I0(GND_net), .I1(n14367[0]), .I2(n153_adj_5492), 
            .I3(n59550), .O(n13443[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_3 (.CI(n59550), .I0(n14367[0]), .I1(n153_adj_5492), 
            .CO(n59551));
    SB_LUT4 add_6208_2_lut (.I0(GND_net), .I1(n11_adj_5493), .I2(n80_adj_5494), 
            .I3(GND_net), .O(n13443[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_13 (.CI(n60408), .I0(n18534[10]), .I1(n901_adj_5481), 
            .CO(n60409));
    SB_CARRY add_6208_2 (.CI(GND_net), .I0(n11_adj_5493), .I1(n80_adj_5494), 
            .CO(n59550));
    SB_LUT4 add_6442_12_lut (.I0(GND_net), .I1(n18534[9]), .I2(n828_adj_5495), 
            .I3(n60407), .O(n18088[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_12 (.CI(n60407), .I0(n18534[9]), .I1(n828_adj_5495), 
            .CO(n60408));
    SB_LUT4 mult_24_i173_2_lut (.I0(\Ki[3] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_5496));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6506_2 (.CI(GND_net), .I0(n38_adj_5487), .I1(n107), .CO(n59168));
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[11]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6442_11_lut (.I0(GND_net), .I1(n18534[8]), .I2(n755_adj_5498), 
            .I3(n60406), .O(n18088[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[12]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6442_11 (.CI(n60406), .I0(n18534[8]), .I1(n755_adj_5498), 
            .CO(n60407));
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[13]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[14]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6442_10_lut (.I0(GND_net), .I1(n18534[7]), .I2(n682_adj_5502), 
            .I3(n60405), .O(n18088[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[15]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i222_2_lut (.I0(\Ki[4] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_5504));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[16]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i63_2_lut (.I0(\Kp[1] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_5506));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i16_2_lut (.I0(\Kp[0] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5507));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i112_2_lut (.I0(\Kp[2] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_5508));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_21_lut (.I0(GND_net), .I1(n15206[18]), .I2(GND_net), 
            .I3(n59528), .O(n14367[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_20_lut (.I0(GND_net), .I1(n15206[17]), .I2(GND_net), 
            .I3(n59527), .O(n14367[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[17]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6250_20 (.CI(n59527), .I0(n15206[17]), .I1(GND_net), 
            .CO(n59528));
    SB_LUT4 add_6250_19_lut (.I0(GND_net), .I1(n15206[16]), .I2(GND_net), 
            .I3(n59526), .O(n14367[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_19 (.CI(n59526), .I0(n15206[16]), .I1(GND_net), 
            .CO(n59527));
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[18]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6250_18_lut (.I0(GND_net), .I1(n15206[15]), .I2(GND_net), 
            .I3(n59525), .O(n14367[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i161_2_lut (.I0(\Kp[3] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_5511));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i161_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6250_18 (.CI(n59525), .I0(n15206[15]), .I1(GND_net), 
            .CO(n59526));
    SB_LUT4 add_6250_17_lut (.I0(GND_net), .I1(n15206[14]), .I2(GND_net), 
            .I3(n59524), .O(n14367[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_17 (.CI(n59524), .I0(n15206[14]), .I1(GND_net), 
            .CO(n59525));
    SB_LUT4 add_6250_16_lut (.I0(GND_net), .I1(n15206[13]), .I2(n1105_adj_5512), 
            .I3(n59523), .O(n14367[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_16 (.CI(n59523), .I0(n15206[13]), .I1(n1105_adj_5512), 
            .CO(n59524));
    SB_LUT4 add_6250_15_lut (.I0(GND_net), .I1(n15206[12]), .I2(n1032_adj_5513), 
            .I3(n59522), .O(n14367[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_15 (.CI(n59522), .I0(n15206[12]), .I1(n1032_adj_5513), 
            .CO(n59523));
    SB_LUT4 add_6250_14_lut (.I0(GND_net), .I1(n15206[11]), .I2(n959_adj_5514), 
            .I3(n59521), .O(n14367[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i71_2_lut (.I0(\Kp[1] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i24_2_lut (.I0(\Kp[0] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5148));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6250_14 (.CI(n59521), .I0(n15206[11]), .I1(n959_adj_5514), 
            .CO(n59522));
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[19]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6250_13_lut (.I0(GND_net), .I1(n15206[10]), .I2(n886_adj_5516), 
            .I3(n59520), .O(n14367[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_13 (.CI(n59520), .I0(n15206[10]), .I1(n886_adj_5516), 
            .CO(n59521));
    SB_LUT4 add_6250_12_lut (.I0(GND_net), .I1(n15206[9]), .I2(n813_adj_5517), 
            .I3(n59519), .O(n14367[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_12 (.CI(n59519), .I0(n15206[9]), .I1(n813_adj_5517), 
            .CO(n59520));
    SB_LUT4 add_6250_11_lut (.I0(GND_net), .I1(n15206[8]), .I2(n740_adj_5518), 
            .I3(n59518), .O(n14367[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i210_2_lut (.I0(\Kp[4] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_5519));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[20]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6250_11 (.CI(n59518), .I0(n15206[8]), .I1(n740_adj_5518), 
            .CO(n59519));
    SB_CARRY add_6442_10 (.CI(n60405), .I0(n18534[7]), .I1(n682_adj_5502), 
            .CO(n60406));
    SB_LUT4 add_6250_10_lut (.I0(GND_net), .I1(n15206[7]), .I2(n667_adj_5521), 
            .I3(n59517), .O(n14367[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_10 (.CI(n59517), .I0(n15206[7]), .I1(n667_adj_5521), 
            .CO(n59518));
    SB_LUT4 i30484_3_lut_4_lut (.I0(\control_mode[0] ), .I1(control_update), 
            .I2(n53108), .I3(\control_mode[1] ), .O(n28076));
    defparam i30484_3_lut_4_lut.LUT_INIT = 16'hc4cc;
    SB_LUT4 add_6250_9_lut (.I0(GND_net), .I1(n15206[6]), .I2(n594_adj_5522), 
            .I3(n59516), .O(n14367[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_9 (.CI(n59516), .I0(n15206[6]), .I1(n594_adj_5522), 
            .CO(n59517));
    SB_LUT4 add_6250_8_lut (.I0(GND_net), .I1(n15206[5]), .I2(n521_adj_5523), 
            .I3(n59515), .O(n14367[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_8 (.CI(n59515), .I0(n15206[5]), .I1(n521_adj_5523), 
            .CO(n59516));
    SB_LUT4 add_6250_7_lut (.I0(GND_net), .I1(n15206[4]), .I2(n448_adj_5524), 
            .I3(n59514), .O(n14367[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6442_9_lut (.I0(GND_net), .I1(n18534[6]), .I2(n609_adj_5525), 
            .I3(n60404), .O(n18088[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_9 (.CI(n60404), .I0(n18534[6]), .I1(n609_adj_5525), 
            .CO(n60405));
    SB_LUT4 add_6442_8_lut (.I0(GND_net), .I1(n18534[5]), .I2(n536_adj_5526), 
            .I3(n60403), .O(n18088[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_7 (.CI(n59514), .I0(n15206[4]), .I1(n448_adj_5524), 
            .CO(n59515));
    SB_LUT4 add_6250_6_lut (.I0(GND_net), .I1(n15206[3]), .I2(n375_adj_5527), 
            .I3(n59513), .O(n14367[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i259_2_lut (.I0(\Kp[5] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_5528));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i308_2_lut (.I0(\Kp[6] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_5529));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6250_6 (.CI(n59513), .I0(n15206[3]), .I1(n375_adj_5527), 
            .CO(n59514));
    SB_LUT4 add_6250_5_lut (.I0(GND_net), .I1(n15206[2]), .I2(n302_adj_5530), 
            .I3(n59512), .O(n14367[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i357_2_lut (.I0(\Kp[7] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_5531));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i357_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6250_5 (.CI(n59512), .I0(n15206[2]), .I1(n302_adj_5530), 
            .CO(n59513));
    SB_LUT4 add_6250_4_lut (.I0(GND_net), .I1(n15206[1]), .I2(n229_adj_5532), 
            .I3(n59511), .O(n14367[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_4 (.CI(n59511), .I0(n15206[1]), .I1(n229_adj_5532), 
            .CO(n59512));
    SB_LUT4 add_6250_3_lut (.I0(GND_net), .I1(n15206[0]), .I2(n156_adj_5533), 
            .I3(n59510), .O(n14367[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_3 (.CI(n59510), .I0(n15206[0]), .I1(n156_adj_5533), 
            .CO(n59511));
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[21]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6250_2_lut (.I0(GND_net), .I1(n14_adj_5535), .I2(n83_adj_5536), 
            .I3(GND_net), .O(n14367[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_2 (.CI(GND_net), .I0(n14_adj_5535), .I1(n83_adj_5536), 
            .CO(n59510));
    SB_CARRY add_6442_8 (.CI(n60403), .I0(n18534[5]), .I1(n536_adj_5526), 
            .CO(n60404));
    SB_LUT4 add_6442_7_lut (.I0(GND_net), .I1(n18534[4]), .I2(n463_adj_5537), 
            .I3(n60402), .O(n18088[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i271_2_lut (.I0(\Ki[5] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_5538));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i406_2_lut (.I0(\Kp[8] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_5539));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i455_2_lut (.I0(\Kp[9] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_5540));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i504_2_lut (.I0(\Kp[10] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_5541));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i553_2_lut (.I0(\Kp[11] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_5542));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i602_2_lut (.I0(\Kp[12] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_5543));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i602_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6442_7 (.CI(n60402), .I0(n18534[4]), .I1(n463_adj_5537), 
            .CO(n60403));
    SB_LUT4 mult_23_i651_2_lut (.I0(\Kp[13] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_5544));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6442_6_lut (.I0(GND_net), .I1(n18534[3]), .I2(n390_adj_5545), 
            .I3(n60401), .O(n18088[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_6 (.CI(n60401), .I0(n18534[3]), .I1(n390_adj_5545), 
            .CO(n60402));
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[22]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6442_5_lut (.I0(GND_net), .I1(n18534[2]), .I2(n317_adj_5547), 
            .I3(n60400), .O(n18088[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_5 (.CI(n60400), .I0(n18534[2]), .I1(n317_adj_5547), 
            .CO(n60401));
    SB_LUT4 mult_23_i700_2_lut (.I0(\Kp[14] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_5548));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5701[23]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i749_2_lut (.I0(\Kp[15] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_5550));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i320_2_lut (.I0(\Ki[6] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_5551));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6442_4_lut (.I0(GND_net), .I1(n18534[1]), .I2(n244_adj_5552), 
            .I3(n60399), .O(n18088[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_4 (.CI(n60399), .I0(n18534[1]), .I1(n244_adj_5552), 
            .CO(n60400));
    SB_LUT4 mult_24_i81_2_lut (.I0(\Ki[1] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i34_2_lut (.I0(\Ki[0] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6442_3_lut (.I0(GND_net), .I1(n18534[0]), .I2(n171_adj_5554), 
            .I3(n60398), .O(n18088[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_3 (.CI(n60398), .I0(n18534[0]), .I1(n171_adj_5554), 
            .CO(n60399));
    SB_LUT4 add_6442_2_lut (.I0(GND_net), .I1(n29_adj_5555), .I2(n98_adj_5556), 
            .I3(GND_net), .O(n18088[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_2 (.CI(GND_net), .I0(n29_adj_5555), .I1(n98_adj_5556), 
            .CO(n60398));
    SB_LUT4 mult_24_i130_2_lut (.I0(\Ki[2] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i179_2_lut (.I0(\Ki[3] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i228_2_lut (.I0(\Ki[4] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i369_2_lut (.I0(\Ki[7] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_5557));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[0]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6586_9_lut (.I0(GND_net), .I1(n20178[6]), .I2(n630), .I3(n60397), 
            .O(n20035[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6586_8_lut (.I0(GND_net), .I1(n20178[5]), .I2(n557), .I3(n60396), 
            .O(n20035[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_8 (.CI(n60396), .I0(n20178[5]), .I1(n557), .CO(n60397));
    SB_LUT4 mult_24_i277_2_lut (.I0(\Ki[5] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6586_7_lut (.I0(GND_net), .I1(n20178[4]), .I2(n484_adj_5559), 
            .I3(n60395), .O(n20035[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_7 (.CI(n60395), .I0(n20178[4]), .I1(n484_adj_5559), 
            .CO(n60396));
    SB_LUT4 mult_24_i326_2_lut (.I0(\Ki[6] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_5560));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i375_2_lut (.I0(\Ki[7] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_5561));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i424_2_lut (.I0(\Ki[8] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_5562));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6586_6_lut (.I0(GND_net), .I1(n20178[3]), .I2(n411_adj_5563), 
            .I3(n60394), .O(n20035[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i418_2_lut (.I0(\Ki[8] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_5564));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[1]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6586_6 (.CI(n60394), .I0(n20178[3]), .I1(n411_adj_5563), 
            .CO(n60395));
    SB_LUT4 unary_minus_33_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[2]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6586_5_lut (.I0(GND_net), .I1(n20178[2]), .I2(n338_adj_5567), 
            .I3(n60393), .O(n20035[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n79282_bdd_4_lut (.I0(n79282), .I1(n535[6]), .I2(n455[6]), 
            .I3(n4736), .O(n79285));
    defparam n79282_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_6586_5 (.CI(n60393), .I0(n20178[2]), .I1(n338_adj_5567), 
            .CO(n60394));
    SB_LUT4 mult_24_i467_2_lut (.I0(\Ki[9] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_5568));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6586_4_lut (.I0(GND_net), .I1(n20178[1]), .I2(n265_adj_5569), 
            .I3(n60392), .O(n20035[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_4 (.CI(n60392), .I0(n20178[1]), .I1(n265_adj_5569), 
            .CO(n60393));
    SB_LUT4 unary_minus_33_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[3]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6586_3_lut (.I0(GND_net), .I1(n20178[0]), .I2(n192_adj_5571), 
            .I3(n60391), .O(n20035[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_10_lut (.I0(GND_net), .I1(n20132[7]), .I2(n700_adj_5572), 
            .I3(n59489), .O(n19974[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_3 (.CI(n60391), .I0(n20178[0]), .I1(n192_adj_5571), 
            .CO(n60392));
    SB_LUT4 add_6586_2_lut (.I0(GND_net), .I1(n50_adj_5573), .I2(n119_adj_5574), 
            .I3(GND_net), .O(n20035[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_2 (.CI(GND_net), .I0(n50_adj_5573), .I1(n119_adj_5574), 
            .CO(n60391));
    SB_LUT4 add_6470_15_lut (.I0(GND_net), .I1(n18922[12]), .I2(n1050_adj_5575), 
            .I3(n60390), .O(n18534[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_9_lut (.I0(GND_net), .I1(n20132[6]), .I2(n627_adj_5576), 
            .I3(n59488), .O(n19974[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_9 (.CI(n59488), .I0(n20132[6]), .I1(n627_adj_5576), 
            .CO(n59489));
    SB_LUT4 add_6470_14_lut (.I0(GND_net), .I1(n18922[11]), .I2(n977_adj_5577), 
            .I3(n60389), .O(n18534[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_8_lut (.I0(GND_net), .I1(n20132[5]), .I2(n554_adj_5578), 
            .I3(n59487), .O(n19974[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_8 (.CI(n59487), .I0(n20132[5]), .I1(n554_adj_5578), 
            .CO(n59488));
    SB_LUT4 add_6580_7_lut (.I0(GND_net), .I1(n20132[4]), .I2(n481_adj_5579), 
            .I3(n59486), .O(n19974[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[4]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6470_14 (.CI(n60389), .I0(n18922[11]), .I1(n977_adj_5577), 
            .CO(n60390));
    SB_CARRY add_6580_7 (.CI(n59486), .I0(n20132[4]), .I1(n481_adj_5579), 
            .CO(n59487));
    SB_LUT4 unary_minus_33_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[5]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i516_2_lut (.I0(\Ki[10] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_5582));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6470_13_lut (.I0(GND_net), .I1(n18922[10]), .I2(n904_adj_5583), 
            .I3(n60388), .O(n18534[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_6_lut (.I0(GND_net), .I1(n20132[3]), .I2(n408_adj_5584), 
            .I3(n59485), .O(n19974[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[6]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6470_13 (.CI(n60388), .I0(n18922[10]), .I1(n904_adj_5583), 
            .CO(n60389));
    SB_LUT4 unary_minus_33_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[7]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_16_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n207[11]), .I3(n58937), .O(n233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_6 (.CI(n59485), .I0(n20132[3]), .I1(n408_adj_5584), 
            .CO(n59486));
    SB_LUT4 add_6580_5_lut (.I0(GND_net), .I1(n20132[2]), .I2(n335_adj_5587), 
            .I3(n59484), .O(n19974[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6470_12_lut (.I0(GND_net), .I1(n18922[9]), .I2(n831_adj_5588), 
            .I3(n60387), .O(n18534[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[8]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6470_12 (.CI(n60387), .I0(n18922[9]), .I1(n831_adj_5588), 
            .CO(n60388));
    SB_LUT4 add_6470_11_lut (.I0(GND_net), .I1(n18922[8]), .I2(n758_adj_5590), 
            .I3(n60386), .O(n18534[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_11 (.CI(n60386), .I0(n18922[8]), .I1(n758_adj_5590), 
            .CO(n60387));
    SB_CARRY add_16_9 (.CI(n58937), .I0(\PID_CONTROLLER.integral [7]), .I1(n207[11]), 
            .CO(n58938));
    SB_CARRY add_6580_5 (.CI(n59484), .I0(n20132[2]), .I1(n335_adj_5587), 
            .CO(n59485));
    SB_LUT4 add_6580_4_lut (.I0(GND_net), .I1(n20132[1]), .I2(n262_adj_5591), 
            .I3(n59483), .O(n19974[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6470_10_lut (.I0(GND_net), .I1(n18922[7]), .I2(n685_adj_5592), 
            .I3(n60385), .O(n18534[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_10 (.CI(n60385), .I0(n18922[7]), .I1(n685_adj_5592), 
            .CO(n60386));
    SB_LUT4 mult_24_i565_2_lut (.I0(\Ki[11] ), .I1(n347_adj_31), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_5593));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6470_9_lut (.I0(GND_net), .I1(n18922[6]), .I2(n612_adj_5594), 
            .I3(n60384), .O(n18534[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_4 (.CI(n59483), .I0(n20132[1]), .I1(n262_adj_5591), 
            .CO(n59484));
    SB_CARRY add_6470_9 (.CI(n60384), .I0(n18922[6]), .I1(n612_adj_5594), 
            .CO(n60385));
    SB_LUT4 mult_23_i61_2_lut (.I0(\Kp[1] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_5595));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6580_3_lut (.I0(GND_net), .I1(n20132[0]), .I2(n189_adj_5596), 
            .I3(n59482), .O(n19974[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_3 (.CI(n59482), .I0(n20132[0]), .I1(n189_adj_5596), 
            .CO(n59483));
    SB_LUT4 mult_23_i14_2_lut (.I0(\Kp[0] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5597));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6580_2_lut (.I0(GND_net), .I1(n47_adj_5598), .I2(n116_adj_5599), 
            .I3(GND_net), .O(n19974[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6470_8_lut (.I0(GND_net), .I1(n18922[5]), .I2(n539_adj_5600), 
            .I3(n60383), .O(n18534[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_2 (.CI(GND_net), .I0(n47_adj_5598), .I1(n116_adj_5599), 
            .CO(n59482));
    SB_CARRY add_6470_8 (.CI(n60383), .I0(n18922[5]), .I1(n539_adj_5600), 
            .CO(n60384));
    SB_LUT4 add_6470_7_lut (.I0(GND_net), .I1(n18922[4]), .I2(n466_adj_5601), 
            .I3(n60382), .O(n18534[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_7 (.CI(n60382), .I0(n18922[4]), .I1(n466_adj_5601), 
            .CO(n60383));
    SB_LUT4 add_6470_6_lut (.I0(GND_net), .I1(n18922[3]), .I2(n393_adj_5602), 
            .I3(n60381), .O(n18534[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_6 (.CI(n60381), .I0(n18922[3]), .I1(n393_adj_5602), 
            .CO(n60382));
    SB_LUT4 add_6289_20_lut (.I0(GND_net), .I1(n15965[17]), .I2(GND_net), 
            .I3(n59481), .O(n15206[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_19_lut (.I0(GND_net), .I1(n15965[16]), .I2(GND_net), 
            .I3(n59480), .O(n15206[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i73_2_lut (.I0(\Ki[1] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_5603));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6470_5_lut (.I0(GND_net), .I1(n18922[2]), .I2(n320_adj_5604), 
            .I3(n60380), .O(n18534[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_5 (.CI(n60380), .I0(n18922[2]), .I1(n320_adj_5604), 
            .CO(n60381));
    SB_LUT4 add_6470_4_lut (.I0(GND_net), .I1(n18922[1]), .I2(n247_adj_5605), 
            .I3(n60379), .O(n18534[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_4 (.CI(n60379), .I0(n18922[1]), .I1(n247_adj_5605), 
            .CO(n60380));
    SB_LUT4 add_6470_3_lut (.I0(GND_net), .I1(n18922[0]), .I2(n174_adj_5606), 
            .I3(n60378), .O(n18534[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_3 (.CI(n60378), .I0(n18922[0]), .I1(n174_adj_5606), 
            .CO(n60379));
    SB_LUT4 mult_23_i110_2_lut (.I0(\Kp[2] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_5607));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6470_2_lut (.I0(GND_net), .I1(n32_adj_5608), .I2(n101_adj_5609), 
            .I3(GND_net), .O(n18534[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i159_2_lut (.I0(\Kp[3] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_5610));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6470_2 (.CI(GND_net), .I0(n32_adj_5608), .I1(n101_adj_5609), 
            .CO(n60378));
    SB_LUT4 add_6496_14_lut (.I0(GND_net), .I1(n19256[11]), .I2(n980_adj_5611), 
            .I3(n60377), .O(n18922[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i208_2_lut (.I0(\Kp[4] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_5612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[9]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6496_13_lut (.I0(GND_net), .I1(n19256[10]), .I2(n907_adj_5614), 
            .I3(n60376), .O(n18922[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_13 (.CI(n60376), .I0(n19256[10]), .I1(n907_adj_5614), 
            .CO(n60377));
    SB_LUT4 add_6496_12_lut (.I0(GND_net), .I1(n19256[9]), .I2(n834_adj_5615), 
            .I3(n60375), .O(n18922[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_12 (.CI(n60375), .I0(n19256[9]), .I1(n834_adj_5615), 
            .CO(n60376));
    SB_LUT4 mult_23_i257_2_lut (.I0(\Kp[5] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_5616));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6496_11_lut (.I0(GND_net), .I1(n19256[8]), .I2(n761_adj_5617), 
            .I3(n60374), .O(n18922[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[10]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6289_19 (.CI(n59480), .I0(n15965[16]), .I1(GND_net), 
            .CO(n59481));
    SB_LUT4 add_6289_18_lut (.I0(GND_net), .I1(n15965[15]), .I2(GND_net), 
            .I3(n59479), .O(n15206[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i306_2_lut (.I0(\Kp[6] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_5619));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6289_18 (.CI(n59479), .I0(n15965[15]), .I1(GND_net), 
            .CO(n59480));
    SB_CARRY add_6496_11 (.CI(n60374), .I0(n19256[8]), .I1(n761_adj_5617), 
            .CO(n60375));
    SB_LUT4 add_6496_10_lut (.I0(GND_net), .I1(n19256[7]), .I2(n688_adj_5620), 
            .I3(n60373), .O(n18922[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i355_2_lut (.I0(\Kp[7] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_5621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i404_2_lut (.I0(\Kp[8] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_5622));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6289_17_lut (.I0(GND_net), .I1(n15965[14]), .I2(GND_net), 
            .I3(n59478), .O(n15206[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i453_2_lut (.I0(\Kp[9] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_5623));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i453_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6496_10 (.CI(n60373), .I0(n19256[7]), .I1(n688_adj_5620), 
            .CO(n60374));
    SB_LUT4 add_16_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n207[10]), .I3(n58936), .O(n233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_17 (.CI(n59478), .I0(n15965[14]), .I1(GND_net), 
            .CO(n59479));
    SB_LUT4 add_6496_9_lut (.I0(GND_net), .I1(n19256[6]), .I2(n615_adj_5624), 
            .I3(n60372), .O(n18922[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_9 (.CI(n60372), .I0(n19256[6]), .I1(n615_adj_5624), 
            .CO(n60373));
    SB_CARRY add_16_8 (.CI(n58936), .I0(\PID_CONTROLLER.integral [6]), .I1(n207[10]), 
            .CO(n58937));
    SB_LUT4 unary_minus_33_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[11]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i502_2_lut (.I0(\Kp[10] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_5626));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6496_8_lut (.I0(GND_net), .I1(n19256[5]), .I2(n542_adj_5627), 
            .I3(n60371), .O(n18922[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i551_2_lut (.I0(\Kp[11] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_5628));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[12]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i600_2_lut (.I0(\Kp[12] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_5630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i600_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_6 (.CI(n58911), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n58912));
    SB_LUT4 add_6289_16_lut (.I0(GND_net), .I1(n15965[13]), .I2(n1108_adj_5631), 
            .I3(n59477), .O(n15206[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i649_2_lut (.I0(\Kp[13] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_5632));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i649_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6289_16 (.CI(n59477), .I0(n15965[13]), .I1(n1108_adj_5631), 
            .CO(n59478));
    SB_CARRY add_6496_8 (.CI(n60371), .I0(n19256[5]), .I1(n542_adj_5627), 
            .CO(n60372));
    SB_LUT4 add_6289_15_lut (.I0(GND_net), .I1(n15965[12]), .I2(n1035_adj_5633), 
            .I3(n59476), .O(n15206[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6496_7_lut (.I0(GND_net), .I1(n19256[4]), .I2(n469_adj_5634), 
            .I3(n60370), .O(n18922[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i698_2_lut (.I0(\Kp[14] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_5635));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[13]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i747_2_lut (.I0(\Kp[15] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_5637));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i747_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6496_7 (.CI(n60370), .I0(n19256[4]), .I1(n469_adj_5634), 
            .CO(n60371));
    SB_LUT4 add_6496_6_lut (.I0(GND_net), .I1(n19256[3]), .I2(n396_adj_5638), 
            .I3(n60369), .O(n18922[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_6 (.CI(n60369), .I0(n19256[3]), .I1(n396_adj_5638), 
            .CO(n60370));
    SB_LUT4 add_6496_5_lut (.I0(GND_net), .I1(n19256[2]), .I2(n323_adj_5639), 
            .I3(n60368), .O(n18922[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_5 (.CI(n60368), .I0(n19256[2]), .I1(n323_adj_5639), 
            .CO(n60369));
    SB_LUT4 add_6496_4_lut (.I0(GND_net), .I1(n19256[1]), .I2(n250_adj_5640), 
            .I3(n60367), .O(n18922[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n207[9]), .I3(n58935), .O(n233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[14]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i122_2_lut (.I0(\Ki[2] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_5642));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i122_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6289_15 (.CI(n59476), .I0(n15965[12]), .I1(n1035_adj_5633), 
            .CO(n59477));
    SB_LUT4 add_6289_14_lut (.I0(GND_net), .I1(n15965[11]), .I2(n962_adj_5643), 
            .I3(n59475), .O(n15206[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_14 (.CI(n59475), .I0(n15965[11]), .I1(n962_adj_5643), 
            .CO(n59476));
    SB_LUT4 add_6289_13_lut (.I0(GND_net), .I1(n15965[10]), .I2(n889_adj_5644), 
            .I3(n59474), .O(n15206[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_4 (.CI(n60367), .I0(n19256[1]), .I1(n250_adj_5640), 
            .CO(n60368));
    SB_LUT4 add_6496_3_lut (.I0(GND_net), .I1(n19256[0]), .I2(n177_adj_5645), 
            .I3(n60366), .O(n18922[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_3 (.CI(n60366), .I0(n19256[0]), .I1(n177_adj_5645), 
            .CO(n60367));
    SB_CARRY add_6289_13 (.CI(n59474), .I0(n15965[10]), .I1(n889_adj_5644), 
            .CO(n59475));
    SB_LUT4 unary_minus_33_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[15]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6496_2_lut (.I0(GND_net), .I1(n35_adj_5647), .I2(n104_adj_5648), 
            .I3(GND_net), .O(n18922[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60327_2_lut (.I0(PWMLimit[23]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75323));
    defparam i60327_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6496_2 (.CI(GND_net), .I0(n35_adj_5647), .I1(n104_adj_5648), 
            .CO(n60366));
    SB_LUT4 add_6601_8_lut (.I0(GND_net), .I1(n20289[5]), .I2(n560_adj_5649), 
            .I3(n60365), .O(n20178[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_12_lut (.I0(GND_net), .I1(n15965[9]), .I2(n816_adj_5650), 
            .I3(n59473), .O(n15206[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[16]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6289_12 (.CI(n59473), .I0(n15965[9]), .I1(n816_adj_5650), 
            .CO(n59474));
    SB_LUT4 mult_24_i171_2_lut (.I0(\Ki[3] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_5652));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6289_11_lut (.I0(GND_net), .I1(n15965[8]), .I2(n743_adj_5653), 
            .I3(n59472), .O(n15206[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6601_7_lut (.I0(GND_net), .I1(n20289[4]), .I2(n487_adj_5654), 
            .I3(n60364), .O(n20178[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_11 (.CI(n59472), .I0(n15965[8]), .I1(n743_adj_5653), 
            .CO(n59473));
    SB_CARRY add_6601_7 (.CI(n60364), .I0(n20289[4]), .I1(n487_adj_5654), 
            .CO(n60365));
    SB_LUT4 add_6601_6_lut (.I0(GND_net), .I1(n20289[3]), .I2(n414_adj_5655), 
            .I3(n60363), .O(n20178[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_6 (.CI(n60363), .I0(n20289[3]), .I1(n414_adj_5655), 
            .CO(n60364));
    SB_LUT4 add_6289_10_lut (.I0(GND_net), .I1(n15965[7]), .I2(n670_adj_5656), 
            .I3(n59471), .O(n15206[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6601_5_lut (.I0(GND_net), .I1(n20289[2]), .I2(n341_adj_5657), 
            .I3(n60362), .O(n20178[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[17]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_16_7 (.CI(n58935), .I0(\PID_CONTROLLER.integral [5]), .I1(n207[9]), 
            .CO(n58936));
    SB_CARRY add_6289_10 (.CI(n59471), .I0(n15965[7]), .I1(n670_adj_5656), 
            .CO(n59472));
    SB_CARRY add_6601_5 (.CI(n60362), .I0(n20289[2]), .I1(n341_adj_5657), 
            .CO(n60363));
    SB_CARRY sub_15_add_2_5 (.CI(n58910), .I0(setpoint[3]), .I1(n17), 
            .CO(n58911));
    SB_LUT4 mult_24_i220_2_lut (.I0(\Ki[4] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_5660));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[18]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6601_4_lut (.I0(GND_net), .I1(n20289[1]), .I2(n268_adj_5662), 
            .I3(n60361), .O(n20178[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_4 (.CI(n60361), .I0(n20289[1]), .I1(n268_adj_5662), 
            .CO(n60362));
    SB_LUT4 unary_minus_33_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[19]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[20]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6601_3_lut (.I0(GND_net), .I1(n20289[0]), .I2(n195_adj_5665), 
            .I3(n60360), .O(n20178[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[21]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i269_2_lut (.I0(\Ki[5] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_5667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i318_2_lut (.I0(\Ki[6] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_5668));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n207[8]), .I3(n58934), .O(n233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_3 (.CI(n60360), .I0(n20289[0]), .I1(n195_adj_5665), 
            .CO(n60361));
    SB_LUT4 add_6289_9_lut (.I0(GND_net), .I1(n15965[6]), .I2(n597_adj_5669), 
            .I3(n59470), .O(n15206[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_9 (.CI(n59470), .I0(n15965[6]), .I1(n597_adj_5669), 
            .CO(n59471));
    SB_LUT4 mult_24_i367_2_lut (.I0(\Ki[7] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_5670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[22]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6601_2_lut (.I0(GND_net), .I1(n53_adj_5672), .I2(n122_adj_5673), 
            .I3(GND_net), .O(n20178[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_2 (.CI(GND_net), .I0(n53_adj_5672), .I1(n122_adj_5673), 
            .CO(n60360));
    SB_LUT4 add_6520_13_lut (.I0(GND_net), .I1(n19540[10]), .I2(n910_adj_5674), 
            .I3(n60359), .O(n19256[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6520_12_lut (.I0(GND_net), .I1(n19540[9]), .I2(n837_adj_5675), 
            .I3(n60358), .O(n19256[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_12 (.CI(n60358), .I0(n19540[9]), .I1(n837_adj_5675), 
            .CO(n60359));
    SB_LUT4 unary_minus_33_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5702[23]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i416_2_lut (.I0(\Ki[8] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_5677));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i416_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_6 (.CI(n58934), .I0(\PID_CONTROLLER.integral [4]), .I1(n207[8]), 
            .CO(n58935));
    SB_LUT4 add_6520_11_lut (.I0(GND_net), .I1(n19540[8]), .I2(n764_adj_5678), 
            .I3(n60357), .O(n19256[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i465_2_lut (.I0(\Ki[9] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_5679));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31191_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45282));   // verilog/motorControl.v(42[14] 73[8])
    defparam i31191_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6289_8_lut (.I0(GND_net), .I1(n15965[5]), .I2(n524_adj_5680), 
            .I3(n59469), .O(n15206[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_8 (.CI(n59469), .I0(n15965[5]), .I1(n524_adj_5680), 
            .CO(n59470));
    SB_LUT4 add_6289_7_lut (.I0(GND_net), .I1(n15965[4]), .I2(n451_adj_5681), 
            .I3(n59468), .O(n15206[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_7 (.CI(n59468), .I0(n15965[4]), .I1(n451_adj_5681), 
            .CO(n59469));
    SB_LUT4 add_6289_6_lut (.I0(GND_net), .I1(n15965[3]), .I2(n378_adj_5682), 
            .I3(n59467), .O(n15206[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_6 (.CI(n59467), .I0(n15965[3]), .I1(n378_adj_5682), 
            .CO(n59468));
    SB_LUT4 add_6289_5_lut (.I0(GND_net), .I1(n15965[2]), .I2(n305_adj_5683), 
            .I3(n59466), .O(n15206[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_5 (.CI(n59466), .I0(n15965[2]), .I1(n305_adj_5683), 
            .CO(n59467));
    SB_LUT4 add_6289_4_lut (.I0(GND_net), .I1(n15965[1]), .I2(n232_adj_5684), 
            .I3(n59465), .O(n15206[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_4 (.CI(n59465), .I0(n15965[1]), .I1(n232_adj_5684), 
            .CO(n59466));
    SB_LUT4 add_6289_3_lut (.I0(GND_net), .I1(n15965[0]), .I2(n159_adj_5685), 
            .I3(n59464), .O(n15206[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_3 (.CI(n59464), .I0(n15965[0]), .I1(n159_adj_5685), 
            .CO(n59465));
    SB_LUT4 mult_23_i59_2_lut (.I0(\Kp[1] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_5686));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6289_2_lut (.I0(GND_net), .I1(n17_adj_5687), .I2(n86_adj_5686), 
            .I3(GND_net), .O(n15206[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_2 (.CI(GND_net), .I0(n17_adj_5687), .I1(n86_adj_5686), 
            .CO(n59464));
    SB_LUT4 mult_23_i12_2_lut (.I0(\Kp[0] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5687));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i12_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6520_11 (.CI(n60357), .I0(n19540[8]), .I1(n764_adj_5678), 
            .CO(n60358));
    SB_LUT4 add_6520_10_lut (.I0(GND_net), .I1(n19540[7]), .I2(n691_adj_5679), 
            .I3(n60356), .O(n19256[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_10 (.CI(n60356), .I0(n19540[7]), .I1(n691_adj_5679), 
            .CO(n60357));
    SB_LUT4 mult_23_i108_2_lut (.I0(\Kp[2] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_5685));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_9_lut (.I0(GND_net), .I1(n19540[6]), .I2(n618_adj_5677), 
            .I3(n60355), .O(n19256[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i120_2_lut (.I0(\Kp[2] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i157_2_lut (.I0(\Kp[3] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_5684));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i206_2_lut (.I0(\Kp[4] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_5683));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i255_2_lut (.I0(\Kp[5] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_5682));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[23]), 
            .I3(n59122), .O(n535[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[22]), 
            .I3(n59121), .O(n535[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_9 (.CI(n60355), .I0(n19540[6]), .I1(n618_adj_5677), 
            .CO(n60356));
    SB_LUT4 mult_23_i304_2_lut (.I0(\Kp[6] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_5681));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_8_lut (.I0(GND_net), .I1(n19540[5]), .I2(n545_adj_5670), 
            .I3(n60354), .O(n19256[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_8 (.CI(n60354), .I0(n19540[5]), .I1(n545_adj_5670), 
            .CO(n60355));
    SB_LUT4 mult_23_i353_2_lut (.I0(\Kp[7] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_5680));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_7_lut (.I0(GND_net), .I1(n19540[4]), .I2(n472_adj_5668), 
            .I3(n60353), .O(n19256[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_7 (.CI(n60353), .I0(n19540[4]), .I1(n472_adj_5668), 
            .CO(n60354));
    SB_LUT4 add_6520_6_lut (.I0(GND_net), .I1(n19540[3]), .I2(n399_adj_5667), 
            .I3(n60352), .O(n19256[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i514_2_lut (.I0(\Ki[10] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_5678));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i514_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_33_add_3_24 (.CI(n59121), .I0(GND_net), .I1(n1_adj_5702[22]), 
            .CO(n59122));
    SB_LUT4 unary_minus_33_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[21]), 
            .I3(n59120), .O(n535[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i563_2_lut (.I0(\Ki[11] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_5675));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i612_2_lut (.I0(\Ki[12] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_5674));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i83_2_lut (.I0(\Kp[1] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_5673));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i36_2_lut (.I0(\Kp[0] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_5672));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i36_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_33_add_3_23 (.CI(n59120), .I0(GND_net), .I1(n1_adj_5702[21]), 
            .CO(n59121));
    SB_LUT4 unary_minus_33_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[20]), 
            .I3(n59119), .O(n535[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_22 (.CI(n59119), .I0(GND_net), .I1(n1_adj_5702[20]), 
            .CO(n59120));
    SB_LUT4 mux_21_i1_3_lut (.I0(n233[0]), .I1(n285[0]), .I2(n284), .I3(GND_net), 
            .O(n310[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[19]), 
            .I3(n59118), .O(n535[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i402_2_lut (.I0(\Kp[8] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_5669));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_33_add_3_21 (.CI(n59118), .I0(GND_net), .I1(n1_adj_5702[19]), 
            .CO(n59119));
    SB_LUT4 unary_minus_33_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[18]), 
            .I3(n59117), .O(n535[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n207[7]), .I3(n58933), .O(n233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_6 (.CI(n60352), .I0(n19540[3]), .I1(n399_adj_5667), 
            .CO(n60353));
    SB_LUT4 add_6520_5_lut (.I0(GND_net), .I1(n19540[2]), .I2(n326_adj_5660), 
            .I3(n60351), .O(n19256[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i132_2_lut (.I0(\Kp[2] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_5665));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i181_2_lut (.I0(\Kp[3] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_5662));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i181_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_33_add_3_20 (.CI(n59117), .I0(GND_net), .I1(n1_adj_5702[18]), 
            .CO(n59118));
    SB_LUT4 unary_minus_33_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[17]), 
            .I3(n59116), .O(n535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_5 (.CI(n60351), .I0(n19540[2]), .I1(n326_adj_5660), 
            .CO(n60352));
    SB_CARRY add_16_5 (.CI(n58933), .I0(\PID_CONTROLLER.integral [3]), .I1(n207[7]), 
            .CO(n58934));
    SB_LUT4 add_16_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n207[6]), .I3(n58932), .O(n233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_4 (.CI(n58909), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n58910));
    SB_CARRY sub_15_add_2_3 (.CI(n58908), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n58909));
    SB_LUT4 add_6520_4_lut (.I0(GND_net), .I1(n19540[1]), .I2(n253_adj_5652), 
            .I3(n60350), .O(n19256[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_19 (.CI(n59116), .I0(GND_net), .I1(n1_adj_5702[17]), 
            .CO(n59117));
    SB_LUT4 mult_23_i230_2_lut (.I0(\Kp[4] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_5657));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i1_3_lut (.I0(n310[0]), .I1(IntegralLimit[0]), .I2(n258), 
            .I3(GND_net), .O(n359));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[16]), 
            .I3(n59115), .O(n535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i2_2_lut (.I0(\Ki[0] ), .I1(n359), .I2(GND_net), .I3(GND_net), 
            .O(n46[0]));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11882_bdd_4_lut (.I0(n11882), .I1(n75323), .I2(setpoint[23]), 
            .I3(n4736), .O(n79534));
    defparam n11882_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_CARRY unary_minus_33_add_3_18 (.CI(n59115), .I0(GND_net), .I1(n1_adj_5702[16]), 
            .CO(n59116));
    SB_LUT4 unary_minus_33_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[15]), 
            .I3(n59114), .O(n535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(\motor_state[0] ), 
            .CO(n58908));
    SB_CARRY add_16_4 (.CI(n58932), .I0(\PID_CONTROLLER.integral [2]), .I1(n207[6]), 
            .CO(n58933));
    SB_LUT4 add_16_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n207[5]), .I3(n58931), .O(n233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_4 (.CI(n60350), .I0(n19540[1]), .I1(n253_adj_5652), 
            .CO(n60351));
    SB_LUT4 add_6520_3_lut (.I0(GND_net), .I1(n19540[0]), .I2(n180_adj_5642), 
            .I3(n60349), .O(n19256[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_19_lut (.I0(GND_net), .I1(n16648[16]), .I2(GND_net), 
            .I3(n59444), .O(n15965[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i451_2_lut (.I0(\Kp[9] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_5656));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_18_lut (.I0(GND_net), .I1(n16648[15]), .I2(GND_net), 
            .I3(n59443), .O(n15965[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i279_2_lut (.I0(\Kp[5] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_5655));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i279_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6326_18 (.CI(n59443), .I0(n16648[15]), .I1(GND_net), 
            .CO(n59444));
    SB_LUT4 mult_23_i328_2_lut (.I0(\Kp[6] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_5654));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_17_lut (.I0(GND_net), .I1(n16648[14]), .I2(GND_net), 
            .I3(n59442), .O(n15965[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_17 (.CI(n59442), .I0(n16648[14]), .I1(GND_net), 
            .CO(n59443));
    SB_LUT4 mult_23_i500_2_lut (.I0(\Kp[10] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_5653));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_33_add_3_17 (.CI(n59114), .I0(GND_net), .I1(n1_adj_5702[15]), 
            .CO(n59115));
    SB_LUT4 unary_minus_33_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[14]), 
            .I3(n59113), .O(n535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_16_lut (.I0(GND_net), .I1(n16648[13]), .I2(n1111_adj_5637), 
            .I3(n59441), .O(n15965[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i549_2_lut (.I0(\Kp[11] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_5650));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6326_16 (.CI(n59441), .I0(n16648[13]), .I1(n1111_adj_5637), 
            .CO(n59442));
    SB_CARRY unary_minus_33_add_3_16 (.CI(n59113), .I0(GND_net), .I1(n1_adj_5702[14]), 
            .CO(n59114));
    SB_LUT4 unary_minus_33_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[13]), 
            .I3(n59112), .O(n535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_3 (.CI(n58931), .I0(\PID_CONTROLLER.integral [1]), .I1(n207[5]), 
            .CO(n58932));
    SB_LUT4 add_6326_15_lut (.I0(GND_net), .I1(n16648[12]), .I2(n1038_adj_5635), 
            .I3(n59440), .O(n15965[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_15 (.CI(n59440), .I0(n16648[12]), .I1(n1038_adj_5635), 
            .CO(n59441));
    SB_LUT4 add_6326_14_lut (.I0(GND_net), .I1(n16648[11]), .I2(n965_adj_5632), 
            .I3(n59439), .O(n15965[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_14 (.CI(n59439), .I0(n16648[11]), .I1(n965_adj_5632), 
            .CO(n59440));
    SB_CARRY unary_minus_33_add_3_15 (.CI(n59112), .I0(GND_net), .I1(n1_adj_5702[13]), 
            .CO(n59113));
    SB_LUT4 mult_23_i377_2_lut (.I0(\Kp[7] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_5649));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_13_lut (.I0(GND_net), .I1(n16648[10]), .I2(n892_adj_5630), 
            .I3(n59438), .O(n15965[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[12]), 
            .I3(n59111), .O(n535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_13 (.CI(n59438), .I0(n16648[10]), .I1(n892_adj_5630), 
            .CO(n59439));
    SB_LUT4 mult_24_i71_2_lut (.I0(\Ki[1] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_5648));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_12_lut (.I0(GND_net), .I1(n16648[9]), .I2(n819_adj_5628), 
            .I3(n59437), .O(n15965[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i24_2_lut (.I0(\Ki[0] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5647));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i120_2_lut (.I0(\Ki[2] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_5645));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6326_12 (.CI(n59437), .I0(n16648[9]), .I1(n819_adj_5628), 
            .CO(n59438));
    SB_LUT4 add_6326_11_lut (.I0(GND_net), .I1(n16648[8]), .I2(n746_adj_5626), 
            .I3(n59436), .O(n15965[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i2_2_lut (.I0(\Kp[0] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n360[0]));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6326_11 (.CI(n59436), .I0(n16648[8]), .I1(n746_adj_5626), 
            .CO(n59437));
    SB_CARRY unary_minus_33_add_3_14 (.CI(n59111), .I0(GND_net), .I1(n1_adj_5702[12]), 
            .CO(n59112));
    SB_LUT4 unary_minus_33_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[11]), 
            .I3(n59110), .O(n535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_10_lut (.I0(GND_net), .I1(n16648[7]), .I2(n673_adj_5623), 
            .I3(n59435), .O(n15965[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_10 (.CI(n59435), .I0(n16648[7]), .I1(n673_adj_5623), 
            .CO(n59436));
    SB_LUT4 add_16_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n207[4]), .I3(GND_net), .O(n233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n207[4]), .CO(n58931));
    SB_LUT4 add_6326_9_lut (.I0(GND_net), .I1(n16648[6]), .I2(n600_adj_5622), 
            .I3(n59434), .O(n15965[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_9 (.CI(n59434), .I0(n16648[6]), .I1(n600_adj_5622), 
            .CO(n59435));
    SB_LUT4 add_6326_8_lut (.I0(GND_net), .I1(n16648[5]), .I2(n527_adj_5621), 
            .I3(n59433), .O(n15965[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i598_2_lut (.I0(\Kp[12] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_5644));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i647_2_lut (.I0(\Kp[13] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_5643));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i169_2_lut (.I0(\Ki[3] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_5640));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i218_2_lut (.I0(\Ki[4] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_5639));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6520_3 (.CI(n60349), .I0(n19540[0]), .I1(n180_adj_5642), 
            .CO(n60350));
    SB_LUT4 mult_24_i267_2_lut (.I0(\Ki[5] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_5638));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6326_8 (.CI(n59433), .I0(n16648[5]), .I1(n527_adj_5621), 
            .CO(n59434));
    SB_LUT4 mult_23_i169_2_lut (.I0(\Kp[3] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_7_lut (.I0(GND_net), .I1(n16648[4]), .I2(n454_adj_5619), 
            .I3(n59432), .O(n15965[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_13 (.CI(n59110), .I0(GND_net), .I1(n1_adj_5702[11]), 
            .CO(n59111));
    SB_CARRY add_6326_7 (.CI(n59432), .I0(n16648[4]), .I1(n454_adj_5619), 
            .CO(n59433));
    SB_LUT4 unary_minus_33_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[10]), 
            .I3(n59109), .O(n535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i218_2_lut (.I0(\Kp[4] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_6_lut (.I0(GND_net), .I1(n16648[3]), .I2(n381_adj_5616), 
            .I3(n59431), .O(n15965[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n58930), .O(n207[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_6 (.CI(n59431), .I0(n16648[3]), .I1(n381_adj_5616), 
            .CO(n59432));
    SB_CARRY unary_minus_33_add_3_12 (.CI(n59109), .I0(GND_net), .I1(n1_adj_5702[10]), 
            .CO(n59110));
    SB_LUT4 unary_minus_33_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[9]), 
            .I3(n59108), .O(n535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_5_lut (.I0(GND_net), .I1(n16648[2]), .I2(n308_adj_5612), 
            .I3(n59430), .O(n15965[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_5 (.CI(n59430), .I0(n16648[2]), .I1(n308_adj_5612), 
            .CO(n59431));
    SB_LUT4 mult_24_i316_2_lut (.I0(\Ki[6] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_5634));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_4_lut (.I0(GND_net), .I1(n16648[1]), .I2(n235_adj_5610), 
            .I3(n59429), .O(n15965[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_4 (.CI(n59429), .I0(n16648[1]), .I1(n235_adj_5610), 
            .CO(n59430));
    SB_LUT4 add_6326_3_lut (.I0(GND_net), .I1(n16648[0]), .I2(n162_adj_5607), 
            .I3(n59428), .O(n15965[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_11 (.CI(n59108), .I0(GND_net), .I1(n1_adj_5702[9]), 
            .CO(n59109));
    SB_LUT4 mult_23_i696_2_lut (.I0(\Kp[14] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_5633));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_2_lut (.I0(GND_net), .I1(n38_adj_32), .I2(n107_adj_5603), 
            .I3(GND_net), .O(n19256[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n58929), .O(n207[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_3 (.CI(n59428), .I0(n16648[0]), .I1(n162_adj_5607), 
            .CO(n59429));
    SB_LUT4 mult_23_i745_2_lut (.I0(\Kp[15] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_5631));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i365_2_lut (.I0(\Ki[7] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_5627));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6326_2_lut (.I0(GND_net), .I1(n20_adj_5597), .I2(n89_adj_5595), 
            .I3(GND_net), .O(n15965[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i414_2_lut (.I0(\Ki[8] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_5624));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i414_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6326_2 (.CI(GND_net), .I0(n20_adj_5597), .I1(n89_adj_5595), 
            .CO(n59428));
    SB_CARRY add_6520_2 (.CI(GND_net), .I0(n38_adj_32), .I1(n107_adj_5603), 
            .CO(n60349));
    SB_LUT4 add_6542_12_lut (.I0(GND_net), .I1(n19778[9]), .I2(n840_adj_5593), 
            .I3(n60348), .O(n19540[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[8]), 
            .I3(n59107), .O(n535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_10 (.CI(n59107), .I0(GND_net), .I1(n1_adj_5702[8]), 
            .CO(n59108));
    SB_LUT4 unary_minus_33_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[7]), 
            .I3(n59106), .O(n535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_9 (.CI(n59106), .I0(GND_net), .I1(n1_adj_5702[7]), 
            .CO(n59107));
    SB_LUT4 mult_24_i463_2_lut (.I0(\Ki[9] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_5620));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i512_2_lut (.I0(\Ki[10] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_5617));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i561_2_lut (.I0(\Ki[11] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_5615));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[6]), 
            .I3(n59105), .O(n535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i610_2_lut (.I0(\Ki[12] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_5614));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i659_2_lut (.I0(\Ki[13] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_5611));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i69_2_lut (.I0(\Ki[1] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_5609));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i69_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_33_add_3_8 (.CI(n59105), .I0(GND_net), .I1(n1_adj_5702[6]), 
            .CO(n59106));
    SB_LUT4 mult_24_i22_2_lut (.I0(\Ki[0] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_5608));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6542_11_lut (.I0(GND_net), .I1(n19778[8]), .I2(n767_adj_5582), 
            .I3(n60347), .O(n19540[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[5]), 
            .I3(n59104), .O(n535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i118_2_lut (.I0(\Ki[2] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_5606));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i167_2_lut (.I0(\Ki[3] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_5605));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_24 (.CI(n58929), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n58930));
    SB_LUT4 mult_24_i216_2_lut (.I0(\Ki[4] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_5604));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_33_add_3_7 (.CI(n59104), .I0(GND_net), .I1(n1_adj_5702[5]), 
            .CO(n59105));
    SB_LUT4 mult_24_i265_2_lut (.I0(\Ki[5] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_5602));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i314_2_lut (.I0(\Ki[6] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_5601));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i363_2_lut (.I0(\Ki[7] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_5600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[4]), 
            .I3(n59103), .O(n535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n58928), .O(n207[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_6 (.CI(n59103), .I0(GND_net), .I1(n1_adj_5702[4]), 
            .CO(n59104));
    SB_LUT4 unary_minus_33_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[3]), 
            .I3(n59102), .O(n535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i79_2_lut (.I0(\Ki[1] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_5599));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i79_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6542_11 (.CI(n60347), .I0(n19778[8]), .I1(n767_adj_5582), 
            .CO(n60348));
    SB_LUT4 mult_24_i32_2_lut (.I0(\Ki[0] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_5598));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6542_10_lut (.I0(GND_net), .I1(n19778[7]), .I2(n694_adj_5568), 
            .I3(n60346), .O(n19540[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_5 (.CI(n59102), .I0(GND_net), .I1(n1_adj_5702[3]), 
            .CO(n59103));
    SB_LUT4 unary_minus_33_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[2]), 
            .I3(n59101), .O(n535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_10 (.CI(n60346), .I0(n19778[7]), .I1(n694_adj_5568), 
            .CO(n60347));
    SB_CARRY unary_minus_33_add_3_4 (.CI(n59101), .I0(GND_net), .I1(n1_adj_5702[2]), 
            .CO(n59102));
    SB_LUT4 mult_24_i128_2_lut (.I0(\Ki[2] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_5596));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i412_2_lut (.I0(\Ki[8] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_5594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i461_2_lut (.I0(\Ki[9] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_5592));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i177_2_lut (.I0(\Ki[3] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_5591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i510_2_lut (.I0(\Ki[10] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_5590));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i559_2_lut (.I0(\Ki[11] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_5588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[1]), 
            .I3(n59100), .O(n535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_3 (.CI(n59100), .I0(GND_net), .I1(n1_adj_5702[1]), 
            .CO(n59101));
    SB_LUT4 add_6542_9_lut (.I0(GND_net), .I1(n19778[6]), .I2(n621_adj_5564), 
            .I3(n60345), .O(n19540[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i226_2_lut (.I0(\Ki[4] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_5587));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6596_9_lut (.I0(GND_net), .I1(n20256[6]), .I2(n630_adj_5562), 
            .I3(n59409), .O(n20132[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6596_8_lut (.I0(GND_net), .I1(n20256[5]), .I2(n557_adj_5561), 
            .I3(n59408), .O(n20132[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_8 (.CI(n59408), .I0(n20256[5]), .I1(n557_adj_5561), 
            .CO(n59409));
    SB_LUT4 add_6596_7_lut (.I0(GND_net), .I1(n20256[4]), .I2(n484_adj_5560), 
            .I3(n59407), .O(n20132[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_7 (.CI(n59407), .I0(n20256[4]), .I1(n484_adj_5560), 
            .CO(n59408));
    SB_CARRY sub_15_add_2_23 (.CI(n58928), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n58929));
    SB_LUT4 add_6596_6_lut (.I0(GND_net), .I1(n20256[3]), .I2(n411), .I3(n59406), 
            .O(n20132[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(n12), 
            .I3(n58927), .O(n207[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5702[0]), 
            .I3(VCC_net), .O(n535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i275_2_lut (.I0(\Ki[5] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_5584));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6542_9 (.CI(n60345), .I0(n19778[6]), .I1(n621_adj_5564), 
            .CO(n60346));
    SB_LUT4 add_6542_8_lut (.I0(GND_net), .I1(n19778[5]), .I2(n548_adj_5557), 
            .I3(n60344), .O(n19540[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_6 (.CI(n59406), .I0(n20256[3]), .I1(n411), .CO(n59407));
    SB_LUT4 add_6596_5_lut (.I0(GND_net), .I1(n20256[2]), .I2(n338), .I3(n59405), 
            .O(n20132[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_5 (.CI(n59405), .I0(n20256[2]), .I1(n338), .CO(n59406));
    SB_LUT4 add_6596_4_lut (.I0(GND_net), .I1(n20256[1]), .I2(n265), .I3(n59404), 
            .O(n20132[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_4 (.CI(n59404), .I0(n20256[1]), .I1(n265), .CO(n59405));
    SB_LUT4 add_6596_3_lut (.I0(GND_net), .I1(n20256[0]), .I2(n192), .I3(n59403), 
            .O(n20132[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_8 (.CI(n60344), .I0(n19778[5]), .I1(n548_adj_5557), 
            .CO(n60345));
    SB_CARRY sub_15_add_2_22 (.CI(n58927), .I0(setpoint[20]), .I1(n12), 
            .CO(n58928));
    SB_LUT4 mult_24_i608_2_lut (.I0(\Ki[12] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_5583));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n58926), .O(n207[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5702[0]), 
            .CO(n59100));
    SB_CARRY add_6596_3 (.CI(n59403), .I0(n20256[0]), .I1(n192), .CO(n59404));
    SB_LUT4 add_6596_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n20132[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n59403));
    SB_LUT4 add_6361_18_lut (.I0(GND_net), .I1(n17259[15]), .I2(GND_net), 
            .I3(n59402), .O(n16648[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6542_7_lut (.I0(GND_net), .I1(n19778[4]), .I2(n475_adj_5551), 
            .I3(n60343), .O(n19540[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i324_2_lut (.I0(\Ki[6] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_5579));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6361_17_lut (.I0(GND_net), .I1(n17259[14]), .I2(GND_net), 
            .I3(n59401), .O(n16648[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_17 (.CI(n59401), .I0(n17259[14]), .I1(GND_net), 
            .CO(n59402));
    SB_LUT4 add_6361_16_lut (.I0(GND_net), .I1(n17259[13]), .I2(n1114_adj_5550), 
            .I3(n59400), .O(n16648[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(n455[23]), .I1(GND_net), .I2(n1_adj_5701[23]), 
            .I3(n59099), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6361_16 (.CI(n59400), .I0(n17259[13]), .I1(n1114_adj_5550), 
            .CO(n59401));
    SB_LUT4 add_6361_15_lut (.I0(GND_net), .I1(n17259[12]), .I2(n1041_adj_5548), 
            .I3(n59399), .O(n16648[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_15 (.CI(n59399), .I0(n17259[12]), .I1(n1041_adj_5548), 
            .CO(n59400));
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[22]), 
            .I3(n59098), .O(n48[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_24 (.CI(n59098), .I0(GND_net), .I1(n1_adj_5701[22]), 
            .CO(n59099));
    SB_LUT4 add_6361_14_lut (.I0(GND_net), .I1(n17259[11]), .I2(n968_adj_5544), 
            .I3(n59398), .O(n16648[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_14 (.CI(n59398), .I0(n17259[11]), .I1(n968_adj_5544), 
            .CO(n59399));
    SB_LUT4 mult_24_i373_2_lut (.I0(\Ki[7] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_5578));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6361_13_lut (.I0(GND_net), .I1(n17259[10]), .I2(n895_adj_5543), 
            .I3(n59397), .O(n16648[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_13 (.CI(n59397), .I0(n17259[10]), .I1(n895_adj_5543), 
            .CO(n59398));
    SB_LUT4 mult_24_i657_2_lut (.I0(\Ki[13] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_5577));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i422_2_lut (.I0(\Ki[8] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_5576));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6361_12_lut (.I0(GND_net), .I1(n17259[9]), .I2(n822_adj_5542), 
            .I3(n59396), .O(n16648[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_7 (.CI(n60343), .I0(n19778[4]), .I1(n475_adj_5551), 
            .CO(n60344));
    SB_CARRY add_6361_12 (.CI(n59396), .I0(n17259[9]), .I1(n822_adj_5542), 
            .CO(n59397));
    SB_LUT4 add_6361_11_lut (.I0(GND_net), .I1(n17259[8]), .I2(n749_adj_5541), 
            .I3(n59395), .O(n16648[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_11 (.CI(n59395), .I0(n17259[8]), .I1(n749_adj_5541), 
            .CO(n59396));
    SB_LUT4 add_6361_10_lut (.I0(GND_net), .I1(n17259[7]), .I2(n676_adj_5540), 
            .I3(n59394), .O(n16648[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_10 (.CI(n59394), .I0(n17259[7]), .I1(n676_adj_5540), 
            .CO(n59395));
    SB_LUT4 add_6361_9_lut (.I0(GND_net), .I1(n17259[6]), .I2(n603_adj_5539), 
            .I3(n59393), .O(n16648[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_9 (.CI(n59393), .I0(n17259[6]), .I1(n603_adj_5539), 
            .CO(n59394));
    SB_LUT4 add_6542_6_lut (.I0(GND_net), .I1(n19778[3]), .I2(n402_adj_5538), 
            .I3(n60342), .O(n19540[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_21 (.CI(n58926), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n58927));
    SB_LUT4 sub_15_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n58925), .O(n207[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[21]), 
            .I3(n59097), .O(n48[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_23 (.CI(n59097), .I0(GND_net), .I1(n1_adj_5701[21]), 
            .CO(n59098));
    SB_LUT4 mult_24_i706_2_lut (.I0(\Ki[14] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_5575));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6361_8_lut (.I0(GND_net), .I1(n17259[5]), .I2(n530_adj_5531), 
            .I3(n59392), .O(n16648[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_8 (.CI(n59392), .I0(n17259[5]), .I1(n530_adj_5531), 
            .CO(n59393));
    SB_CARRY add_6542_6 (.CI(n60342), .I0(n19778[3]), .I1(n402_adj_5538), 
            .CO(n60343));
    SB_LUT4 add_6361_7_lut (.I0(GND_net), .I1(n17259[4]), .I2(n457_adj_5529), 
            .I3(n59391), .O(n16648[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i81_2_lut (.I0(\Kp[1] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_5574));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i81_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6361_7 (.CI(n59391), .I0(n17259[4]), .I1(n457_adj_5529), 
            .CO(n59392));
    SB_LUT4 mult_23_i34_2_lut (.I0(\Kp[0] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_5573));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6361_6_lut (.I0(GND_net), .I1(n17259[3]), .I2(n384_adj_5528), 
            .I3(n59390), .O(n16648[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_20 (.CI(n58925), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n58926));
    SB_LUT4 sub_15_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n58924), .O(n207[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[20]), 
            .I3(n59096), .O(n48[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_6 (.CI(n59390), .I0(n17259[3]), .I1(n384_adj_5528), 
            .CO(n59391));
    SB_LUT4 add_6361_5_lut (.I0(GND_net), .I1(n17259[2]), .I2(n311_adj_5519), 
            .I3(n59389), .O(n16648[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i471_2_lut (.I0(\Ki[9] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_5572));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i130_2_lut (.I0(\Kp[2] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_5571));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6361_5 (.CI(n59389), .I0(n17259[2]), .I1(n311_adj_5519), 
            .CO(n59390));
    SB_CARRY unary_minus_27_add_3_22 (.CI(n59096), .I0(GND_net), .I1(n1_adj_5701[20]), 
            .CO(n59097));
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[19]), 
            .I3(n59095), .O(n486)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6361_4_lut (.I0(GND_net), .I1(n17259[1]), .I2(n238_adj_5511), 
            .I3(n59388), .O(n16648[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_21 (.CI(n59095), .I0(GND_net), .I1(n1_adj_5701[19]), 
            .CO(n59096));
    SB_CARRY add_6361_4 (.CI(n59388), .I0(n17259[1]), .I1(n238_adj_5511), 
            .CO(n59389));
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[18]), 
            .I3(n59094), .O(n48[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_20 (.CI(n59094), .I0(GND_net), .I1(n1_adj_5701[18]), 
            .CO(n59095));
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[17]), 
            .I3(n59093), .O(n48[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6361_3_lut (.I0(GND_net), .I1(n17259[0]), .I2(n165_adj_5508), 
            .I3(n59387), .O(n16648[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_3 (.CI(n59387), .I0(n17259[0]), .I1(n165_adj_5508), 
            .CO(n59388));
    SB_LUT4 add_6361_2_lut (.I0(GND_net), .I1(n23_adj_5507), .I2(n92_adj_5506), 
            .I3(GND_net), .O(n16648[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_19 (.CI(n59093), .I0(GND_net), .I1(n1_adj_5701[17]), 
            .CO(n59094));
    SB_CARRY add_6361_2 (.CI(GND_net), .I0(n23_adj_5507), .I1(n92_adj_5506), 
            .CO(n59387));
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[16]), 
            .I3(n59092), .O(n48[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_18 (.CI(n59092), .I0(GND_net), .I1(n1_adj_5701[16]), 
            .CO(n59093));
    SB_LUT4 add_6542_5_lut (.I0(GND_net), .I1(n19778[2]), .I2(n329_adj_5504), 
            .I3(n60341), .O(n19540[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_19 (.CI(n58924), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n58925));
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[15]), 
            .I3(n59091), .O(n48[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i179_2_lut (.I0(\Kp[3] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_5569));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i228_2_lut (.I0(\Kp[4] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_5567));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_27_add_3_17 (.CI(n59091), .I0(GND_net), .I1(n1_adj_5701[15]), 
            .CO(n59092));
    SB_LUT4 mult_23_i277_2_lut (.I0(\Kp[5] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_5563));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[14]), 
            .I3(n59090), .O(n48[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_16 (.CI(n59090), .I0(GND_net), .I1(n1_adj_5701[14]), 
            .CO(n59091));
    SB_LUT4 mult_23_i326_2_lut (.I0(\Kp[6] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_5559));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[13]), 
            .I3(n59089), .O(n48[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_5 (.CI(n60341), .I0(n19778[2]), .I1(n329_adj_5504), 
            .CO(n60342));
    SB_CARRY unary_minus_27_add_3_15 (.CI(n59089), .I0(GND_net), .I1(n1_adj_5701[13]), 
            .CO(n59090));
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[12]), 
            .I3(n59088), .O(n48[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n59088), .I0(GND_net), .I1(n1_adj_5701[12]), 
            .CO(n59089));
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i375_2_lut (.I0(\Kp[7] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i424_2_lut (.I0(\Kp[8] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i67_2_lut (.I0(\Ki[1] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_5556));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[11]), 
            .I3(n59087), .O(n48[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_13 (.CI(n59087), .I0(GND_net), .I1(n1_adj_5701[11]), 
            .CO(n59088));
    SB_LUT4 add_6542_4_lut (.I0(GND_net), .I1(n19778[1]), .I2(n256_adj_5496), 
            .I3(n60340), .O(n19540[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i20_2_lut (.I0(\Ki[0] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5555));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i116_2_lut (.I0(\Ki[2] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_5554));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6542_4 (.CI(n60340), .I0(n19778[1]), .I1(n256_adj_5496), 
            .CO(n60341));
    SB_LUT4 add_6542_3_lut (.I0(GND_net), .I1(n19778[0]), .I2(n183_adj_5490), 
            .I3(n60339), .O(n19540[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_3 (.CI(n60339), .I0(n19778[0]), .I1(n183_adj_5490), 
            .CO(n60340));
    SB_LUT4 add_6542_2_lut (.I0(GND_net), .I1(n41_adj_5488), .I2(n110), 
            .I3(GND_net), .O(n19540[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_2 (.CI(GND_net), .I0(n41_adj_5488), .I1(n110), .CO(n60339));
    SB_LUT4 add_6394_17_lut (.I0(GND_net), .I1(n17802[14]), .I2(GND_net), 
            .I3(n59369), .O(n17259[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6614_7_lut (.I0(GND_net), .I1(n69227), .I2(n490_adj_5429), 
            .I3(n60338), .O(n20289[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_16_lut (.I0(GND_net), .I1(n17802[13]), .I2(n1117_adj_5425), 
            .I3(n59368), .O(n17259[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i312_2_lut (.I0(\Ki[6] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_5537));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6394_16 (.CI(n59368), .I0(n17802[13]), .I1(n1117_adj_5425), 
            .CO(n59369));
    SB_LUT4 add_6394_15_lut (.I0(GND_net), .I1(n17802[12]), .I2(n1044), 
            .I3(n59367), .O(n17259[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_15 (.CI(n59367), .I0(n17802[12]), .I1(n1044), .CO(n59368));
    SB_LUT4 add_6394_14_lut (.I0(GND_net), .I1(n17802[11]), .I2(n971), 
            .I3(n59366), .O(n17259[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i57_2_lut (.I0(\Kp[1] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_5536));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6614_6_lut (.I0(GND_net), .I1(n20372[3]), .I2(n417_adj_5422), 
            .I3(n60337), .O(n20289[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6614_6 (.CI(n60337), .I0(n20372[3]), .I1(n417_adj_5422), 
            .CO(n60338));
    SB_LUT4 add_6614_5_lut (.I0(GND_net), .I1(n20372[2]), .I2(n344_adj_5419), 
            .I3(n60336), .O(n20289[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6614_5 (.CI(n60336), .I0(n20372[2]), .I1(n344_adj_5419), 
            .CO(n60337));
    SB_LUT4 mult_23_i10_2_lut (.I0(\Kp[0] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_5535));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6614_4_lut (.I0(GND_net), .I1(n20372[1]), .I2(n271_adj_5415), 
            .I3(n60335), .O(n20289[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[10]), 
            .I3(n59086), .O(n48[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_14 (.CI(n59366), .I0(n17802[11]), .I1(n971), .CO(n59367));
    SB_LUT4 mult_24_i165_2_lut (.I0(\Ki[3] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_5552));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i165_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6614_4 (.CI(n60335), .I0(n20372[1]), .I1(n271_adj_5415), 
            .CO(n60336));
    SB_LUT4 add_6614_3_lut (.I0(GND_net), .I1(n20372[0]), .I2(n198_adj_5413), 
            .I3(n60334), .O(n20289[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_13_lut (.I0(GND_net), .I1(n17802[10]), .I2(n898), 
            .I3(n59365), .O(n17259[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n58923), .O(n207[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_13 (.CI(n59365), .I0(n17802[10]), .I1(n898), .CO(n59366));
    SB_CARRY sub_15_add_2_18 (.CI(n58923), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n58924));
    SB_LUT4 sub_15_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n58922), .O(n207[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_12_lut (.I0(GND_net), .I1(n17802[9]), .I2(n825), 
            .I3(n59364), .O(n17259[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_17 (.CI(n58922), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n58923));
    SB_LUT4 sub_15_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n58921), .O(n207[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_12 (.CI(n59364), .I0(n17802[9]), .I1(n825), .CO(n59365));
    SB_CARRY sub_15_add_2_16 (.CI(n58921), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n58922));
    SB_LUT4 sub_15_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n58920), .O(n207[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_11_lut (.I0(GND_net), .I1(n17802[8]), .I2(n752), 
            .I3(n59363), .O(n17259[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_15 (.CI(n58920), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n58921));
    SB_LUT4 sub_15_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(n10_adj_33), 
            .I3(n58919), .O(n207[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_11 (.CI(n59363), .I0(n17802[8]), .I1(n752), .CO(n59364));
    SB_CARRY add_6614_3 (.CI(n60334), .I0(n20372[0]), .I1(n198_adj_5413), 
            .CO(n60335));
    SB_CARRY unary_minus_27_add_3_12 (.CI(n59086), .I0(GND_net), .I1(n1_adj_5701[10]), 
            .CO(n59087));
    SB_LUT4 add_6614_2_lut (.I0(GND_net), .I1(n56_adj_5411), .I2(n125_adj_5410), 
            .I3(GND_net), .O(n20289[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6614_2 (.CI(GND_net), .I0(n56_adj_5411), .I1(n125_adj_5410), 
            .CO(n60334));
    SB_LUT4 mult_23_i106_2_lut (.I0(\Kp[2] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_5533));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i106_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_14 (.CI(n58919), .I0(setpoint[12]), .I1(n10_adj_33), 
            .CO(n58920));
    SB_LUT4 sub_15_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(n42994), 
            .I3(n58918), .O(n207[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_10_lut (.I0(GND_net), .I1(n17802[7]), .I2(n679), 
            .I3(n59362), .O(n17259[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[9]), 
            .I3(n59085), .O(n48[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_13 (.CI(n58918), .I0(setpoint[11]), .I1(n42994), 
            .CO(n58919));
    SB_LUT4 sub_15_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n58917), .O(n207[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_10 (.CI(n59362), .I0(n17802[7]), .I1(n679), .CO(n59363));
    SB_CARRY unary_minus_27_add_3_11 (.CI(n59085), .I0(GND_net), .I1(n1_adj_5701[9]), 
            .CO(n59086));
    SB_LUT4 add_6394_9_lut (.I0(GND_net), .I1(n17802[6]), .I2(n606), .I3(n59361), 
            .O(n17259[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_9 (.CI(n59361), .I0(n17802[6]), .I1(n606), .CO(n59362));
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[8]), 
            .I3(n59084), .O(n48[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_10 (.CI(n59084), .I0(GND_net), .I1(n1_adj_5701[8]), 
            .CO(n59085));
    SB_LUT4 mult_24_i214_2_lut (.I0(\Ki[4] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_5547));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6394_8_lut (.I0(GND_net), .I1(n17802[5]), .I2(n533), .I3(n59360), 
            .O(n17259[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_8 (.CI(n59360), .I0(n17802[5]), .I1(n533), .CO(n59361));
    SB_LUT4 add_6394_7_lut (.I0(GND_net), .I1(n17802[4]), .I2(n460_adj_5404), 
            .I3(n59359), .O(n17259[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i263_2_lut (.I0(\Ki[5] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_5545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6394_7 (.CI(n59359), .I0(n17802[4]), .I1(n460_adj_5404), 
            .CO(n59360));
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[7]), 
            .I3(n59083), .O(n48[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_6_lut (.I0(GND_net), .I1(n17802[3]), .I2(n387_adj_5402), 
            .I3(n59358), .O(n17259[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_6 (.CI(n59358), .I0(n17802[3]), .I1(n387_adj_5402), 
            .CO(n59359));
    SB_LUT4 add_6394_5_lut (.I0(GND_net), .I1(n17802[2]), .I2(n314_adj_5401), 
            .I3(n59357), .O(n17259[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_5 (.CI(n59357), .I0(n17802[2]), .I1(n314_adj_5401), 
            .CO(n59358));
    SB_LUT4 add_6394_4_lut (.I0(GND_net), .I1(n17802[1]), .I2(n241_adj_5400), 
            .I3(n59356), .O(n17259[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_4 (.CI(n59356), .I0(n17802[1]), .I1(n241_adj_5400), 
            .CO(n59357));
    SB_LUT4 add_6394_3_lut (.I0(GND_net), .I1(n17802[0]), .I2(n168), .I3(n59355), 
            .O(n17259[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_3 (.CI(n59355), .I0(n17802[0]), .I1(n168), .CO(n59356));
    SB_LUT4 add_6394_2_lut (.I0(GND_net), .I1(n26_adj_5398), .I2(n95), 
            .I3(GND_net), .O(n17259[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i155_2_lut (.I0(\Kp[3] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_5532));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i155_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6394_2 (.CI(GND_net), .I0(n26_adj_5398), .I1(n95), .CO(n59355));
    SB_LUT4 mult_23_i204_2_lut (.I0(\Kp[4] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_5530));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i253_2_lut (.I0(\Kp[5] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_5527));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i361_2_lut (.I0(\Ki[7] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_5526));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i410_2_lut (.I0(\Ki[8] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_5525));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i302_2_lut (.I0(\Kp[6] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_5524));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i351_2_lut (.I0(\Kp[7] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_5523));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i400_2_lut (.I0(\Kp[8] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_5522));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n79534_bdd_4_lut (.I0(n79534), .I1(n535[23]), .I2(n455[23]), 
            .I3(n4736), .O(n79537));
    defparam n79534_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i449_2_lut (.I0(\Kp[9] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_5521));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i449_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_12 (.CI(n58917), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n58918));
    SB_LUT4 mult_23_i498_2_lut (.I0(\Kp[10] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_5518));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i547_2_lut (.I0(\Kp[11] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_5517));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i596_2_lut (.I0(\Kp[12] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_5516));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i596_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_27_add_3_9 (.CI(n59083), .I0(GND_net), .I1(n1_adj_5701[7]), 
            .CO(n59084));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[6]), 
            .I3(n59082), .O(n48[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i645_2_lut (.I0(\Kp[13] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_5514));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i694_2_lut (.I0(\Kp[14] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_5513));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i743_2_lut (.I0(\Kp[15] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_5512));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i743_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_27_add_3_8 (.CI(n59082), .I0(GND_net), .I1(n1_adj_5701[6]), 
            .CO(n59083));
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[5]), 
            .I3(n59081), .O(n48[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_7 (.CI(n59081), .I0(GND_net), .I1(n1_adj_5701[5]), 
            .CO(n59082));
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[4]), 
            .I3(n59080), .O(n48[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_6 (.CI(n59080), .I0(GND_net), .I1(n1_adj_5701[4]), 
            .CO(n59081));
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[3]), 
            .I3(n59079), .O(n48[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n59079), .I0(GND_net), .I1(n1_adj_5701[3]), 
            .CO(n59080));
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[2]), 
            .I3(n59078), .O(n48[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i44713_2_lut_3_lut_4_lut (.I0(\Ki[1] ), .I1(n339), .I2(\Ki[0] ), 
            .I3(n37117), .O(n58789));   // verilog/motorControl.v(61[29:40])
    defparam i44713_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i44711_2_lut_3_lut_4_lut (.I0(\Ki[1] ), .I1(n339), .I2(\Ki[0] ), 
            .I3(n37117), .O(n20492[0]));   // verilog/motorControl.v(61[29:40])
    defparam i44711_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_6610_8_lut (.I0(GND_net), .I1(n20350[5]), .I2(n560), .I3(n59338), 
            .O(n20256[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6610_7_lut (.I0(GND_net), .I1(n20350[4]), .I2(n487), .I3(n59337), 
            .O(n20256[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6610_7 (.CI(n59337), .I0(n20350[4]), .I1(n487), .CO(n59338));
    SB_LUT4 add_6610_6_lut (.I0(GND_net), .I1(n20350[3]), .I2(n414), .I3(n59336), 
            .O(n20256[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_4 (.CI(n59078), .I0(GND_net), .I1(n1_adj_5701[2]), 
            .CO(n59079));
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5701[1]), 
            .I3(n59077), .O(n48[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6610_6 (.CI(n59336), .I0(n20350[3]), .I1(n414), .CO(n59337));
    SB_LUT4 add_6610_5_lut (.I0(GND_net), .I1(n20350[2]), .I2(n341), .I3(n59335), 
            .O(n20256[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6610_5 (.CI(n59335), .I0(n20350[2]), .I1(n341), .CO(n59336));
    SB_LUT4 add_6610_4_lut (.I0(GND_net), .I1(n20350[1]), .I2(n268), .I3(n59334), 
            .O(n20256[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n59077), .I0(GND_net), .I1(n1_adj_5701[1]), 
            .CO(n59078));
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(n45309), .I1(GND_net), .I2(n1_adj_5701[0]), 
            .I3(VCC_net), .O(n75139)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_6610_4 (.CI(n59334), .I0(n20350[1]), .I1(n268), .CO(n59335));
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5701[0]), 
            .CO(n59077));
    SB_LUT4 i1_3_lut_4_lut (.I0(\Ki[2] ), .I1(n339), .I2(n58789), .I3(n20501[0]), 
            .O(n20492[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 add_6610_3_lut (.I0(GND_net), .I1(n20350[0]), .I2(n195), .I3(n59333), 
            .O(n20256[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6610_3 (.CI(n59333), .I0(n20350[0]), .I1(n195), .CO(n59334));
    SB_LUT4 add_6610_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n20256[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6610_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n59333));
    SB_LUT4 i44724_3_lut_4_lut (.I0(\Ki[2] ), .I1(n339), .I2(n58789), 
            .I3(n20501[0]), .O(n4_adj_5291));   // verilog/motorControl.v(61[29:40])
    defparam i44724_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_6425_16_lut (.I0(GND_net), .I1(n18281[13]), .I2(n1120), 
            .I3(n59332), .O(n17802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6425_15_lut (.I0(GND_net), .I1(n18281[12]), .I2(n1047), 
            .I3(n59331), .O(n17802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_15 (.CI(n59331), .I0(n18281[12]), .I1(n1047), .CO(n59332));
    SB_LUT4 add_6425_14_lut (.I0(GND_net), .I1(n18281[11]), .I2(n974), 
            .I3(n59330), .O(n17802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_14 (.CI(n59330), .I0(n18281[11]), .I1(n974), .CO(n59331));
    SB_LUT4 add_6425_13_lut (.I0(GND_net), .I1(n18281[10]), .I2(n901), 
            .I3(n59329), .O(n17802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_13 (.CI(n59329), .I0(n18281[10]), .I1(n901), .CO(n59330));
    SB_LUT4 add_6425_12_lut (.I0(GND_net), .I1(n18281[9]), .I2(n828), 
            .I3(n59328), .O(n17802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_12 (.CI(n59328), .I0(n18281[9]), .I1(n828), .CO(n59329));
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(n11922[0]), .I2(n12498[0]), 
            .I3(n58976), .O(n455[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6425_11_lut (.I0(GND_net), .I1(n18281[8]), .I2(n755), 
            .I3(n59327), .O(n17802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_11 (.CI(n59327), .I0(n18281[8]), .I1(n755), .CO(n59328));
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(n360[22]), .I2(n46[22]), 
            .I3(n58975), .O(n455[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6425_10_lut (.I0(GND_net), .I1(n18281[7]), .I2(n682), 
            .I3(n59326), .O(n17802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_10 (.CI(n59326), .I0(n18281[7]), .I1(n682), .CO(n59327));
    SB_CARRY add_25_24 (.CI(n58975), .I0(n360[22]), .I1(n46[22]), .CO(n58976));
    SB_LUT4 add_6425_9_lut (.I0(GND_net), .I1(n18281[6]), .I2(n609), .I3(n59325), 
            .O(n17802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_9 (.CI(n59325), .I0(n18281[6]), .I1(n609), .CO(n59326));
    SB_LUT4 add_6425_8_lut (.I0(GND_net), .I1(n18281[5]), .I2(n536_adj_5326), 
            .I3(n59324), .O(n17802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_8 (.CI(n59324), .I0(n18281[5]), .I1(n536_adj_5326), 
            .CO(n59325));
    SB_LUT4 add_6425_7_lut (.I0(GND_net), .I1(n18281[4]), .I2(n463_adj_5324), 
            .I3(n59323), .O(n17802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_7 (.CI(n59323), .I0(n18281[4]), .I1(n463_adj_5324), 
            .CO(n59324));
    SB_LUT4 add_6425_6_lut (.I0(GND_net), .I1(n18281[3]), .I2(n390_adj_5323), 
            .I3(n59322), .O(n17802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_6 (.CI(n59322), .I0(n18281[3]), .I1(n390_adj_5323), 
            .CO(n59323));
    SB_LUT4 add_6425_5_lut (.I0(GND_net), .I1(n18281[2]), .I2(n317), .I3(n59321), 
            .O(n17802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_5 (.CI(n59321), .I0(n18281[2]), .I1(n317), .CO(n59322));
    SB_LUT4 add_6425_4_lut (.I0(GND_net), .I1(n18281[1]), .I2(n244_adj_5318), 
            .I3(n59320), .O(n17802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_4 (.CI(n59320), .I0(n18281[1]), .I1(n244_adj_5318), 
            .CO(n59321));
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(n360[21]), .I2(n46[21]), 
            .I3(n58974), .O(n455[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6425_3_lut (.I0(GND_net), .I1(n18281[0]), .I2(n171), .I3(n59319), 
            .O(n17802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_3 (.CI(n59319), .I0(n18281[0]), .I1(n171), .CO(n59320));
    SB_CARRY add_25_23 (.CI(n58974), .I0(n360[21]), .I1(n46[21]), .CO(n58975));
    SB_LUT4 add_6425_2_lut (.I0(GND_net), .I1(n29_adj_5317), .I2(n98), 
            .I3(GND_net), .O(n17802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_2 (.CI(GND_net), .I0(n29_adj_5317), .I1(n98), .CO(n59319));
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(n360[20]), .I2(n46[20]), 
            .I3(n58973), .O(n455[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_22 (.CI(n58973), .I0(n360[20]), .I1(n46[20]), .CO(n58974));
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(n360[19]), .I2(n46[19]), 
            .I3(n58972), .O(n460)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_21 (.CI(n58972), .I0(n360[19]), .I1(n46[19]), .CO(n58973));
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(n360[18]), .I2(n46[18]), 
            .I3(n58971), .O(n461)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_20 (.CI(n58971), .I0(n360[18]), .I1(n46[18]), .CO(n58972));
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(n360[17]), .I2(n46[17]), 
            .I3(n58970), .O(n462)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_19 (.CI(n58970), .I0(n360[17]), .I1(n46[17]), .CO(n58971));
    SB_LUT4 mult_24_i459_2_lut (.I0(\Ki[9] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_5502));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(n360[16]), .I2(n46[16]), 
            .I3(n58969), .O(n455[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_18 (.CI(n58969), .I0(n360[16]), .I1(n46[16]), .CO(n58970));
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(n360[15]), .I2(n46[15]), 
            .I3(n58968), .O(n455[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n59076), .O(n285[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_17 (.CI(n58968), .I0(n360[15]), .I1(n46[15]), .CO(n58969));
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n59075), .O(n285[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_15_lut (.I0(GND_net), .I1(n18700[12]), .I2(n1050), 
            .I3(n59303), .O(n18281[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n59075), .I0(GND_net), .I1(n1[22]), 
            .CO(n59076));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n59074), .O(n285[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(n360[14]), .I2(n46[14]), 
            .I3(n58967), .O(n455[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_16 (.CI(n58967), .I0(n360[14]), .I1(n46[14]), .CO(n58968));
    SB_CARRY unary_minus_20_add_3_23 (.CI(n59074), .I0(GND_net), .I1(n1[21]), 
            .CO(n59075));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n59073), .O(n285[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_14_lut (.I0(GND_net), .I1(n18700[11]), .I2(n977), 
            .I3(n59302), .O(n18281[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n59073), .I0(GND_net), .I1(n1[20]), 
            .CO(n59074));
    SB_CARRY add_6454_14 (.CI(n59302), .I0(n18700[11]), .I1(n977), .CO(n59303));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n59072), .O(n285[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n59072), .I0(GND_net), .I1(n1[19]), 
            .CO(n59073));
    SB_LUT4 mult_23_i267_2_lut (.I0(\Kp[5] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(n360[13]), .I2(n46[13]), 
            .I3(n58966), .O(n455[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_15 (.CI(n58966), .I0(n360[13]), .I1(n46[13]), .CO(n58967));
    SB_LUT4 add_6454_13_lut (.I0(GND_net), .I1(n18700[10]), .I2(n904), 
            .I3(n59301), .O(n18281[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_13 (.CI(n59301), .I0(n18700[10]), .I1(n904), .CO(n59302));
    SB_LUT4 add_6454_12_lut (.I0(GND_net), .I1(n18700[9]), .I2(n831), 
            .I3(n59300), .O(n18281[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_12 (.CI(n59300), .I0(n18700[9]), .I1(n831), .CO(n59301));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n59071), .O(n291)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_20 (.CI(n59071), .I0(GND_net), .I1(n1[18]), 
            .CO(n59072));
    SB_LUT4 add_6454_11_lut (.I0(GND_net), .I1(n18700[8]), .I2(n758), 
            .I3(n59299), .O(n18281[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n59070), .O(n285[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(n360[12]), .I2(n46[12]), 
            .I3(n58965), .O(n467)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n59070), .I0(GND_net), .I1(n1[17]), 
            .CO(n59071));
    SB_CARRY add_25_14 (.CI(n58965), .I0(n360[12]), .I1(n46[12]), .CO(n58966));
    SB_CARRY add_6454_11 (.CI(n59299), .I0(n18700[8]), .I1(n758), .CO(n59300));
    SB_LUT4 add_6454_10_lut (.I0(GND_net), .I1(n18700[7]), .I2(n685), 
            .I3(n59298), .O(n18281[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_10 (.CI(n59298), .I0(n18700[7]), .I1(n685), .CO(n59299));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n59069), .O(n285[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n59069), .I0(GND_net), .I1(n1[16]), 
            .CO(n59070));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n59068), .O(n285[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_9_lut (.I0(GND_net), .I1(n18700[6]), .I2(n612), .I3(n59297), 
            .O(n18281[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_9 (.CI(n59297), .I0(n18700[6]), .I1(n612), .CO(n59298));
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(n360[11]), .I2(n46[11]), 
            .I3(n58964), .O(n455[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_8_lut (.I0(GND_net), .I1(n18700[5]), .I2(n539_adj_5301), 
            .I3(n59296), .O(n18281[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_8 (.CI(n59296), .I0(n18700[5]), .I1(n539_adj_5301), 
            .CO(n59297));
    SB_CARRY add_25_13 (.CI(n58964), .I0(n360[11]), .I1(n46[11]), .CO(n58965));
    SB_LUT4 add_6454_7_lut (.I0(GND_net), .I1(n18700[4]), .I2(n466_adj_5300), 
            .I3(n59295), .O(n18281[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i44622_2_lut_3_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n62_adj_5427), 
            .I3(GND_net), .O(n20372[0]));   // verilog/motorControl.v(61[20:26])
    defparam i44622_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_CARRY add_6454_7 (.CI(n59295), .I0(n18700[4]), .I1(n466_adj_5300), 
            .CO(n59296));
    SB_LUT4 add_6454_6_lut (.I0(GND_net), .I1(n18700[3]), .I2(n393), .I3(n59294), 
            .O(n18281[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(n360[10]), .I2(n46[10]), 
            .I3(n58963), .O(n455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_6 (.CI(n59294), .I0(n18700[3]), .I1(n393), .CO(n59295));
    SB_LUT4 add_6454_5_lut (.I0(GND_net), .I1(n18700[2]), .I2(n320), .I3(n59293), 
            .O(n18281[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_5 (.CI(n59293), .I0(n18700[2]), .I1(n320), .CO(n59294));
    SB_LUT4 add_6454_4_lut (.I0(GND_net), .I1(n18700[1]), .I2(n247_adj_5296), 
            .I3(n59292), .O(n18281[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_4 (.CI(n59292), .I0(n18700[1]), .I1(n247_adj_5296), 
            .CO(n59293));
    SB_LUT4 mult_24_i508_2_lut (.I0(\Ki[10] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_5498));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6454_3_lut (.I0(GND_net), .I1(n18700[0]), .I2(n174), .I3(n59291), 
            .O(n18281[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_3 (.CI(n59291), .I0(n18700[0]), .I1(n174), .CO(n59292));
    SB_LUT4 add_6454_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n18281[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n59291));
    SB_CARRY add_25_12 (.CI(n58963), .I0(n360[10]), .I1(n46[10]), .CO(n58964));
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(n360[9]), .I2(n46[9]), .I3(n58962), 
            .O(n455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_11 (.CI(n58962), .I0(n360[9]), .I1(n46[9]), .CO(n58963));
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(n360[8]), .I2(n46[8]), .I3(n58961), 
            .O(n455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_10 (.CI(n58961), .I0(n360[8]), .I1(n46[8]), .CO(n58962));
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(n360[7]), .I2(n46[7]), .I3(n58960), 
            .O(n455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i557_2_lut (.I0(\Ki[11] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_5495));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1802 (.I0(\Kp[1] ), .I1(n207[22]), .I2(n62_adj_5427), 
            .I3(n71550), .O(n20372[1]));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_4_lut_adj_1802.LUT_INIT = 16'h7f80;
    SB_CARRY add_25_9 (.CI(n58960), .I0(n360[7]), .I1(n46[7]), .CO(n58961));
    SB_CARRY unary_minus_20_add_3_17 (.CI(n59068), .I0(GND_net), .I1(n1[15]), 
            .CO(n59069));
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(n360[6]), .I2(n46[6]), .I3(n58959), 
            .O(n455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n59067), .O(n285[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i316_2_lut (.I0(\Kp[6] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i55_2_lut (.I0(\Kp[1] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_5494));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i8_2_lut (.I0(\Kp[0] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5493));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i8_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_25_8 (.CI(n58959), .I0(n360[6]), .I1(n46[6]), .CO(n58960));
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(n360[5]), .I2(n46[5]), .I3(n58958), 
            .O(n455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_7 (.CI(n58958), .I0(n360[5]), .I1(n46[5]), .CO(n58959));
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(n360[4]), .I2(n46[4]), .I3(n58957), 
            .O(n475)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6622_7_lut (.I0(GND_net), .I1(n69694), .I2(n490), .I3(n59276), 
            .O(n20350[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6622_6_lut (.I0(GND_net), .I1(n20418[3]), .I2(n417), .I3(n59275), 
            .O(n20350[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i104_2_lut (.I0(\Kp[2] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_5492));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i153_2_lut (.I0(\Kp[3] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_5491));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i73_2_lut (.I0(\Kp[1] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i26_2_lut (.I0(\Kp[0] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_5487));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i202_2_lut (.I0(\Kp[4] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_5486));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i122_2_lut (.I0(\Kp[2] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i251_2_lut (.I0(\Kp[5] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_5485));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i171_2_lut (.I0(\Kp[3] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_5484));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i300_2_lut (.I0(\Kp[6] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_5483));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i220_2_lut (.I0(\Kp[4] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i349_2_lut (.I0(\Kp[7] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_5482));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i606_2_lut (.I0(\Ki[12] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_5481));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i655_2_lut (.I0(\Ki[13] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_5480));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i269_2_lut (.I0(\Kp[5] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_5479));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i398_2_lut (.I0(\Kp[8] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_5478));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i318_2_lut (.I0(\Kp[6] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_5477));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i447_2_lut (.I0(\Kp[9] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_5476));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i367_2_lut (.I0(\Kp[7] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_5475));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i496_2_lut (.I0(\Kp[10] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_5474));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i416_2_lut (.I0(\Kp[8] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i545_2_lut (.I0(\Kp[11] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_5473));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i594_2_lut (.I0(\Kp[12] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_5472));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i704_2_lut (.I0(\Ki[14] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_5471));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i753_2_lut (.I0(\Ki[15] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_5470));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i643_2_lut (.I0(\Kp[13] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_5469));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i692_2_lut (.I0(\Kp[14] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_5468));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i65_2_lut (.I0(\Ki[1] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_5466));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i18_2_lut (.I0(\Ki[0] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_5465));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i741_2_lut (.I0(\Kp[15] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_5464));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i465_2_lut (.I0(\Kp[9] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i365_2_lut (.I0(\Kp[7] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i514_2_lut (.I0(\Kp[10] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i563_2_lut (.I0(\Kp[11] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i612_2_lut (.I0(\Kp[12] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i414_2_lut (.I0(\Kp[8] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i114_2_lut (.I0(\Ki[2] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_5463));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i463_2_lut (.I0(\Kp[9] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i53_2_lut (.I0(\Kp[1] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_5462));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i6_2_lut (.I0(\Kp[0] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5461));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i102_2_lut (.I0(\Kp[2] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_5460));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i151_2_lut (.I0(\Kp[3] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_5459));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i200_2_lut (.I0(\Kp[4] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_5458));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i163_2_lut (.I0(\Ki[3] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_5457));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i249_2_lut (.I0(\Kp[5] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_5456));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i298_2_lut (.I0(\Kp[6] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_5455));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i347_2_lut (.I0(\Kp[7] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_5454));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i396_2_lut (.I0(\Kp[8] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_5453));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i445_2_lut (.I0(\Kp[9] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_5452));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i494_2_lut (.I0(\Kp[10] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_5451));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i543_2_lut (.I0(\Kp[11] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_5450));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i512_2_lut (.I0(\Kp[10] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i561_2_lut (.I0(\Kp[11] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i592_2_lut (.I0(\Kp[12] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_5448));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60100_3_lut_4_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(n233[2]), .O(n75956));   // verilog/motorControl.v(58[23:46])
    defparam i60100_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n11882_bdd_4_lut_63393 (.I0(n11882), .I1(n75258), .I2(setpoint[5]), 
            .I3(n4736), .O(n79276));
    defparam n11882_bdd_4_lut_63393.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(GND_net), .O(n6_adj_5235));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_23_i641_2_lut (.I0(\Kp[13] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_5446));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i690_2_lut (.I0(\Kp[14] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_5445));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i739_2_lut (.I0(\Kp[15] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_5444));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n233[3]), 
            .I2(n233[2]), .I3(GND_net), .O(n6_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i60168_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n233[3]), .I2(n233[2]), 
            .I3(IntegralLimit[2]), .O(n76024));   // verilog/motorControl.v(56[14:36])
    defparam i60168_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n79276_bdd_4_lut (.I0(n79276), .I1(n535[5]), .I2(n455[5]), 
            .I3(n4736), .O(n79279));
    defparam n79276_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_9_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), 
            .I2(setpoint[2]), .I3(GND_net), .O(n6_adj_5227));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i60332_3_lut_4_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), .I2(setpoint[2]), 
            .I3(PWMLimit[2]), .O(n76188));   // verilog/motorControl.v(45[16:33])
    defparam i60332_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i60260_3_lut_4_lut (.I0(setpoint[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(setpoint[2]), .O(n76116));   // verilog/motorControl.v(47[25:43])
    defparam i60260_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(setpoint[3]), .I1(n535[3]), 
            .I2(n535[2]), .I3(GND_net), .O(n6_adj_5281));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 n11882_bdd_4_lut_63601 (.I0(n11882), .I1(n75294), .I2(setpoint[22]), 
            .I3(n4736), .O(n79498));
    defparam n11882_bdd_4_lut_63601.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i212_2_lut (.I0(\Ki[4] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_5442));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59638_2_lut (.I0(PWMLimit[7]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75260));
    defparam i59638_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i8_3_lut (.I0(n233[7]), .I1(n285[7]), .I2(n284), .I3(GND_net), 
            .O(n310[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i8_3_lut (.I0(n310[7]), .I1(IntegralLimit[7]), .I2(n258), 
            .I3(GND_net), .O(n352));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i63_2_lut (.I0(\Ki[1] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i16_2_lut (.I0(\Ki[0] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5399));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i112_2_lut (.I0(\Ki[2] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i261_2_lut (.I0(\Ki[5] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_5441));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i161_2_lut (.I0(\Ki[3] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_5396));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i420_2_lut (.I0(\Ki[8] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_5395));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i210_2_lut (.I0(\Ki[4] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_5392));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i259_2_lut (.I0(\Ki[5] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_5391));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i469_2_lut (.I0(\Ki[9] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_5390));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i14_3_lut (.I0(n233[13]), .I1(n285[13]), .I2(n284), 
            .I3(GND_net), .O(n310[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i14_3_lut (.I0(n310[13]), .I1(IntegralLimit[13]), .I2(n258), 
            .I3(GND_net), .O(n346));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i518_2_lut (.I0(\Ki[10] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_5389));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i308_2_lut (.I0(\Ki[6] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_5388));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i6_3_lut_3_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(GND_net), .O(n6_adj_5428));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_24_i357_2_lut (.I0(\Ki[7] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i51_2_lut (.I0(\Kp[1] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_5381));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i4_2_lut (.I0(\Kp[0] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5380));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i100_2_lut (.I0(\Kp[2] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_5379));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n79498_bdd_4_lut (.I0(n79498), .I1(n535[22]), .I2(n455[22]), 
            .I3(n4736), .O(n79501));
    defparam n79498_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i406_2_lut (.I0(\Ki[8] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i310_2_lut (.I0(\Ki[6] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_5440));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i455_2_lut (.I0(\Ki[9] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i504_2_lut (.I0(\Ki[10] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i553_2_lut (.I0(\Ki[11] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59808_3_lut_4_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(n455[2]), .O(n75664));   // verilog/motorControl.v(65[25:41])
    defparam i59808_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i602_2_lut (.I0(\Ki[12] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i651_2_lut (.I0(\Ki[13] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i359_2_lut (.I0(\Ki[7] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_5439));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i408_2_lut (.I0(\Ki[8] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_5438));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i457_2_lut (.I0(\Ki[9] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_5437));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i700_2_lut (.I0(\Ki[14] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i506_2_lut (.I0(\Ki[10] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_5436));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i555_2_lut (.I0(\Ki[11] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_5435));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i749_2_lut (.I0(\Ki[15] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i604_2_lut (.I0(\Ki[12] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_5434));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i149_2_lut (.I0(\Kp[3] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_5376));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11882_bdd_4_lut_63571 (.I0(n11882), .I1(n75293), .I2(setpoint[21]), 
            .I3(n4736), .O(n79492));
    defparam n11882_bdd_4_lut_63571.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i653_2_lut (.I0(\Ki[13] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_5433));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n79492_bdd_4_lut (.I0(n79492), .I1(n535[21]), .I2(n455[21]), 
            .I3(n4736), .O(n79495));
    defparam n79492_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i702_2_lut (.I0(\Ki[14] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_5432));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i751_2_lut (.I0(\Ki[15] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11882_bdd_4_lut_63388 (.I0(n11882), .I1(n75257), .I2(setpoint[4]), 
            .I3(n4736), .O(n79270));
    defparam n11882_bdd_4_lut_63388.LUT_INIT = 16'he4aa;
    SB_LUT4 n11882_bdd_4_lut_63566 (.I0(n11882), .I1(n75292), .I2(setpoint[20]), 
            .I3(n4736), .O(n79486));
    defparam n11882_bdd_4_lut_63566.LUT_INIT = 16'he4aa;
    SB_LUT4 n79486_bdd_4_lut (.I0(n79486), .I1(n535[20]), .I2(n455[20]), 
            .I3(n4736), .O(n79489));
    defparam n79486_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n79270_bdd_4_lut (.I0(n79270), .I1(n535[4]), .I2(n475), .I3(n4736), 
            .O(n79273));
    defparam n79270_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11882_bdd_4_lut_63561 (.I0(n11882), .I1(n75291), .I2(setpoint[19]), 
            .I3(n4736), .O(n79480));
    defparam n11882_bdd_4_lut_63561.LUT_INIT = 16'he4aa;
    SB_LUT4 n79480_bdd_4_lut (.I0(n79480), .I1(n535[19]), .I2(n460), .I3(n4736), 
            .O(n79483));
    defparam n79480_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11882_bdd_4_lut_63383 (.I0(n11882), .I1(n75256), .I2(setpoint[3]), 
            .I3(n4736), .O(n79264));
    defparam n11882_bdd_4_lut_63383.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_21_i7_3_lut (.I0(n233[6]), .I1(n285[6]), .I2(n284), .I3(GND_net), 
            .O(n310[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n79264_bdd_4_lut (.I0(n79264), .I1(n535[3]), .I2(n455[3]), 
            .I3(n4736), .O(n79267));
    defparam n79264_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_22_i7_3_lut (.I0(n310[6]), .I1(IntegralLimit[6]), .I2(n258), 
            .I3(GND_net), .O(n353));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i61_2_lut (.I0(\Ki[1] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i14_2_lut (.I0(\Ki[0] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5373));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11882_bdd_4_lut_63556 (.I0(n11882), .I1(n75289), .I2(setpoint[18]), 
            .I3(n4736), .O(n79474));
    defparam n11882_bdd_4_lut_63556.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i110_2_lut (.I0(\Ki[2] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i159_2_lut (.I0(\Ki[3] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_5372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i208_2_lut (.I0(\Ki[4] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_5371));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i257_2_lut (.I0(\Ki[5] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i306_2_lut (.I0(\Ki[6] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i355_2_lut (.I0(\Ki[7] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n79474_bdd_4_lut (.I0(n79474), .I1(n535[18]), .I2(n461), .I3(n4736), 
            .O(n79477));
    defparam n79474_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i404_2_lut (.I0(\Ki[8] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i453_2_lut (.I0(\Ki[9] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i502_2_lut (.I0(\Ki[10] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i551_2_lut (.I0(\Ki[11] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i600_2_lut (.I0(\Ki[12] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i79_2_lut (.I0(\Kp[1] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11882_bdd_4_lut_63378 (.I0(n11882), .I1(n75255), .I2(setpoint[2]), 
            .I3(n4736), .O(n79258));
    defparam n11882_bdd_4_lut_63378.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i32_2_lut (.I0(\Kp[0] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_5420));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i649_2_lut (.I0(\Ki[13] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i198_2_lut (.I0(\Kp[4] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_5370));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i698_2_lut (.I0(\Ki[14] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n79258_bdd_4_lut (.I0(n79258), .I1(n535[2]), .I2(n455[2]), 
            .I3(n4736), .O(n79261));
    defparam n79258_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i747_2_lut (.I0(\Ki[15] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11882_bdd_4_lut_63551 (.I0(n11882), .I1(n75288), .I2(setpoint[17]), 
            .I3(n4736), .O(n79468));
    defparam n11882_bdd_4_lut_63551.LUT_INIT = 16'he4aa;
    SB_LUT4 n79468_bdd_4_lut (.I0(n79468), .I1(n535[17]), .I2(n462), .I3(n4736), 
            .O(n79471));
    defparam n79468_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11882_bdd_4_lut_63546 (.I0(n11882), .I1(n75287), .I2(setpoint[16]), 
            .I3(n4736), .O(n79462));
    defparam n11882_bdd_4_lut_63546.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i128_2_lut (.I0(\Kp[2] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i17_3_lut (.I0(n233[16]), .I1(n285[16]), .I2(n284), 
            .I3(GND_net), .O(n310[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i17_3_lut (.I0(n310[16]), .I1(IntegralLimit[16]), .I2(n258), 
            .I3(GND_net), .O(n343));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n79462_bdd_4_lut (.I0(n79462), .I1(n535[16]), .I2(n455[16]), 
            .I3(n4736), .O(n79465));
    defparam n79462_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i44527_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n340), .I2(\Ki[1] ), 
            .I3(n37307), .O(n20418[0]));   // verilog/motorControl.v(61[29:40])
    defparam i44527_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_21_i16_3_lut (.I0(n233[15]), .I1(n285[15]), .I2(n284), 
            .I3(GND_net), .O(n310[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44529_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n340), .I2(\Ki[1] ), 
            .I3(n37307), .O(n58586));   // verilog/motorControl.v(61[29:40])
    defparam i44529_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mux_22_i16_3_lut (.I0(n310[15]), .I1(IntegralLimit[15]), .I2(n258), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_21_i13_3_lut (.I0(n233[12]), .I1(n285[12]), .I2(n284), 
            .I3(GND_net), .O(n322));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i12_3_lut (.I0(n233[11]), .I1(n285[11]), .I2(n284), 
            .I3(GND_net), .O(n310[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i12_3_lut (.I0(n310[11]), .I1(IntegralLimit[11]), .I2(n258), 
            .I3(GND_net), .O(n348));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11882_bdd_4_lut_63373 (.I0(n11882), .I1(n75254), .I2(setpoint[1]), 
            .I3(n4736), .O(n79246));
    defparam n11882_bdd_4_lut_63373.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_21_i10_3_lut (.I0(n233[9]), .I1(n285[9]), .I2(n284), .I3(GND_net), 
            .O(n310[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i10_3_lut (.I0(n310[9]), .I1(IntegralLimit[9]), .I2(n258), 
            .I3(GND_net), .O(n350));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n79246_bdd_4_lut (.I0(n79246), .I1(n535[1]), .I2(n455[1]), 
            .I3(n4736), .O(n79249));
    defparam n79246_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1803 (.I0(\Ki[2] ), .I1(n340), .I2(n58814), 
            .I3(n20492[0]), .O(n20467));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_1803.LUT_INIT = 16'h8778;
    SB_LUT4 mult_23_i610_2_lut (.I0(\Kp[12] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i659_2_lut (.I0(\Kp[13] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i9_3_lut (.I0(n233[8]), .I1(n285[8]), .I2(n284), .I3(GND_net), 
            .O(n310[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i9_3_lut (.I0(n310[8]), .I1(IntegralLimit[8]), .I2(n258), 
            .I3(GND_net), .O(n351));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44747_3_lut_4_lut (.I0(\Ki[2] ), .I1(n340), .I2(n58814), 
            .I3(n20492[0]), .O(n4_adj_5288));   // verilog/motorControl.v(61[29:40])
    defparam i44747_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i44736_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n339), .I2(n340), 
            .I3(\Ki[1] ), .O(n58814));   // verilog/motorControl.v(61[29:40])
    defparam i44736_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i44734_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n339), .I2(n340), 
            .I3(\Ki[1] ), .O(n20468));   // verilog/motorControl.v(61[29:40])
    defparam i44734_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i247_2_lut (.I0(\Kp[5] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_5366));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i85_2_lut (.I0(\Ki[1] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1804 (.I0(counter[6]), .I1(counter[3]), .I2(counter[0]), 
            .I3(counter[4]), .O(n69713));   // verilog/motorControl.v(27[8:42])
    defparam i3_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n69713), .I1(counter[8]), .I2(counter[5]), .I3(counter[2]), 
            .O(n18_adj_5695));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(counter[7]), .I1(n18_adj_5695), .I2(counter[1]), 
            .I3(counter[10]), .O(n20_adj_5696));
    defparam i9_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut (.I0(n44726), .I1(n25921), .I2(n508), .I3(GND_net), 
            .O(n4_adj_5467));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_2_lut (.I0(counter[9]), .I1(counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5697));   // verilog/motorControl.v(27[8:42])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(n7_adj_5697), .I1(counter[12]), .I2(counter[13]), 
            .I3(n20_adj_5696), .O(counter_31__N_3714));   // verilog/motorControl.v(27[8:42])
    defparam i4_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i59720_2_lut_4_lut (.I0(n455[21]), .I1(n535[21]), .I2(n455[9]), 
            .I3(n535[9]), .O(n75576));
    defparam i59720_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_21_i15_3_lut (.I0(n233[14]), .I1(n285[14]), .I2(n284), 
            .I3(GND_net), .O(n310[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i15_3_lut (.I0(n310[14]), .I1(IntegralLimit[14]), .I2(n258), 
            .I3(GND_net), .O(n345));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i77_2_lut (.I0(\Ki[1] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_5417));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i134_2_lut (.I0(\Ki[2] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i30_2_lut (.I0(\Ki[0] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_5416));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_3_lut (.I0(\Kp[2] ), .I1(\Kp[1] ), .I2(\Kp[0] ), 
            .I3(GND_net), .O(n69342));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i44584_2_lut_3_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n58648));   // verilog/motorControl.v(61[20:26])
    defparam i44584_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i59753_2_lut_4_lut (.I0(n455[16]), .I1(n535[16]), .I2(n455[7]), 
            .I3(n535[7]), .O(n75609));
    defparam i59753_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n11882_bdd_4_lut_63363 (.I0(n11882), .I1(n75241), .I2(setpoint[0]), 
            .I3(n4736), .O(n79222));
    defparam n11882_bdd_4_lut_63363.LUT_INIT = 16'he4aa;
    SB_LUT4 n79222_bdd_4_lut (.I0(n79222), .I1(n535[0]), .I2(n455[0]), 
            .I3(n4736), .O(n79225));
    defparam n79222_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i59796_2_lut (.I0(PWMLimit[8]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75261));
    defparam i59796_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i177_2_lut (.I0(\Kp[3] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59904_2_lut_4_lut (.I0(n455[8]), .I1(n48[8]), .I2(n475), 
            .I3(n48[4]), .O(n75760));
    defparam i59904_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i77_2_lut (.I0(\Kp[1] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i183_2_lut (.I0(\Ki[3] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i30_2_lut (.I0(\Kp[0] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i126_2_lut (.I0(\Kp[2] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_5365));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i175_2_lut (.I0(\Kp[3] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_5364));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i224_2_lut (.I0(\Kp[4] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_5363));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i273_2_lut (.I0(\Kp[5] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_5361));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i322_2_lut (.I0(\Kp[6] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_5360));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59879_2_lut_4_lut (.I0(n455[16]), .I1(n48[16]), .I2(n455[7]), 
            .I3(n48[7]), .O(n75735));
    defparam i59879_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i60008_2_lut_4_lut (.I0(deadband[9]), .I1(n455[9]), .I2(deadband[8]), 
            .I3(n455[8]), .O(n75864));
    defparam i60008_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i60001_2_lut_4_lut (.I0(deadband[11]), .I1(n455[11]), .I2(deadband[7]), 
            .I3(n455[7]), .O(n75857));
    defparam i60001_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i371_2_lut (.I0(\Kp[7] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_5359));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i420_2_lut (.I0(\Kp[8] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i469_2_lut (.I0(\Kp[9] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i518_2_lut (.I0(\Kp[10] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i6_3_lut (.I0(n233[5]), .I1(n285[5]), .I2(n284), .I3(GND_net), 
            .O(n310[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i6_3_lut (.I0(n310[5]), .I1(IntegralLimit[5]), .I2(n258), 
            .I3(GND_net), .O(n354));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i59_2_lut (.I0(\Ki[1] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i12_2_lut (.I0(\Ki[0] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5357));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i108_2_lut (.I0(\Ki[2] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i296_2_lut (.I0(\Kp[6] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_5356));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i157_2_lut (.I0(\Ki[3] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i206_2_lut (.I0(\Ki[4] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_5354));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i255_2_lut (.I0(\Ki[5] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i304_2_lut (.I0(\Ki[6] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_5353));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i353_2_lut (.I0(\Ki[7] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i402_2_lut (.I0(\Ki[8] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i451_2_lut (.I0(\Ki[9] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i500_2_lut (.I0(\Ki[10] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i549_2_lut (.I0(\Ki[11] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i598_2_lut (.I0(\Ki[12] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i647_2_lut (.I0(\Ki[13] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60170_2_lut_4_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(setpoint[9]), 
            .I3(n535[9]), .O(n76026));
    defparam i60170_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i696_2_lut (.I0(\Ki[14] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i745_2_lut (.I0(\Ki[15] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i5_3_lut (.I0(n233[4]), .I1(n285[4]), .I2(n284), .I3(GND_net), 
            .O(n310[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60188_2_lut_4_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(setpoint[7]), 
            .I3(n535[7]), .O(n76044));
    defparam i60188_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_22_i5_3_lut (.I0(n310[4]), .I1(IntegralLimit[4]), .I2(n258), 
            .I3(GND_net), .O(n355));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i57_2_lut (.I0(\Ki[1] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i10_2_lut (.I0(\Ki[0] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_5348));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i106_2_lut (.I0(\Ki[2] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i155_2_lut (.I0(\Ki[3] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59646_2_lut (.I0(PWMLimit[9]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75262));
    defparam i59646_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59819_2_lut_4_lut (.I0(PWMLimit[19]), .I1(n460), .I2(PWMLimit[15]), 
            .I3(n455[15]), .O(n75675));
    defparam i59819_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i204_2_lut (.I0(\Ki[4] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_5344));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i253_2_lut (.I0(\Ki[5] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i302_2_lut (.I0(\Ki[6] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_5342));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i351_2_lut (.I0(\Ki[7] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i400_2_lut (.I0(\Ki[8] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59795_2_lut (.I0(PWMLimit[10]), .I1(n5076), .I2(GND_net), 
            .I3(GND_net), .O(n75263));
    defparam i59795_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i449_2_lut (.I0(\Ki[9] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i498_2_lut (.I0(\Ki[10] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59846_2_lut_4_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(PWMLimit[4]), 
            .I3(n475), .O(n75702));
    defparam i59846_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i24_3_lut_3_lut (.I0(setpoint[11]), .I1(setpoint[12]), 
            .I2(PWMLimit[12]), .I3(GND_net), .O(n24_adj_5248));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i547_2_lut (.I0(\Ki[11] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60298_2_lut_4_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), .I2(PWMLimit[13]), 
            .I3(setpoint[13]), .O(n76154));
    defparam i60298_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i596_2_lut (.I0(\Ki[12] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i645_2_lut (.I0(\Ki[13] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i26_3_lut_3_lut (.I0(setpoint[13]), .I1(setpoint[17]), 
            .I2(PWMLimit[17]), .I3(GND_net), .O(n26));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60306_2_lut_4_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), .I2(PWMLimit[14]), 
            .I3(setpoint[14]), .O(n76162));
    defparam i60306_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i694_2_lut (.I0(\Ki[14] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i743_2_lut (.I0(\Ki[15] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i28_3_lut_3_lut (.I0(setpoint[14]), .I1(setpoint[15]), 
            .I2(PWMLimit[15]), .I3(GND_net), .O(n28));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60038_2_lut_4_lut (.I0(n233[21]), .I1(n285[21]), .I2(n233[9]), 
            .I3(n285[9]), .O(n75894));
    defparam i60038_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i75_2_lut (.I0(\Kp[1] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i28_2_lut (.I0(\Kp[0] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5328));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i60104_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n233[21]), .I2(IntegralLimit[9]), 
            .I3(n233[9]), .O(n75960));
    defparam i60104_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i60063_2_lut_4_lut (.I0(n233[16]), .I1(n285[16]), .I2(n233[7]), 
            .I3(n285[7]), .O(n75919));
    defparam i60063_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i60120_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n233[16]), .I2(IntegralLimit[7]), 
            .I3(n233[7]), .O(n75976));
    defparam i60120_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i232_2_lut (.I0(\Ki[4] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n344_c));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_21_i23_3_lut (.I0(n233[22]), .I1(n285[22]), .I2(n284), 
            .I3(GND_net), .O(n310[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_3_lut (.I0(n310[22]), .I1(IntegralLimit[22]), .I2(n258), 
            .I3(GND_net), .O(n337));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i46_2_lut (.I0(\Ki[0] ), .I1(n337), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_5292));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i187_2_lut (.I0(\Ki[3] ), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n277));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i187_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i18_3_lut (.I0(n233[17]), .I1(n285[17]), .I2(n284), 
            .I3(GND_net), .O(n310[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i18_3_lut (.I0(n310[17]), .I1(IntegralLimit[17]), .I2(n258), 
            .I3(GND_net), .O(n342));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i22_3_lut (.I0(n233[21]), .I1(n285[21]), .I2(n284), 
            .I3(GND_net), .O(n313));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (\a_new[1] , \b_new[1] , debounce_cnt_N_3833, 
            ENCODER1_B_N_keep, n1779, ENCODER1_A_N_keep, b_prev, GND_net, 
            n1786, n1788, n1790, n1792, n1794, n1796, \encoder1_position[25] , 
            \encoder1_position[24] , \encoder1_position[23] , \encoder1_position[22] , 
            \encoder1_position[21] , \encoder1_position[20] , \encoder1_position[19] , 
            \encoder1_position[18] , \encoder1_position[17] , \encoder1_position[16] , 
            \encoder1_position[15] , \encoder1_position[14] , \encoder1_position[13] , 
            \encoder1_position[12] , \encoder1_position[11] , \encoder1_position[10] , 
            \encoder1_position[9] , \encoder1_position[8] , \encoder1_position[7] , 
            \encoder1_position[6] , \encoder1_position[5] , \encoder1_position[4] , 
            \encoder1_position[3] , \encoder1_position[2] , n1822, n1824, 
            VCC_net, n30013, a_prev, n29959, n29958, n1784, position_31__N_3836) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    output \b_new[1] ;
    output debounce_cnt_N_3833;
    input ENCODER1_B_N_keep;
    input n1779;
    input ENCODER1_A_N_keep;
    output b_prev;
    input GND_net;
    output n1786;
    output n1788;
    output n1790;
    output n1792;
    output n1794;
    output n1796;
    output \encoder1_position[25] ;
    output \encoder1_position[24] ;
    output \encoder1_position[23] ;
    output \encoder1_position[22] ;
    output \encoder1_position[21] ;
    output \encoder1_position[20] ;
    output \encoder1_position[19] ;
    output \encoder1_position[18] ;
    output \encoder1_position[17] ;
    output \encoder1_position[16] ;
    output \encoder1_position[15] ;
    output \encoder1_position[14] ;
    output \encoder1_position[13] ;
    output \encoder1_position[12] ;
    output \encoder1_position[11] ;
    output \encoder1_position[10] ;
    output \encoder1_position[9] ;
    output \encoder1_position[8] ;
    output \encoder1_position[7] ;
    output \encoder1_position[6] ;
    output \encoder1_position[5] ;
    output \encoder1_position[4] ;
    output \encoder1_position[3] ;
    output \encoder1_position[2] ;
    output n1822;
    output n1824;
    input VCC_net;
    input n30013;
    output a_prev;
    input n29959;
    input n29958;
    output n1784;
    output position_31__N_3836;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire direction_N_3840;
    wire [31:0]n133;
    
    wire n60218, n60217, n60216, n60215, n60214, n60213, n60212, 
        n60211, n60210, n60209, n60208, n60207, n60206, n60205, 
        n60204, n60203, n60202, n60201, n60200, n60199, n60198, 
        n60197, n60196, n60195, n60194, n60193, n60192, n60191, 
        n60190, n60189, n60188;
    
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 position_2041_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1786), .I3(n60218), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2041_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1788), .I3(n60217), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_32 (.CI(n60217), .I0(direction_N_3840), 
            .I1(n1788), .CO(n60218));
    SB_LUT4 position_2041_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1790), .I3(n60216), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_31 (.CI(n60216), .I0(direction_N_3840), 
            .I1(n1790), .CO(n60217));
    SB_LUT4 position_2041_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1792), .I3(n60215), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_30 (.CI(n60215), .I0(direction_N_3840), 
            .I1(n1792), .CO(n60216));
    SB_LUT4 position_2041_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1794), .I3(n60214), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_29 (.CI(n60214), .I0(direction_N_3840), 
            .I1(n1794), .CO(n60215));
    SB_LUT4 position_2041_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1796), .I3(n60213), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_28 (.CI(n60213), .I0(direction_N_3840), 
            .I1(n1796), .CO(n60214));
    SB_LUT4 position_2041_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[25] ), .I3(n60212), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_27 (.CI(n60212), .I0(direction_N_3840), 
            .I1(\encoder1_position[25] ), .CO(n60213));
    SB_LUT4 position_2041_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[24] ), .I3(n60211), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_26 (.CI(n60211), .I0(direction_N_3840), 
            .I1(\encoder1_position[24] ), .CO(n60212));
    SB_LUT4 position_2041_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[23] ), .I3(n60210), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_25 (.CI(n60210), .I0(direction_N_3840), 
            .I1(\encoder1_position[23] ), .CO(n60211));
    SB_LUT4 position_2041_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[22] ), .I3(n60209), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_24 (.CI(n60209), .I0(direction_N_3840), 
            .I1(\encoder1_position[22] ), .CO(n60210));
    SB_LUT4 position_2041_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[21] ), .I3(n60208), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_23 (.CI(n60208), .I0(direction_N_3840), 
            .I1(\encoder1_position[21] ), .CO(n60209));
    SB_LUT4 position_2041_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[20] ), .I3(n60207), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_22 (.CI(n60207), .I0(direction_N_3840), 
            .I1(\encoder1_position[20] ), .CO(n60208));
    SB_LUT4 position_2041_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[19] ), .I3(n60206), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_21 (.CI(n60206), .I0(direction_N_3840), 
            .I1(\encoder1_position[19] ), .CO(n60207));
    SB_LUT4 position_2041_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[18] ), .I3(n60205), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_20 (.CI(n60205), .I0(direction_N_3840), 
            .I1(\encoder1_position[18] ), .CO(n60206));
    SB_LUT4 position_2041_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[17] ), .I3(n60204), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_19 (.CI(n60204), .I0(direction_N_3840), 
            .I1(\encoder1_position[17] ), .CO(n60205));
    SB_LUT4 position_2041_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[16] ), .I3(n60203), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_18 (.CI(n60203), .I0(direction_N_3840), 
            .I1(\encoder1_position[16] ), .CO(n60204));
    SB_LUT4 position_2041_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[15] ), .I3(n60202), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_17 (.CI(n60202), .I0(direction_N_3840), 
            .I1(\encoder1_position[15] ), .CO(n60203));
    SB_LUT4 position_2041_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[14] ), .I3(n60201), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_16 (.CI(n60201), .I0(direction_N_3840), 
            .I1(\encoder1_position[14] ), .CO(n60202));
    SB_LUT4 position_2041_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[13] ), .I3(n60200), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_15 (.CI(n60200), .I0(direction_N_3840), 
            .I1(\encoder1_position[13] ), .CO(n60201));
    SB_LUT4 position_2041_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[12] ), .I3(n60199), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_14 (.CI(n60199), .I0(direction_N_3840), 
            .I1(\encoder1_position[12] ), .CO(n60200));
    SB_LUT4 position_2041_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[11] ), .I3(n60198), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_13 (.CI(n60198), .I0(direction_N_3840), 
            .I1(\encoder1_position[11] ), .CO(n60199));
    SB_LUT4 position_2041_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[10] ), .I3(n60197), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_12 (.CI(n60197), .I0(direction_N_3840), 
            .I1(\encoder1_position[10] ), .CO(n60198));
    SB_LUT4 position_2041_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[9] ), .I3(n60196), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_11 (.CI(n60196), .I0(direction_N_3840), 
            .I1(\encoder1_position[9] ), .CO(n60197));
    SB_LUT4 position_2041_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[8] ), .I3(n60195), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_10 (.CI(n60195), .I0(direction_N_3840), 
            .I1(\encoder1_position[8] ), .CO(n60196));
    SB_LUT4 position_2041_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[7] ), .I3(n60194), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_9 (.CI(n60194), .I0(direction_N_3840), 
            .I1(\encoder1_position[7] ), .CO(n60195));
    SB_LUT4 position_2041_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[6] ), .I3(n60193), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_8 (.CI(n60193), .I0(direction_N_3840), 
            .I1(\encoder1_position[6] ), .CO(n60194));
    SB_LUT4 position_2041_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[5] ), .I3(n60192), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_7 (.CI(n60192), .I0(direction_N_3840), 
            .I1(\encoder1_position[5] ), .CO(n60193));
    SB_LUT4 position_2041_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[4] ), .I3(n60191), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_6 (.CI(n60191), .I0(direction_N_3840), 
            .I1(\encoder1_position[4] ), .CO(n60192));
    SB_LUT4 position_2041_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[3] ), .I3(n60190), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_5 (.CI(n60190), .I0(direction_N_3840), 
            .I1(\encoder1_position[3] ), .CO(n60191));
    SB_LUT4 position_2041_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[2] ), .I3(n60189), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_4 (.CI(n60189), .I0(direction_N_3840), 
            .I1(\encoder1_position[2] ), .CO(n60190));
    SB_LUT4 position_2041_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1822), .I3(n60188), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_3 (.CI(n60188), .I0(direction_N_3840), 
            .I1(n1822), .CO(n60189));
    SB_LUT4 position_2041_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1824), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n1824), 
            .CO(n60188));
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n30013));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29959));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1784), .C(n1779), .D(n29958));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i0 (.Q(n1824), .C(n1779), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i31 (.Q(n1786), .C(n1779), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i30 (.Q(n1788), .C(n1779), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i29 (.Q(n1790), .C(n1779), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i28 (.Q(n1792), .C(n1779), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i27 (.Q(n1794), .C(n1779), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i26 (.Q(n1796), .C(n1779), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i25 (.Q(\encoder1_position[25] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i24 (.Q(\encoder1_position[24] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i23 (.Q(\encoder1_position[23] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i22 (.Q(\encoder1_position[22] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i21 (.Q(\encoder1_position[21] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i20 (.Q(\encoder1_position[20] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i19 (.Q(\encoder1_position[19] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i18 (.Q(\encoder1_position[18] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i17 (.Q(\encoder1_position[17] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i16 (.Q(\encoder1_position[16] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i15 (.Q(\encoder1_position[15] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i14 (.Q(\encoder1_position[14] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i13 (.Q(\encoder1_position[13] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i12 (.Q(\encoder1_position[12] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i11 (.Q(\encoder1_position[11] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i10 (.Q(\encoder1_position[10] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i9 (.Q(\encoder1_position[9] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i8 (.Q(\encoder1_position[8] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i7 (.Q(\encoder1_position[7] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i6 (.Q(\encoder1_position[6] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i5 (.Q(\encoder1_position[5] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i4 (.Q(\encoder1_position[4] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i3 (.Q(\encoder1_position[3] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i2 (.Q(\encoder1_position[2] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i1 (.Q(n1822), .C(n1779), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module coms
//

module coms (VCC_net, clk16MHz, \Kp[6] , \data_out_frame[7] , \FRAME_MATCHER.i_31__N_2509 , 
            encoder0_position_scaled, byte_transmit_counter, \data_out_frame[25] , 
            \data_out_frame[24] , n2874, \data_out_frame[8] , n66744, 
            n66703, \FRAME_MATCHER.state[3] , reset, rx_data, \data_in_frame[11] , 
            \Kp[5] , GND_net, \Kp[4] , \data_out_frame[1][6] , \data_out_frame[3][6] , 
            \data_out_frame[6] , \data_out_frame[23] , \data_out_frame[18] , 
            \data_out_frame[22] , n67085, n79, \data_out_frame[4] , 
            \data_out_frame[5] , \Kp[3] , \data_out_frame[21] , n25419, 
            \data_out_frame[20] , n67203, n26999, \Kp[2] , displacement, 
            DE_c, \Kp[1] , \data_out_frame[17] , pwm_setpoint, IntegralLimit, 
            n24045, LED_c, \data_out_frame[1][5] , n30193, \data_in_frame[6] , 
            n30190, n30187, n30184, n30181, \data_out_frame[16] , 
            n30178, n26619, \data_out_frame[1][3] , n69502, \data_out_frame[15] , 
            \data_out_frame[19] , \data_out_frame[14] , setpoint, n62277, 
            n62302, n30175, n29359, \data_in_frame[12][6] , \data_in_frame[19] , 
            \data_in_frame[16] , deadband, \data_out_frame[13] , n66700, 
            n30172, n8, n67425, \data_in_frame[16][7] , \data_out_frame[1][7] , 
            \data_out_frame[3][7] , n28392, n30169, \data_in_frame[5] , 
            n66699, n72460, n72458, n66577, n66698, \data_out_frame[9] , 
            n66697, n66696, n66695, n66694, n27, n66693, n66692, 
            n66691, \data_out_frame[10] , n66690, n66689, n66688, 
            n66687, n66686, n66685, \data_out_frame[1][0] , n66684, 
            n66683, \data_out_frame[11] , n66682, n66681, n66680, 
            n66679, n66678, n66677, n66676, n66675, \data_out_frame[12] , 
            n66674, n66673, n66672, n66671, n66670, n66669, \data_in_frame[15][5] , 
            n66668, n30166, n66667, \FRAME_MATCHER.i[1] , \data_in_frame[14] , 
            \FRAME_MATCHER.i[2] , n66666, n25421, n30163, n30160, 
            n30157, n30154, \data_in_frame[14][2] , n30151, n66665, 
            n67274, n30148, \FRAME_MATCHER.i[0] , n62281, \data_in_frame[14][4] , 
            n69075, \data_in_frame[14][5] , \data_in_frame[14][6] , \data_in_frame[14][7] , 
            \data_in_frame[13][2] , n66664, \data_in_frame[13][4] , n30145, 
            \data_in_frame[4] , \data_in_frame[13][5] , \data_in_frame[13][6] , 
            n30141, n30138, n8_adj_5, n30135, \data_in_frame[13][7] , 
            n30132, n23094, n30129, n67599, n30126, n30123, n67361, 
            \data_in_frame[12][2] , \data_in_frame[12][3] , PWMLimit, 
            n35, \data_in_frame[12][5] , n462, n36361, \data_in_frame[12][4] , 
            n105, control_mode, control_update, n24, n30, n27184, 
            \data_out_frame[0][4] , \data_out_frame[3][4] , \data_out_frame[0][2] , 
            n66663, \data_out_frame[0][3] , \data_out_frame[3][3] , n66662, 
            n66661, n66660, n66659, n66658, n66657, n66656, n66655, 
            n66654, n66653, n66652, \data_out_frame[1][1] , \data_out_frame[3][1] , 
            n66651, \Kp[7] , \Kp[8] , \Kp[9] , n66650, n66649, \Kp[10] , 
            \Kp[11] , \Kp[12] , n66648, n66647, n66646, \Kp[13] , 
            \Kp[14] , \Kp[15] , \Ki[1] , \Ki[2] , \Ki[3] , n66645, 
            n66644, n66643, n66642, \Ki[4] , \Ki[5] , n66641, \Ki[6] , 
            \Ki[7] , n66580, n66581, n66582, \Ki[8] , \Ki[9] , \Ki[10] , 
            n66583, \Ki[11] , n66584, n66585, n66586, \Ki[12] , 
            n66588, n30873, n29288, n66589, n66590, \Ki[13] , \Ki[14] , 
            \Ki[15] , n66591, n66592, n66593, n66594, n66595, n66596, 
            n66578, n30883, n29278, n30007, \FRAME_MATCHER.rx_data_ready_prev , 
            n30003, neopxl_color, n30002, n30001, n30000, n29999, 
            n29998, n29997, n29996, n29995, n29994, n29993, n75275, 
            n29991, n29990, n29989, n29988, n29987, n29984, \control_mode[5] , 
            n29983, \control_mode[6] , n29979, \control_mode[7] , n29976, 
            \current_limit[1] , n29975, \current_limit[2] , n29974, 
            \current_limit[3] , n29973, \current_limit[4] , n29972, 
            \current_limit[5] , n29943, \current_limit[0] , n29941, 
            \Ki[0] , \Kp[0] , n66597, n66598, n66599, n66600, n66601, 
            n66602, n29271, n66603, n66604, n66605, n66606, n66607, 
            n66576, n66608, n29263, n66609, n29261, n66610, n66611, 
            n66612, n66613, n66614, n66615, n66616, n29253, n66617, 
            n29251, n66618, n66619, n66620, n66621, n66743, n66742, 
            n66741, n38, n460, n486, n40, n41637, n66852, n34, 
            n36, n66740, n66739, n30786, \current_limit[8] , n45283, 
            encoder1_position_scaled, n53108, n42994, n30785, \current_limit[9] , 
            n30781, \current_limit[10] , n30779, \current_limit[12] , 
            n65900, \data_in_frame[18] , n65896, n65892, n65888, \motor_state_23__N_91[12] , 
            n15, n10, n29731, n29734, n30740, n65884, n29740, 
            n30734, n29746, \data_in_frame[19][2] , n30727, \data_in_frame[17] , 
            n29749, \data_in_frame[19][3] , n29752, \data_in_frame[19][4] , 
            n29756, \data_in_frame[19][5] , n30678, n30666, \data_in_frame[9] , 
            n66738, n30632, n30249, n29759, \data_in_frame[19][6] , 
            n30252, n30255, n29763, \data_in_frame[19][7] , n30258, 
            n30261, n30264, n30619, n30616, n66737, \data_in_frame[20][0] , 
            \data_in_frame[20][1] , \data_in_frame[20][2] , \data_in_frame[20][4] , 
            n29794, \data_in_frame[21] , n29797, n30267, n30603, n29800, 
            n29803, n30593, n29806, n30589, n30588, n29809, n30585, 
            n29812, n29815, n29818, \data_in_frame[22] , n66142, n30349, 
            \data_in_frame[13][0] , n30355, n30362, n30365, n30368, 
            n30372, n30375, n66736, n66735, n30382, n30388, n30392, 
            n30395, n30398, n65878, \data_in_frame[16][0] , n30432, 
            n65874, n65870, n65842, n65866, n65960, n30458, n65998, 
            n65994, n65990, n30517, n66734, n29821, n29824, n29827, 
            n29830, n29833, n29836, n29839, n29842, \data_in_frame[23] , 
            n29845, n65966, n30469, n29863, n65964, n65962, n29872, 
            n26875, \data_in_frame[1][1] , \data_in_frame[1][2] , \data_in_frame[1][3] , 
            \data_in_frame[1][5] , \data_in_frame[1][6] , \data_in_frame[1][7] , 
            n66733, n66732, n66731, n66730, n66729, n66728, n66727, 
            n66726, n26311, n66725, n66724, n66723, n26475, n29387, 
            n66722, n66721, n66720, n66719, n66718, n66717, n66716, 
            n66715, n66714, n66713, n66712, n66711, n29374, n66710, 
            n66622, n66623, n29755, \current_limit[6] , n31022, n29244, 
            n31023, n29243, n66624, n66625, n66626, n66627, n66628, 
            n66629, n29236, n31031, n29235, n66587, n66630, n31034, 
            n29232, n66709, n82, n28703, n28672, n66708, n66707, 
            n31038, n29369, n31039, n29231, n66631, n66632, n66633, 
            n66634, n66635, n66636, n31046, n29224, n66579, n66637, 
            n66638, n66639, n66640, n61795, n66706, n31088, n29367, 
            n29727, \current_limit[7] , n31093, n29366, n66705, n66704, 
            n66702, n66701, n15_adj_6, rx_data_ready, n15_adj_7, \motor_state_23__N_91[8] , 
            n25590, n66867, n66869, n66862, \current[7] , \current[6] , 
            \current[5] , n67584, \current[4] , n461, n38_adj_8, n75815, 
            n6, n3476, n66945, ID, n79417, n79243, n1, n5, n67259, 
            n27089, n69485, n67194, n6_adj_9, n69065, n16, n67500, 
            n67135, n69463, n27243, n26760, n61396, n67238, n67596, 
            n67235, n89, n4, Kp_23__N_1389, n25921, \current[3] , 
            \current[2] , \current[1] , \current[0] , \current[15] , 
            n8_adj_10, n67578, n8_adj_11, n67243, n61406, n67213, 
            n28715, n75246, n27203, n66853, \current[11] , \current[10] , 
            \current[9] , \current[8] , n28730, n75250, n28717, n10_adj_12, 
            n66872, n66866, n79237, tx_active, n23025, n79447, n51, 
            n22, n260, tx_o, r_SM_Main, n29956, r_Clock_Count, n5220, 
            n27_adj_13, n67730, n6_adj_14, tx_enable, r_Clock_Count_adj_26, 
            baudrate, n28240, n67800, \r_SM_Main[2]_adj_23 , r_Rx_Data, 
            RX_N_2, \o_Rx_DV_N_3488[8] , n5217, n66790, \r_SM_Main[1]_adj_24 , 
            n28117, n70292, n29937, n29936, n29934, n29915, n29914, 
            n29910, n29906, n30762, n62510, n30758, \r_Bit_Index[0] , 
            n70662, n34_adj_25, \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , 
            n70340, n70356, n70276, n70324, n70308, n70388, n70372) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    input clk16MHz;
    output \Kp[6] ;
    output [7:0]\data_out_frame[7] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input [23:0]encoder0_position_scaled;
    output [7:0]byte_transmit_counter;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[24] ;
    input n2874;
    output [7:0]\data_out_frame[8] ;
    input n66744;
    input n66703;
    output \FRAME_MATCHER.state[3] ;
    input reset;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[11] ;
    output \Kp[5] ;
    input GND_net;
    output \Kp[4] ;
    output \data_out_frame[1][6] ;
    output \data_out_frame[3][6] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[22] ;
    input n67085;
    output n79;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output \Kp[3] ;
    output [7:0]\data_out_frame[21] ;
    input n25419;
    output [7:0]\data_out_frame[20] ;
    input n67203;
    input n26999;
    output \Kp[2] ;
    input [23:0]displacement;
    output DE_c;
    output \Kp[1] ;
    output [7:0]\data_out_frame[17] ;
    input [23:0]pwm_setpoint;
    output [23:0]IntegralLimit;
    input n24045;
    output LED_c;
    output \data_out_frame[1][5] ;
    input n30193;
    output [7:0]\data_in_frame[6] ;
    input n30190;
    input n30187;
    input n30184;
    input n30181;
    output [7:0]\data_out_frame[16] ;
    input n30178;
    output n26619;
    output \data_out_frame[1][3] ;
    output n69502;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[14] ;
    output [23:0]setpoint;
    output n62277;
    input n62302;
    input n30175;
    input n29359;
    output \data_in_frame[12][6] ;
    output [7:0]\data_in_frame[19] ;
    output [7:0]\data_in_frame[16] ;
    output [23:0]deadband;
    output [7:0]\data_out_frame[13] ;
    input n66700;
    input n30172;
    input n8;
    input n67425;
    output \data_in_frame[16][7] ;
    output \data_out_frame[1][7] ;
    output \data_out_frame[3][7] ;
    output n28392;
    input n30169;
    output [7:0]\data_in_frame[5] ;
    input n66699;
    input n72460;
    input n72458;
    input n66577;
    input n66698;
    output [7:0]\data_out_frame[9] ;
    input n66697;
    input n66696;
    input n66695;
    input n66694;
    input n27;
    input n66693;
    input n66692;
    input n66691;
    output [7:0]\data_out_frame[10] ;
    input n66690;
    input n66689;
    input n66688;
    input n66687;
    input n66686;
    input n66685;
    output \data_out_frame[1][0] ;
    input n66684;
    input n66683;
    output [7:0]\data_out_frame[11] ;
    input n66682;
    input n66681;
    input n66680;
    input n66679;
    input n66678;
    input n66677;
    input n66676;
    input n66675;
    output [7:0]\data_out_frame[12] ;
    input n66674;
    input n66673;
    input n66672;
    input n66671;
    input n66670;
    input n66669;
    output \data_in_frame[15][5] ;
    input n66668;
    input n30166;
    input n66667;
    output \FRAME_MATCHER.i[1] ;
    output [7:0]\data_in_frame[14] ;
    output \FRAME_MATCHER.i[2] ;
    input n66666;
    input n25421;
    input n30163;
    input n30160;
    input n30157;
    input n30154;
    output \data_in_frame[14][2] ;
    input n30151;
    input n66665;
    output n67274;
    input n30148;
    output \FRAME_MATCHER.i[0] ;
    output n62281;
    output \data_in_frame[14][4] ;
    output n69075;
    output \data_in_frame[14][5] ;
    output \data_in_frame[14][6] ;
    output \data_in_frame[14][7] ;
    output \data_in_frame[13][2] ;
    input n66664;
    output \data_in_frame[13][4] ;
    input n30145;
    output [7:0]\data_in_frame[4] ;
    output \data_in_frame[13][5] ;
    output \data_in_frame[13][6] ;
    input n30141;
    input n30138;
    output n8_adj_5;
    input n30135;
    output \data_in_frame[13][7] ;
    input n30132;
    output n23094;
    input n30129;
    input n67599;
    input n30126;
    input n30123;
    output n67361;
    output \data_in_frame[12][2] ;
    output \data_in_frame[12][3] ;
    output [23:0]PWMLimit;
    output n35;
    output \data_in_frame[12][5] ;
    input n462;
    output n36361;
    output \data_in_frame[12][4] ;
    input n105;
    output [7:0]control_mode;
    input control_update;
    output n24;
    output n30;
    output n27184;
    output \data_out_frame[0][4] ;
    output \data_out_frame[3][4] ;
    output \data_out_frame[0][2] ;
    input n66663;
    output \data_out_frame[0][3] ;
    output \data_out_frame[3][3] ;
    input n66662;
    input n66661;
    input n66660;
    input n66659;
    input n66658;
    input n66657;
    input n66656;
    input n66655;
    input n66654;
    input n66653;
    input n66652;
    output \data_out_frame[1][1] ;
    output \data_out_frame[3][1] ;
    input n66651;
    output \Kp[7] ;
    output \Kp[8] ;
    output \Kp[9] ;
    input n66650;
    input n66649;
    output \Kp[10] ;
    output \Kp[11] ;
    output \Kp[12] ;
    input n66648;
    input n66647;
    input n66646;
    output \Kp[13] ;
    output \Kp[14] ;
    output \Kp[15] ;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    input n66645;
    input n66644;
    input n66643;
    input n66642;
    output \Ki[4] ;
    output \Ki[5] ;
    input n66641;
    output \Ki[6] ;
    output \Ki[7] ;
    input n66580;
    input n66581;
    input n66582;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    input n66583;
    output \Ki[11] ;
    input n66584;
    input n66585;
    input n66586;
    output \Ki[12] ;
    input n66588;
    input n30873;
    input n29288;
    input n66589;
    input n66590;
    output \Ki[13] ;
    output \Ki[14] ;
    output \Ki[15] ;
    input n66591;
    input n66592;
    input n66593;
    input n66594;
    input n66595;
    input n66596;
    input n66578;
    input n30883;
    input n29278;
    input n30007;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    input n30003;
    output [23:0]neopxl_color;
    input n30002;
    input n30001;
    input n30000;
    input n29999;
    input n29998;
    input n29997;
    input n29996;
    input n29995;
    input n29994;
    input n29993;
    input n75275;
    input n29991;
    input n29990;
    input n29989;
    input n29988;
    input n29987;
    input n29984;
    output \control_mode[5] ;
    input n29983;
    output \control_mode[6] ;
    input n29979;
    output \control_mode[7] ;
    input n29976;
    output \current_limit[1] ;
    input n29975;
    output \current_limit[2] ;
    input n29974;
    output \current_limit[3] ;
    input n29973;
    output \current_limit[4] ;
    input n29972;
    output \current_limit[5] ;
    input n29943;
    output \current_limit[0] ;
    input n29941;
    output \Ki[0] ;
    output \Kp[0] ;
    input n66597;
    input n66598;
    input n66599;
    input n66600;
    input n66601;
    input n66602;
    input n29271;
    input n66603;
    input n66604;
    input n66605;
    input n66606;
    input n66607;
    input n66576;
    input n66608;
    input n29263;
    input n66609;
    input n29261;
    input n66610;
    input n66611;
    input n66612;
    input n66613;
    input n66614;
    input n66615;
    input n66616;
    input n29253;
    input n66617;
    input n29251;
    input n66618;
    input n66619;
    input n66620;
    input n66621;
    input n66743;
    input n66742;
    input n66741;
    input n38;
    input n460;
    input n486;
    output n40;
    output n41637;
    output n66852;
    input n34;
    output n36;
    input n66740;
    input n66739;
    input n30786;
    output \current_limit[8] ;
    output n45283;
    input [23:0]encoder1_position_scaled;
    output n53108;
    output n42994;
    input n30785;
    output \current_limit[9] ;
    input n30781;
    output \current_limit[10] ;
    input n30779;
    output \current_limit[12] ;
    input n65900;
    output [7:0]\data_in_frame[18] ;
    input n65896;
    input n65892;
    input n65888;
    input \motor_state_23__N_91[12] ;
    output n15;
    output n10;
    input n29731;
    input n29734;
    input n30740;
    input n65884;
    input n29740;
    input n30734;
    input n29746;
    output \data_in_frame[19][2] ;
    input n30727;
    output [7:0]\data_in_frame[17] ;
    input n29749;
    output \data_in_frame[19][3] ;
    input n29752;
    output \data_in_frame[19][4] ;
    input n29756;
    output \data_in_frame[19][5] ;
    input n30678;
    input n30666;
    output [7:0]\data_in_frame[9] ;
    input n66738;
    input n30632;
    input n30249;
    input n29759;
    output \data_in_frame[19][6] ;
    input n30252;
    input n30255;
    input n29763;
    output \data_in_frame[19][7] ;
    input n30258;
    input n30261;
    input n30264;
    input n30619;
    input n30616;
    input n66737;
    output \data_in_frame[20][0] ;
    output \data_in_frame[20][1] ;
    output \data_in_frame[20][2] ;
    output \data_in_frame[20][4] ;
    input n29794;
    output [7:0]\data_in_frame[21] ;
    input n29797;
    input n30267;
    input n30603;
    input n29800;
    input n29803;
    input n30593;
    input n29806;
    input n30589;
    input n30588;
    input n29809;
    input n30585;
    input n29812;
    input n29815;
    input n29818;
    output [7:0]\data_in_frame[22] ;
    input n66142;
    input n30349;
    output \data_in_frame[13][0] ;
    input n30355;
    input n30362;
    input n30365;
    input n30368;
    input n30372;
    input n30375;
    input n66736;
    input n66735;
    input n30382;
    input n30388;
    input n30392;
    input n30395;
    input n30398;
    input n65878;
    output \data_in_frame[16][0] ;
    input n30432;
    input n65874;
    input n65870;
    input n65842;
    input n65866;
    input n65960;
    input n30458;
    input n65998;
    input n65994;
    input n65990;
    input n30517;
    input n66734;
    input n29821;
    input n29824;
    input n29827;
    input n29830;
    input n29833;
    input n29836;
    input n29839;
    input n29842;
    output [7:0]\data_in_frame[23] ;
    input n29845;
    input n65966;
    input n30469;
    input n29863;
    input n65964;
    input n65962;
    input n29872;
    output n26875;
    output \data_in_frame[1][1] ;
    output \data_in_frame[1][2] ;
    output \data_in_frame[1][3] ;
    output \data_in_frame[1][5] ;
    output \data_in_frame[1][6] ;
    output \data_in_frame[1][7] ;
    input n66733;
    input n66732;
    input n66731;
    input n66730;
    input n66729;
    input n66728;
    input n66727;
    input n66726;
    input n26311;
    input n66725;
    input n66724;
    input n66723;
    output n26475;
    input n29387;
    input n66722;
    input n66721;
    input n66720;
    input n66719;
    input n66718;
    input n66717;
    input n66716;
    input n66715;
    input n66714;
    input n66713;
    input n66712;
    input n66711;
    input n29374;
    input n66710;
    input n66622;
    input n66623;
    input n29755;
    output \current_limit[6] ;
    input n31022;
    input n29244;
    input n31023;
    input n29243;
    input n66624;
    input n66625;
    input n66626;
    input n66627;
    input n66628;
    input n66629;
    input n29236;
    input n31031;
    input n29235;
    input n66587;
    input n66630;
    input n31034;
    input n29232;
    input n66709;
    input n82;
    output n28703;
    output n28672;
    input n66708;
    input n66707;
    input n31038;
    input n29369;
    input n31039;
    input n29231;
    input n66631;
    input n66632;
    input n66633;
    input n66634;
    input n66635;
    input n66636;
    input n31046;
    input n29224;
    input n66579;
    input n66637;
    input n66638;
    input n66639;
    input n66640;
    output n61795;
    input n66706;
    input n31088;
    input n29367;
    input n29727;
    output \current_limit[7] ;
    input n31093;
    input n29366;
    input n66705;
    input n66704;
    input n66702;
    input n66701;
    output n15_adj_6;
    output rx_data_ready;
    output n15_adj_7;
    output \motor_state_23__N_91[8] ;
    output n25590;
    output n66867;
    output n66869;
    output n66862;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    output n67584;
    input \current[4] ;
    input n461;
    output n38_adj_8;
    output n75815;
    output n6;
    output n3476;
    output n66945;
    input [7:0]ID;
    input n79417;
    input n79243;
    input n1;
    input n5;
    output n67259;
    input n27089;
    input n69485;
    output n67194;
    input n6_adj_9;
    output n69065;
    output n16;
    input n67500;
    output n67135;
    output n69463;
    output n27243;
    input n26760;
    input n61396;
    output n67238;
    output n67596;
    output n67235;
    output n89;
    output n4;
    output Kp_23__N_1389;
    output n25921;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    input \current[15] ;
    output n8_adj_10;
    input n67578;
    output n8_adj_11;
    output n67243;
    output n61406;
    output n67213;
    output n28715;
    output n75246;
    output n27203;
    output n66853;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    output n28730;
    output n75250;
    input n28717;
    input n10_adj_12;
    output n66872;
    output n66866;
    input n79237;
    output tx_active;
    output n23025;
    output n79447;
    output n51;
    input n22;
    output n260;
    output tx_o;
    output [2:0]r_SM_Main;
    input n29956;
    output [8:0]r_Clock_Count;
    input n5220;
    output n27_adj_13;
    input n67730;
    output n6_adj_14;
    output tx_enable;
    output [7:0]r_Clock_Count_adj_26;
    input [31:0]baudrate;
    output n28240;
    output n67800;
    output \r_SM_Main[2]_adj_23 ;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[8] ;
    input n5217;
    input n66790;
    output \r_SM_Main[1]_adj_24 ;
    output n28117;
    output n70292;
    input n29937;
    input n29936;
    input n29934;
    input n29915;
    input n29914;
    input n29910;
    input n29906;
    input n30762;
    input n62510;
    input n30758;
    output \r_Bit_Index[0] ;
    output n70662;
    output n34_adj_25;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n70340;
    output n70356;
    output n70276;
    output n70324;
    output n70308;
    output n70388;
    output n70372;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n30243;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    
    wire n30240, Kp_23__N_612, Kp_23__N_1748;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    
    wire n30044, n30237;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n79426, n79429, n2_adj_4734, n2_adj_4735, n30234, n67126, 
        n3, n6_c, n62464, n3_adj_4736, n79420, n67451, n62476, 
        n3_adj_4737, n28674, n30320, n30045, n61789, n67055, n3_adj_4738, 
        n30046, n28394, n72477, n6_adj_4739, n67052, n3_adj_4740, 
        n61954, n62261, n67210, n67480, n27298, n67139, n14, n61312, 
        n10_c, n72478;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n67716, n72476, n30047, n67075, n79453, n75296, n61422, 
        n66953, n18, n27096, n20, n79363, n79135, n77507, n61681, 
        n16_c, n62428, n67485, n10_adj_4741;
    wire [7:0]\data_in_frame[11]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30316, n67512, n67572, n67453, n20_adj_4742, n67277, n26203, 
        n19, n26661, n61445, n21, n62290, n61412, n8_c, n62368, 
        n3_adj_4743, n30048, n67061, n67432, n3_adj_4744, n2_adj_4745, 
        tx_transmit_N_3416, \FRAME_MATCHER.i_31__N_2511 , n1_c, n6_adj_4746, 
        n66848, n27318, n2_adj_4747, n2_adj_4748, n30049, n2_adj_4749, 
        n2_adj_4750, n2_adj_4751, n67435, n26232, n12, n67557, n2_adj_4752, 
        n2_adj_4753, n2_adj_4754, n30050, n2_adj_4755, n30231, n6_adj_4756, 
        n3_adj_4757, n30228, n30225, n30222, n30219;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n29953;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_4758, n30215, n30212, n30209, n30206, n30203, n30200, 
        n30197, n2_adj_4759, n30051, LED_N_3408, LED_N_3407, n2_adj_4760, 
        n27770, \FRAME_MATCHER.i_31__N_2513 , n29211, n30052, n3_adj_4761, 
        n5_c, n2_adj_4762, n29962, n30053, n30054, n2_adj_4763, 
        n79423, n5_adj_4764, n25458, n69352, n3_adj_4765, n2_adj_4766, 
        n2_adj_4767, n62332, n3_adj_4768, n24041, n67132, n69736, 
        n3_adj_4769, n67503, n67509, n10_adj_4770, n2_adj_4771, n61447, 
        n3_adj_4772, n61324, n2_adj_4773, n2_adj_4774, n2_adj_4775, 
        n69543, n62253, n26829, n26517, n67176, n67158, n62013, 
        n61333, n12_adj_4776, n2_adj_4777, n67477, n2_adj_4778, n2_adj_4779, 
        n2_adj_4780, n30055, n61386, n61472, n2_adj_4781, n2_adj_4782, 
        n30056, n62285, n67252, n61824, n6_adj_4783, n61503, n2_adj_4784, 
        n2_adj_4785, n67010, n26089, n2_adj_4786, n26607, n2_adj_4787, 
        n7, n67058, n67326, n26060, n67388, n10_adj_4788, n66929, 
        n26645, n6_adj_4789, n67046, n61362, n30057, n61517, n67049, 
        n40_c, n67207, n38_c, n2_adj_4790, n30_c, n66967, n44, 
        n2_adj_4791, n69868, n42, n26, n67506, n43, n27258, n41, 
        n2_adj_4792, n67280, n44_adj_4793, n61320, n14_adj_4794, n9, 
        n67216;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    
    wire n30058, n60995, n26943, n67222, n6_adj_4795, n2_adj_4796, 
        n2_adj_4797, n2_adj_4798, n30059;
    wire [23:0]n4932;
    
    wire n61434, n30095, n79408, n79411, n67491, n2068, n30094, 
        n66886, n30093, n28131, n1720, n2_adj_4799, n30092, n2_adj_4800, 
        n7_adj_4802, n62080, n8_adj_4803, n67271, n2_adj_4804, n79402, 
        n2_adj_4805, n79435, n75277;
    wire [7:0]\data_in_frame[16]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30091, n79375, n79201, n77345, n30090, n2_adj_4806, n30089, 
        n2_adj_4807, n79405;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n30088, n79396, n2_adj_4808, n67332, n10_adj_4809, n68641, 
        n24023, n8_adj_4810, n7_adj_4811, n28327, n28651, n60249, 
        n75190, n28329, n60248, n75189, n79399, n28331, n60247, 
        n75181, n2_adj_4812, n6_adj_4813, n28333, n60246, n75171, 
        n28337, n60245, n75168, n2_adj_4814, n7_adj_4815, n30087, 
        n61577, n67291, n79459, n75267, n2_adj_4816, n2_adj_4817, 
        n2_adj_4818, n2_adj_4819, n2_adj_4820, n2_adj_4821, n2_adj_4822, 
        n2_adj_4823, n30086, n2_adj_4824, n2_adj_4825, n2_adj_4826, 
        n2_adj_4827, n2_adj_4828, n2_adj_4829, n2_adj_4830, n2_adj_4831, 
        n28339, n60244, n75167, n28341, n60243, n75145, n28443, 
        n28343, n60242, n75144, n30085, n28345, n60241, n75133, 
        n72465, n61378, n62336, n72466, n72464, n28347, n60240, 
        n75132, n2_adj_4832, n2_adj_4833, n2_adj_4834, n2_adj_4835, 
        n2_adj_4836, n2_adj_4837, n2_adj_4838, n2_adj_4839, n2_adj_4840, 
        n2_adj_4841, n2_adj_4842, n2_adj_4843, n2_adj_4844, n2_adj_4845, 
        n2_adj_4846, n28349, n60239, n75131, n67335, n2_adj_4847, 
        n28351, n60238, n75127, n30310, n79507, n75276, n28353, 
        n60237, n75124, n79141, n77369, n30084, n28355, n60236, 
        n75103, n30083, n2_adj_4848, n2_adj_4849, n28357, n60235, 
        n75100, n79390, n72529, n30082, n2_adj_4850, n67524, n67344, 
        n18_adj_4851, n28359, n60234, n75099, n66926, n16_adj_4852, 
        n30081, n61164, n66878, n20_adj_4853, n28361, n60233, n75092, 
        n28363, n60232, n75090, n67527, n67474, n69481, n67167, 
        n69703, \FRAME_MATCHER.i_31__N_2507 , n75063, n30080, n75064, 
        n2_adj_4854, n28365, n60231, n75084, n4_c, n67094, n75065, 
        n75068, n28367, n60230, n75083, n28369, n60229, n75082, 
        n28371, n60228, n75081, n28373, n60227, n75080, n28375, 
        n60226, n75076;
    wire [7:0]\data_in_frame[14]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30079, n2_adj_4855, n75069, n75073, n28377, n60225, n75075, 
        n30078, n28379, n60224, n6_adj_4856, n28381, n60223, n28383, 
        n60222, n28385, n60221, n28387, n60220, n28389, n60219;
    wire [31:0]n133;
    
    wire n161, n30077, n61294, n12_adj_4857, n30306, n30076;
    wire [7:0]\data_in_frame[19]_c ;   // verilog/coms.v(99[12:25])
    
    wire n29743, n67001, n30075, n30074, n16_adj_4858, n17, n30073, 
        n69880, n21_adj_4859;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    
    wire n30072, n30071, n30070, n67286, n20_adj_4860, n17_adj_4861, 
        n24_c, n62273, n30069, n67161, n8_adj_4862, n29980, n67438, 
        n12_adj_4863, n30068, n3_adj_4864, n30067, n67358, n6_adj_4865, 
        n67429, n67305, n67188, n61327, n10_adj_4866, n28692, n45, 
        n30066, n27159, n61384, n79372, n79366, n72550, n79360;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n79354, n79177, n7_adj_4868;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n79231, n79342, n79219, n79336, n79339, n26064, n67536, 
        n67347, n10_adj_4869, n66961, n79330;
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    
    wire n30775, n30065, n67593, n10_adj_4870, n67548, n66906, n30120, 
        n66935, n26480, n12_adj_4871, n30777, n8_adj_4872, n30778, 
        n30064, n37668, n30063, n67542, n67587, n6_adj_4873, n36341, 
        n67551, n10_adj_4874, n1130, n6_adj_4875, n79189, n72454, 
        n4_adj_4876, n67036, n30062, n14_adj_4877, n67400, n15_c, 
        n61380, n30004, n30009, n30014, n1168, n30097, n27213, 
        n67367, n67379, n10_adj_4878, n30060, n30061, n30017, n27058, 
        n33, n14_adj_4879, n10_adj_4880, n23, n1951, n4452, n1954, 
        n1957, n68793, n71998, \FRAME_MATCHER.i_31__N_2514 , n68593, 
        n66896, n67102, n10_adj_4883, n66948, n27006, n12_adj_4884, 
        n8_adj_4885, n72449, n72602, n72603, n72276, n72275, n72281, 
        n72282, n72300, n72299, n72455, n72456, n72582, n72581, 
        n72524, n72525, n72576, n72575, n72551, n72552, n72495, 
        n72494, n72554, n72555, n72468, n72467, n72563, n72564, 
        n72570, n72569, n72599, n72600, n72606, n72605, n1655, 
        n75282, n72501, n72502, n72500, n75279, n79111, n77433, 
        n1_adj_4886, n75196, n1699, n1193, n67397, n10_adj_4887, 
        n28400, n72507, n30043, n72508, n72506, n30042, n30041, 
        n30040, n30039, n30038, n67530, n30037, n30036, n30035, 
        n30034, n30033, n30032, n30031, n30030, n67355, n30029, 
        n30028, n30027, n30026, n30025, n30024, n30023, n30022, 
        n30021, n30020, n67533, n67590, n75273, n79642, n79165, 
        n77467, n79213, n7_adj_4888, n66957, n30300, n29992, n67004, 
        n77811, n79630, n30296, n29985;
    wire [7:0]control_mode_c;   // verilog/TinyFPGA_B.v(246[14:26])
    
    wire n29951;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n29944, n29942, n29940, n29939, n29938, n29935, n2_adj_4889;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n26197, n2_adj_4890, n2_adj_4891, n2_adj_4892, n2_adj_4893, 
        n2_adj_4894, n2_adj_4895, n2_adj_4896, n2_adj_4897, n2_adj_4898, 
        n2_adj_4899, n2_adj_4900, n2_adj_4901, n2_adj_4902, n2_adj_4903, 
        n2_adj_4904, n2_adj_4905, n2_adj_4906, n2_adj_4907, n2_adj_4908, 
        n2_adj_4909, n2_adj_4910, n2_adj_4911, n2_adj_4912, n2_adj_4913, 
        n26724, n79207, n7_adj_4914, n67016, n14_adj_4915, n20_adj_4916, 
        n18_adj_4917, n22_c, n69691, n67391, n16_adj_4918, n67545, 
        n17_adj_4919, n28325, n28676;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    
    wire n66088, n69308, n15_adj_4920, n2_adj_4921, n2_adj_4922, n2_adj_4923, 
        n12_adj_4924, n14_adj_4925, n68705, n2_adj_4926, n2_adj_4927, 
        n2_adj_4928, n8_adj_4929, n26813, n10_adj_4930, n26190, n26752, 
        n2_adj_4931, n2_adj_4932, n2_adj_4933, n27292, n34_c, n7_adj_4936, 
        n2_adj_4938, n2_adj_4939, n24_adj_4940, n38_adj_4941, n67313, 
        n36_adj_4942, n66092, n32, n40_adj_4943, n35_adj_4944, n75232, 
        n60595, n30774, n30773, n30772, n30770, n30768, n30766, 
        n30763, n30737, n30736, n30733, n30732, n30730, n30725, 
        n30723, n30722, n30699, n30681, n30679, n30665, n30664, 
        n30663, n30662, n30661, n30660, n30659, n30658, n30657;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n30656, n30655, n30654, n30653, n30652, n30651, n30650, 
        n30649;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n30648, n30647, n30646, n30645, n30644, n30643, n30642, 
        n30641;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n67249, n30640, n30639, n30638, n30637, n30636, n30635, 
        n30634, n30633, n30631, n30630, n30626, n30624, n29766, 
        n29769, n29772, n29776, n29779, n29782, n65834, n29788, 
        n65838, n30270, n30273, n30280, n30286, n30290, n30293, 
        n66022, n66068, n30323, n30326, n66112, n66144, n30339, 
        n30342, n30346, n30352, n30359, n2_adj_4947, n2_adj_4948, 
        n30378, n62342, n62473, n26551, n61016, n30385, n771, 
        \FRAME_MATCHER.i_31__N_2508 , n25859, n30402, n30405, n30408, 
        n30412, n15_adj_4949, n30418, n30422, n30425, n30445, n30448, 
        n2_adj_4950, n26345, n67043, n61494, n26053, n66130, n66084, 
        n66132, n29876, n29879, n66128, n67111, n26418, n29885;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    
    wire n29888, n26687, n26848, n9_adj_4951, n29891, n29894, n29897, 
        n29900, n29903, n29907, n29911, n29916, n29919, n67013, 
        n10_adj_4952, n29922, n29925, n35_adj_4953, n2_adj_4954, n28658, 
        n2_adj_4955, n2_adj_4956, n2_adj_4957, n2_adj_4958, n68795, 
        n29928, n29931, n2_adj_4959, n2_adj_4960, n26592, n10_adj_4961, 
        n79682, n27429, n2048, n2049, n20639, n65734, \FRAME_MATCHER.i_31__N_2512 , 
        n2060, n27432, n2_adj_4962, n2_adj_4963, n2_adj_4964, n2_adj_4965, 
        n2_adj_4966, n2_adj_4967, n2_adj_4968, n2_adj_4969, n2_adj_4970, 
        n2_adj_4971, n2_adj_4972, n2_adj_4973, n2_adj_4974, n2_adj_4975, 
        n2_adj_4976, n2_adj_4977, n26364, n71760, n67581, n66922, 
        n67129, n67441, n26721, n67456, n2_adj_4978, n2_adj_4979, 
        n2_adj_4980, n6_adj_4981, n2_adj_4982, n2_adj_4983, n2_adj_4984, 
        n2_adj_4985, n2_adj_4986, n2_adj_4987, n2_adj_4988, Kp_23__N_767, 
        n26986, n2_adj_4989, n2_adj_4990, n2_adj_4991, n2_adj_4992, 
        n2_adj_4993, n2_adj_4994, n2_adj_4995, n2_adj_4996, n2_adj_4997, 
        n44662, Kp_23__N_993, n67229, n2_adj_4998, n2_adj_4999, n2_adj_5000, 
        n2_adj_5001, n6_adj_5002, n2_adj_5003, n2_adj_5004, n2_adj_5005, 
        n2_adj_5006, n2_adj_5007, n2_adj_5008, n2_adj_5009, n2_adj_5010, 
        n2_adj_5011, n2_adj_5012, n2_adj_5013, n2_adj_5014, n3_adj_5015, 
        n66761, n66762, n66763, n66764, n66760, n66765, n3_adj_5016, 
        n66766, n66767, n29201;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n29195, n66768, n66769, n66770, n66758, n66759, n3_adj_5017, 
        n66771, n66772, n66773, n1_adj_5018, n66751, n1_adj_5019, 
        n66752, n2_adj_5020, n1_adj_5021, n66753, n1_adj_5022, n66754, 
        n1_adj_5023, n66749, n1_adj_5024, n66755, n1_adj_5025, n66756, 
        n2_adj_5026, n2_adj_5027, n1_adj_5028, n66750, n2_adj_5029, 
        n2_adj_5030, n6_adj_5032, n27164, n6_adj_5033, n62268, n6_adj_5034, 
        n59006, n66748, n59005, n59004, n59003, n59002, n59001, 
        n59000, n6_adj_5036, n62356, n71704, n27052, n67067, Kp_23__N_799, 
        n66860, n67338, n66868, n67412, n67554, n67105, n67462, 
        n27048, n26585, n10_adj_5037, n24270, n67560, n67406, n79528, 
        n26818, n26317, n27225, n26246, n26331, Kp_23__N_974, n26776, 
        n79159, n7_adj_5038, n6_adj_5040, n67468, n26959, n69576, 
        n24167, n67284, n67385, n67539, n67149, n67329, n67262, 
        n79522, n6_adj_5042, n72450, n77461, n77462, n79147, n79516, 
        n26783, n20634, n23017, n3303, n62383, n69522, n71754, 
        n67341, n67497, n61755, n67373, n72001, n71620, n69866, 
        n27045, n62404, n69568, n67301, n67170, n71938, n71942, 
        n71836, n66932, n71840, n62406, n71846, n67316, n67283, 
        n62365, n71852, n61366, n67382, n71858, n1955, n66893, 
        n61424, n67298, n67152, n71864, n67191, n67064, n69350, 
        n24227, n69224, n66970, n6_adj_5045, n69042, n66889, n67310, 
        n67246, n6_adj_5047, n5_adj_5049, n25879, n25749, n27994, 
        n67232, n69098, n67364, n71812, n25868, n26872, n66985, 
        n71818, n62266, n62313, n71824, n69062, n26796, n26292, 
        n25493, n71892, n71898, n67471, n69479, n71920, n69235, 
        n68596, n10_adj_5050, n25915, n79510, n16_adj_5051, n17_adj_5052, 
        n67569, n67422, n14_adj_5053, n62400, n25956, n62392, n26675, 
        n10_adj_5054, n10_adj_5055, n62348, n10_adj_5056, n14_adj_5057, 
        n25909, n20_adj_5058, n25779, n19_adj_5059, n72176, n61300, 
        n72057, n18_adj_5060, n6_adj_5061, n62329, n62003, n67488, 
        n67519, n68666, n62307, n66942, n67416, n71738, n71668, 
        n62327, n19_adj_5062, n14_adj_5063, n15_adj_5064, n69302, 
        n16_adj_5065, n17_adj_5066, n61404, n10_adj_5067, n61345, 
        n66854, n4_adj_5068, n4_adj_5069, n45392, n6_adj_5070, n69824, 
        n79183, n7_adj_5071, n67265, n6_adj_5072, n67028, n25507, 
        n6_adj_5073, n71966, n71970, n71974, n26261, n67563, n67566, 
        n71980, n67079, n61427, n67179, n67268, n67117, n27073, 
        n67091, n71948, n67322, n67114, n71954, n71766, n79504, 
        n67459, n62034, n26100, n18_adj_5074, n16_adj_5075, n30_adj_5076, 
        n20_adj_5077, n8_adj_5078, n66835, n69589, n7_adj_5079, n67225, 
        n67294, n62321, n26323, n67409, n7_adj_5081, n26655, n67032, 
        n71990, n71996, n67019, n67403, n25469, n71776, n7_adj_5082, 
        n71782, n69556, n67419, n4_adj_5083, n27_adj_5084, n71658, 
        n26779, n67198, n66918, n67099, n44_adj_5085, n35_adj_5086, 
        n66991, n26282, n72045, n27117, n67173, n24274, n26299, 
        n6_adj_5088, n26286, n26139, n67142, n69356, n10_adj_5089, 
        n62438, n67352, n6_adj_5090, n67146, n71590, n71596, n71600, 
        n71602, n71608, n67515, n71614, n71796, n68717, n66988, 
        n69802, n26296, n6_adj_5092, n66964, n14_adj_5093, n66974, 
        n15_adj_5094, n67465, n61339, n67070, n67185, n26718, n67182, 
        n71682, n71684, Kp_23__N_753, n71690, n66982, n71694, n71706, 
        n71712, n71700, n72487, n72485, n72486, n15_adj_5095, n14_adj_5096, 
        n69633, n69451, n72192, n69421, n24_adj_5097, n25, n23_adj_5098, 
        n10_adj_5099, n8_adj_5100, n71628, n10_adj_5101, n71630, n71632, 
        n69188, n8_adj_5102, n71636, n10_adj_5103, n71638, n71640, 
        n71642, n71908, n71644, n71916, n71646, n71648, n71886, 
        Kp_23__N_1607, n71650, n69696, n71654, n71568, n71656, n44_adj_5104, 
        n42_adj_5105, n43_adj_5106, n41_adj_5107, n40_adj_5108, n39, 
        n50, n45_adj_5109, n71502, n79456, n79228, n79216, n79441, 
        n79450, n79444, n79210, n79204, n79198, n79186, n79180, 
        n79174, n79438, n12_adj_5111, n10_adj_5112, n11, n79432, 
        n9_adj_5113, Kp_23__N_748, n67025, n79162, n66998, n10_adj_5114, 
        n23_adj_5115, n22_adj_5116, n27_adj_5117, n71866, n79156, 
        n79144, n79138, n26_adj_5118, n79132, n65, n29, n31, n75118, 
        n79108;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n29_adj_5120, n23_adj_5121;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n68353;
    
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30243));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30240));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15830_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [6]), 
            .I3(\Kp[6] ), .O(n30044));   // verilog/coms.v(130[12] 305[6])
    defparam i15830_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30237));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63516 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n79426));
    defparam byte_transmit_counter_0__bdd_4_lut_63516.LUT_INIT = 16'he4aa;
    SB_LUT4 n79426_bdd_4_lut (.I0(n79426), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n79429));
    defparam n79426_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4734), .S(n66744));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4735), .S(n66703));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30234));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_223_i3_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n67126), .I3(\data_out_frame[25] [6]), 
            .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_787_Select_222_i3_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_c), .I3(n62464), .O(n3_adj_4736));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63511 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n79420));
    defparam byte_transmit_counter_0__bdd_4_lut_63511.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_220_i3_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n67451), .I3(n62476), .O(n3_adj_4737));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i16106_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n30320));
    defparam i16106_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15831_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [5]), 
            .I3(\Kp[5] ), .O(n30045));   // verilog/coms.v(130[12] 305[6])
    defparam i15831_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_219_i3_3_lut (.I0(n61789), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n67055), .I3(GND_net), .O(n3_adj_4738));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_219_i3_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i15832_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [4]), 
            .I3(\Kp[4] ), .O(n30046));   // verilog/coms.v(130[12] 305[6])
    defparam i15832_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14181_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n28394));   // verilog/coms.v(109[34:55])
    defparam i14181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56621_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72477));
    defparam i56621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_218_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_4739), .I3(n67052), 
            .O(n3_adj_4740));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_218_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[23] [0]), .I1(n61954), .I2(GND_net), 
            .I3(GND_net), .O(n67052));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\data_out_frame[18] [5]), .I1(n62261), 
            .I2(GND_net), .I3(GND_net), .O(n67210));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut (.I0(n67480), .I1(n27298), .I2(n67139), .I3(\data_out_frame[22] [6]), 
            .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n61312), .I1(n14), .I2(n10_c), .I3(n67085), 
            .O(n61954));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i56622_4_lut (.I0(n72477), .I1(n28394), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n72478));
    defparam i56622_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n67716), .O(n79));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i56620_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72476));
    defparam i56620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15833_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [3]), 
            .I3(\Kp[3] ), .O(n30047));   // verilog/coms.v(130[12] 305[6])
    defparam i15833_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_out_frame[21] [0]), .I1(n25419), 
            .I2(GND_net), .I3(GND_net), .O(n67075));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i59751_2_lut (.I0(n79453), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n75296));
    defparam i59751_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut_adj_1080 (.I0(n67075), .I1(\data_out_frame[22] [7]), 
            .I2(n61422), .I3(n66953), .O(n18));
    defparam i7_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n27096), .I1(n18), .I2(n61954), .I3(n67210), 
            .O(n20));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i61651_3_lut (.I0(n79363), .I1(n79135), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n77507));
    defparam i61651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut (.I0(n61681), .I1(n20), .I2(n16_c), .I3(\data_out_frame[20] [7]), 
            .O(n67451));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(n62428), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n62464));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n67203), .I1(\data_out_frame[20] [5]), .I2(n67451), 
            .I3(n67485), .O(n10_adj_4741));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i16102_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[11]_c [6]), .O(n30316));
    defparam i16102_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(\data_out_frame[22] [7]), .I1(n67512), 
            .I2(GND_net), .I3(GND_net), .O(n67480));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut (.I0(n26999), .I1(n67572), .I2(\data_out_frame[23] [1]), 
            .I3(n67453), .O(n20_adj_4742));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1083 (.I0(n67277), .I1(\data_out_frame[21] [1]), 
            .I2(n26203), .I3(n67480), .O(n19));
    defparam i7_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1084 (.I0(n67210), .I1(\data_out_frame[23] [2]), 
            .I2(n26661), .I3(n61445), .O(n21));
    defparam i9_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut (.I0(n21), .I1(n19), .I2(n20_adj_4742), .I3(GND_net), 
            .O(n62290));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(n61789), .I1(n61412), .I2(n67126), .I3(GND_net), 
            .O(n8_c));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_217_i3_4_lut (.I0(n62368), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_c), .I3(n62290), .O(n3_adj_4743));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_217_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i15834_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [2]), 
            .I3(\Kp[2] ), .O(n30048));   // verilog/coms.v(130[12] 305[6])
    defparam i15834_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_216_i3_4_lut (.I0(n67061), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n67432), .I3(n62368), .O(n3_adj_4744));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_216_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [4]), 
            .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4745));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 select_1745_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_c));   // verilog/coms.v(148[4] 304[11])
    defparam select_1745_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1085 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_4746), .I3(n66848), .O(n27318));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1085.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [3]), 
            .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4747));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4748));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15835_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [1]), 
            .I3(\Kp[1] ), .O(n30049));   // verilog/coms.v(130[12] 305[6])
    defparam i15835_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4749));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4750));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n67055));
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4751));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut (.I0(n67055), .I1(n67435), .I2(\data_out_frame[25] [4]), 
            .I3(n26232), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1088 (.I0(\data_out_frame[25] [3]), .I1(n12), .I2(n67557), 
            .I3(\data_out_frame[25] [5]), .O(n62368));
    defparam i6_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1089 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[17] [7]), 
            .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4752));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1089.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4753));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4754));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15836_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n30050));   // verilog/coms.v(130[12] 305[6])
    defparam i15836_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1090 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[17] [4]), 
            .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4755));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'ha088;
    SB_DFFE data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30231));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_215_i3_4_lut (.I0(n62368), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_4756), .I3(n24045), .O(n3_adj_4757));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFE data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30228));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30225));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30222));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30219));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n29953));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4758));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30215));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30212));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30209));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30206));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30203));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30200));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30197));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4759));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15837_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11]_c [6]), 
            .I3(IntegralLimit[22]), .O(n30051));   // verilog/coms.v(130[12] 305[6])
    defparam i15837_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i30522_2_lut (.I0(LED_c), .I1(LED_N_3408), .I2(GND_net), .I3(GND_net), 
            .O(LED_N_3407));   // verilog/coms.v(253[15] 255[9])
    defparam i30522_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 select_787_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4760));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14997_4_lut (.I0(n2874), .I1(LED_N_3407), .I2(n27770), .I3(\FRAME_MATCHER.i_31__N_2513 ), 
            .O(n29211));   // verilog/coms.v(130[12] 305[6])
    defparam i14997_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i22968_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11]_c [5]), 
            .I3(IntegralLimit[21]), .O(n30052));   // verilog/coms.v(130[12] 305[6])
    defparam i22968_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_1743_Select_0_i3_3_lut (.I0(LED_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n3_adj_4761));   // verilog/coms.v(148[4] 304[11])
    defparam select_1743_Select_0_i3_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1091 (.I0(LED_c), .I1(n3_adj_4761), .I2(Kp_23__N_1748), 
            .I3(Kp_23__N_612), .O(n5_c));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1091.LUT_INIT = 16'hfcec;
    SB_LUT4 select_787_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4762));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
           .D(n29962));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15839_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11]_c [4]), 
            .I3(IntegralLimit[20]), .O(n30053));   // verilog/coms.v(130[12] 305[6])
    defparam i15839_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30193));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30190));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15840_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11]_c [3]), 
            .I3(IntegralLimit[19]), .O(n30054));   // verilog/coms.v(130[12] 305[6])
    defparam i15840_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30187));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4763));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30184));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30181));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n79420_bdd_4_lut (.I0(n79420), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n79423));
    defparam n79420_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4764));
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_213_i3_4_lut (.I0(n5_adj_4764), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n25458), .I3(n69352), .O(n3_adj_4765));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_213_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_787_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4766));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4767));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1093 (.I0(\FRAME_MATCHER.state[3] ), .I1(n62332), 
            .I2(\data_out_frame[24] [2]), .I3(\data_out_frame[24] [3]), 
            .O(n3_adj_4768));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1093.LUT_INIT = 16'h8228;
    SB_LUT4 select_787_Select_211_i3_4_lut (.I0(n24041), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n67132), .I3(n69736), .O(n3_adj_4769));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_211_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i4_4_lut_adj_1094 (.I0(n67503), .I1(\data_out_frame[24] [0]), 
            .I2(\data_out_frame[24] [1]), .I3(n67509), .O(n10_adj_4770));
    defparam i4_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4771));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30178));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_210_i3_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n10_adj_4770), .I3(n61447), 
            .O(n3_adj_4772));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(n26999), .I1(n61324), .I2(GND_net), 
            .I3(GND_net), .O(n66953));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1096 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[16] [4]), 
            .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4773));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1096.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4774));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut (.I0(n26619), .I1(n66953), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n61681));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4775));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1097 (.I0(n69543), .I1(\data_out_frame[20] [0]), 
            .I2(n67277), .I3(n62253), .O(n26829));
    defparam i1_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(n61681), .I1(n26517), .I2(GND_net), 
            .I3(GND_net), .O(n67176));
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1099 (.I0(n26829), .I1(n67158), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n69352));
    defparam i2_3_lut_adj_1099.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1100 (.I0(n62013), .I1(n67176), .I2(n26829), 
            .I3(n61333), .O(n12_adj_4776));
    defparam i5_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4777));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i6_4_lut_adj_1101 (.I0(n69502), .I1(n12_adj_4776), .I2(n67477), 
            .I3(\data_out_frame[22] [1]), .O(n69736));
    defparam i6_4_lut_adj_1101.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(n69736), .I1(n69352), .I2(GND_net), 
            .I3(GND_net), .O(n62332));
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4778));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4779));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4780));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23166_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11]_c [2]), 
            .I3(IntegralLimit[18]), .O(n30055));   // verilog/coms.v(130[12] 305[6])
    defparam i23166_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut (.I0(n61386), .I1(\data_out_frame[19] [5]), .I2(n61472), 
            .I3(GND_net), .O(n62253));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4781));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4782));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15842_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11]_c [1]), 
            .I3(IntegralLimit[17]), .O(n30056));   // verilog/coms.v(130[12] 305[6])
    defparam i15842_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1103 (.I0(n62285), .I1(n67252), .I2(n61824), 
            .I3(\data_out_frame[21] [7]), .O(n67509));
    defparam i3_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[23] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4783));
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1105 (.I0(n67509), .I1(n62253), .I2(n61503), 
            .I3(n6_adj_4783), .O(n24041));
    defparam i4_4_lut_adj_1105.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4784));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4785));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1106 (.I0(\data_out_frame[15] [3]), .I1(n67010), 
            .I2(n26089), .I3(GND_net), .O(n61386));
    defparam i2_3_lut_adj_1106.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4786));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1107 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[22] [0]), 
            .I2(n61386), .I3(GND_net), .O(n62285));
    defparam i2_3_lut_adj_1107.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26607));
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4787));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n67132));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1110 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[15] [0]), 
            .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n7));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1110.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n67058));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1112 (.I0(n67326), .I1(\data_out_frame[8] [6]), 
            .I2(n26060), .I3(n67388), .O(n10_adj_4788));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n66929), .I1(n10_adj_4788), .I2(\data_out_frame[6] [6]), 
            .I3(GND_net), .O(n26089));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut (.I0(\data_out_frame[15] [3]), .I1(n26645), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4789));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1113 (.I0(\data_out_frame[17] [5]), .I1(n67046), 
            .I2(n6_adj_4789), .I3(n26089), .O(n61362));
    defparam i1_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_out_frame[19] [3]), .I1(n61362), 
            .I2(GND_net), .I3(GND_net), .O(n67252));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i15843_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11]_c [0]), 
            .I3(IntegralLimit[16]), .O(n30057));   // verilog/coms.v(130[12] 305[6])
    defparam i15843_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16_4_lut (.I0(n61517), .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[14] [3]), 
            .I3(n67049), .O(n40_c));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(n67207), .I1(\data_out_frame[17] [7]), .I2(\data_out_frame[18] [2]), 
            .I3(\data_out_frame[19] [4]), .O(n38_c));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4790));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20_4_lut (.I0(n67252), .I1(n40_c), .I2(n30_c), .I3(n66967), 
            .O(n44));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4791));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18_4_lut (.I0(\data_out_frame[17] [0]), .I1(n69868), .I2(\data_out_frame[17] [5]), 
            .I3(\data_out_frame[17] [4]), .O(n42));
    defparam i18_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[19] [5]), .I1(n38_c), .I2(n26), 
            .I3(n67506), .O(n43));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(\data_out_frame[17] [3]), .I1(n27258), .I2(n62277), 
            .I3(\data_out_frame[17] [6]), .O(n41));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4792));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n67512));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1115 (.I0(n67280), .I1(n44_adj_4793), .I2(n27258), 
            .I3(n61320), .O(n14_adj_4794));
    defparam i6_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(n67512), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1117 (.I0(n9), .I1(n14_adj_4794), .I2(n67216), 
            .I3(n62302), .O(n61324));
    defparam i7_4_lut_adj_1117.LUT_INIT = 16'h9669;
    SB_LUT4 i15844_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n30058));   // verilog/coms.v(130[12] 305[6])
    defparam i15844_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_out_frame[18] [3]), .I1(n60995), 
            .I2(GND_net), .I3(GND_net), .O(n61422));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1119 (.I0(n61422), .I1(n26943), .I2(n67222), 
            .I3(n6_adj_4795), .O(n26517));
    defparam i4_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30175));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4796));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4797), .S(n29359));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4798));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15845_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12][6] ), 
            .I3(IntegralLimit[14]), .O(n30059));   // verilog/coms.v(130[12] 305[6])
    defparam i15845_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_1087_i1_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n4932[0]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_out_frame[20] [4]), .I1(n26517), 
            .I2(GND_net), .I3(GND_net), .O(n61434));
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n67506));
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 i15881_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [1]), 
            .I3(deadband[1]), .O(n30095));   // verilog/coms.v(130[12] 305[6])
    defparam i15881_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63506 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n79408));
    defparam byte_transmit_counter_0__bdd_4_lut_63506.LUT_INIT = 16'he4aa;
    SB_LUT4 n79408_bdd_4_lut (.I0(n79408), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n79411));
    defparam n79408_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1122 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n67491));
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h6666;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2068), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i15880_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n30094));   // verilog/coms.v(130[12] 305[6])
    defparam i15880_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66886));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i15879_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n30093));   // verilog/coms.v(130[12] 305[6])
    defparam i15879_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n28131), 
            .D(n4932[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1124 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(GND_net), .I3(GND_net), .O(n67046));
    defparam i1_2_lut_adj_1124.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4799), .S(n66700));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i21586_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n30092));   // verilog/coms.v(130[12] 305[6])
    defparam i21586_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30172));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4800));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1125 (.I0(n66886), .I1(\data_out_frame[15] [7]), 
            .I2(n8), .I3(n67491), .O(n7_adj_4802));
    defparam i1_4_lut_adj_1125.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1126 (.I0(n67425), .I1(n7_adj_4802), .I2(n62080), 
            .I3(n8_adj_4803), .O(n61333));
    defparam i5_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1127 (.I0(\data_out_frame[18] [1]), .I1(n67425), 
            .I2(n67271), .I3(n67222), .O(n69502));
    defparam i3_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4804));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63496 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n79402));
    defparam byte_transmit_counter_0__bdd_4_lut_63496.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1128 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [0]), 
            .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4805));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1128.LUT_INIT = 16'ha088;
    SB_LUT4 i59716_2_lut (.I0(n79435), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n75277));
    defparam i59716_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15877_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16]_c [5]), 
            .I3(deadband[5]), .O(n30091));   // verilog/coms.v(130[12] 305[6])
    defparam i15877_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i61489_3_lut (.I0(n79375), .I1(n79201), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n77345));
    defparam i61489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15876_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16]_c [6]), 
            .I3(deadband[6]), .O(n30090));   // verilog/coms.v(130[12] 305[6])
    defparam i15876_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4806));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15875_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16][7] ), 
            .I3(deadband[7]), .O(n30089));   // verilog/coms.v(130[12] 305[6])
    defparam i15875_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4807));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n79402_bdd_4_lut (.I0(n79402), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n79405));
    defparam n79402_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14179_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n28392));   // verilog/coms.v(109[34:55])
    defparam i14179_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30169));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15874_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n30088));   // verilog/coms.v(130[12] 305[6])
    defparam i15874_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63491 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n79396));
    defparam byte_transmit_counter_0__bdd_4_lut_63491.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4808), .S(n66699));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1129 (.I0(n67332), .I1(\data_out_frame[22] [2]), 
            .I2(\data_out_frame[20] [0]), .I3(n67506), .O(n10_adj_4809));
    defparam i4_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1130 (.I0(n67010), .I1(n10_adj_4809), .I2(\data_out_frame[17] [6]), 
            .I3(GND_net), .O(n68641));
    defparam i5_3_lut_adj_1130.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1131 (.I0(n68641), .I1(n26619), .I2(n24023), 
            .I3(GND_net), .O(n8_adj_4810));
    defparam i3_3_lut_adj_1131.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_adj_1132 (.I0(\data_out_frame[22] [1]), .I1(n61324), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4811));
    defparam i2_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_33_lut  (.I0(n75190), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n60249), .O(n28327)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_32_lut  (.I0(n75189), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n60248), .O(n28329)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_32  (.CI(n60248), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n60249));
    SB_LUT4 n79396_bdd_4_lut (.I0(n79396), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n79399));
    defparam n79396_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_31_lut  (.I0(n75181), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n60247), .O(n28331)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_31  (.CI(n60247), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n60248));
    SB_LUT4 i2_4_lut (.I0(n61434), .I1(n7_adj_4811), .I2(\data_out_frame[21] [7]), 
            .I3(n8_adj_4810), .O(n67158));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4812));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1133 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [4]), 
            .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n6_adj_4813));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1133.LUT_INIT = 16'ha088;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_30_lut  (.I0(n75171), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n60246), .O(n28333)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_30  (.CI(n60246), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n60247));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_29_lut  (.I0(n75168), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n60245), .O(n28337)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_787_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4814));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_4_lut (.I0(n72460), .I1(n72458), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[0]), 
            .O(n7_adj_4815));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15873_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n30087));   // verilog/coms.v(130[12] 305[6])
    defparam i15873_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(n61447), .I1(n61577), .I2(GND_net), 
            .I3(GND_net), .O(n67291));
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i59793_2_lut (.I0(n79459), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n75267));
    defparam i59793_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4816), .S(n66577));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4817), .S(n66698));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4818), .S(n66697));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4819), .S(n66696));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4820), .S(n66695));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4821), .S(n66694));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4822), .S(n27));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4823), .S(n66693));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15872_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n30086));   // verilog/coms.v(130[12] 305[6])
    defparam i15872_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4824), .S(n66692));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4825), .S(n66691));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4826), .S(n66690));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4827), .S(n66689));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4828), .S(n66688));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4829), .S(n66687));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4830), .S(n66686));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4831), .S(n66685));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_29  (.CI(n60245), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n60246));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_28_lut  (.I0(n75167), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n60244), .O(n28339)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_28  (.CI(n60244), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n60245));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_27_lut  (.I0(n75145), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n60243), .O(n28341)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i14230_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n28443));   // verilog/coms.v(109[34:55])
    defparam i14230_2_lut.LUT_INIT = 16'hbbbb;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_27  (.CI(n60243), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n60244));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_26_lut  (.I0(n75144), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n60242), .O(n28343)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_26  (.CI(n60242), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n60243));
    SB_LUT4 i15871_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n30085));   // verilog/coms.v(130[12] 305[6])
    defparam i15871_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_25_lut  (.I0(n75133), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n60241), .O(n28345)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i56609_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72465));
    defparam i56609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1135 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n61378), .I3(GND_net), .O(n61445));
    defparam i2_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_25  (.CI(n60241), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n60242));
    SB_LUT4 i1_2_lut_adj_1136 (.I0(\data_out_frame[16] [1]), .I1(n61445), 
            .I2(GND_net), .I3(GND_net), .O(n62336));
    defparam i1_2_lut_adj_1136.LUT_INIT = 16'h6666;
    SB_LUT4 i56610_4_lut (.I0(n72465), .I1(n28443), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][0] ), .O(n72466));
    defparam i56610_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i56608_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72464));
    defparam i56608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_24_lut  (.I0(n75132), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n60240), .O(n28347)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_24  (.CI(n60240), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n60241));
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4832), .S(n66684));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4833), .S(n66683));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4834), .S(n66682));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4835), .S(n66681));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4836), .S(n66680));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4837), .S(n66679));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4838), .S(n66678));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4839), .S(n66677));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4840), .S(n66676));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4841), .S(n66675));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4842), .S(n66674));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4843), .S(n66673));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4844), .S(n66672));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4845), .S(n66671));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4846), .S(n66670));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_23_lut  (.I0(n75131), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n60239), .O(n28349)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_23  (.CI(n60239), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n60240));
    SB_LUT4 i1_2_lut_adj_1137 (.I0(\data_out_frame[17] [5]), .I1(n26645), 
            .I2(GND_net), .I3(GND_net), .O(n67335));
    defparam i1_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4847), .S(n66669));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_22_lut  (.I0(n75127), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n60238), .O(n28351)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_22  (.CI(n60238), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n60239));
    SB_LUT4 i16096_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[11]_c [4]), .O(n30310));
    defparam i16096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i59756_2_lut (.I0(n79507), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n75276));
    defparam i59756_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_21_lut  (.I0(n75124), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n60237), .O(n28353)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_21  (.CI(n60237), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n60238));
    SB_LUT4 i61513_3_lut (.I0(n79405), .I1(n79141), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n77369));
    defparam i61513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21967_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n30084));   // verilog/coms.v(130[12] 305[6])
    defparam i21967_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_20_lut  (.I0(n75103), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n60236), .O(n28355)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i15869_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15][5] ), 
            .I3(deadband[13]), .O(n30083));   // verilog/coms.v(130[12] 305[6])
    defparam i15869_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26619));
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4848), .S(n66668));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30166));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_20  (.CI(n60236), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n60237));
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4849), .S(n66667));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_19_lut  (.I0(n75100), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n60235), .O(n28357)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63486 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n79390));
    defparam byte_transmit_counter_0__bdd_4_lut_63486.LUT_INIT = 16'he4aa;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_19  (.CI(n60235), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n60236));
    SB_LUT4 n79390_bdd_4_lut (.I0(n79390), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n72529));
    defparam n79390_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15868_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n30082));   // verilog/coms.v(130[12] 305[6])
    defparam i15868_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1139 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [2]), 
            .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4850));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1139.LUT_INIT = 16'ha088;
    SB_LUT4 i7_4_lut_adj_1140 (.I0(n67524), .I1(n67344), .I2(\data_out_frame[12] [0]), 
            .I3(\data_out_frame[10] [7]), .O(n18_adj_4851));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_18_lut  (.I0(n75099), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n60234), .O(n28359)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_18  (.CI(n60234), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n60235));
    SB_LUT4 i5_2_lut (.I0(n66926), .I1(\data_out_frame[6] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4852));   // verilog/coms.v(74[16:27])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15867_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n30081));   // verilog/coms.v(130[12] 305[6])
    defparam i15867_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9_4_lut_adj_1141 (.I0(n61164), .I1(n18_adj_4851), .I2(\data_out_frame[13] [7]), 
            .I3(n66878), .O(n20_adj_4853));   // verilog/coms.v(74[16:27])
    defparam i9_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_17_lut  (.I0(n75092), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n60233), .O(n28361)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_17  (.CI(n60233), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n60234));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_16_lut  (.I0(n75090), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n60232), .O(n28363)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i10_4_lut_adj_1142 (.I0(n67527), .I1(n20_adj_4853), .I2(n16_adj_4852), 
            .I3(n67474), .O(n69481));   // verilog/coms.v(74[16:27])
    defparam i10_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1143 (.I0(\data_out_frame[12] [3]), .I1(n69481), 
            .I2(n67474), .I3(n67167), .O(n69703));
    defparam i3_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i59481_2_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75063));   // verilog/coms.v(158[12:15])
    defparam i59481_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15866_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n30080));   // verilog/coms.v(130[12] 305[6])
    defparam i15866_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i59835_2_lut (.I0(\FRAME_MATCHER.i[2] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75064));   // verilog/coms.v(158[12:15])
    defparam i59835_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4854), .S(n66666));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_16  (.CI(n60232), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n60233));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_15_lut  (.I0(n75084), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n60231), .O(n28365)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i2_4_lut_adj_1144 (.I0(n25421), .I1(n4_c), .I2(n69703), .I3(n67094), 
            .O(n44_adj_4793));   // verilog/coms.v(77[16:27])
    defparam i2_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i59485_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75065));   // verilog/coms.v(158[12:15])
    defparam i59485_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i59552_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75068));   // verilog/coms.v(158[12:15])
    defparam i59552_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_15  (.CI(n60231), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n60232));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_14_lut  (.I0(n75083), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n60230), .O(n28367)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_out_frame[16] [3]), .I1(n44_adj_4793), 
            .I2(GND_net), .I3(GND_net), .O(n27096));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_14  (.CI(n60230), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n60231));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_13_lut  (.I0(n75082), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n60229), .O(n28369)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30163));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_13  (.CI(n60229), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n60230));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_12_lut  (.I0(n75081), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n60228), .O(n28371)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_12  (.CI(n60228), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n60229));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_11_lut  (.I0(n75080), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n60227), .O(n28373)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_11  (.CI(n60227), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n60228));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_10_lut  (.I0(n75076), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n60226), .O(n28375)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i22175_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14]_c [1]), 
            .I3(deadband[17]), .O(n30079));   // verilog/coms.v(130[12] 305[6])
    defparam i22175_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_10  (.CI(n60226), .I0(n28651), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n60227));
    SB_DFFE data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30160));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1146 (.I0(\data_out_frame[19] [0]), .I1(n62261), 
            .I2(GND_net), .I3(GND_net), .O(n67280));
    defparam i1_2_lut_adj_1146.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4855));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59486_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75069));   // verilog/coms.v(158[12:15])
    defparam i59486_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30157));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59553_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75073));   // verilog/coms.v(158[12:15])
    defparam i59553_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_9_lut  (.I0(n75075), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n60225), .O(n28377)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i59556_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75075));   // verilog/coms.v(158[12:15])
    defparam i59556_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30154));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_9  (.CI(n60225), .I0(n28651), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n60226));
    SB_LUT4 i15864_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][2] ), 
            .I3(deadband[18]), .O(n30078));   // verilog/coms.v(130[12] 305[6])
    defparam i15864_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_8_lut  (.I0(n75073), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n60224), .O(n28379)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30151));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_8  (.CI(n60224), .I0(n28651), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n60225));
    SB_LUT4 i4_4_lut_adj_1147 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[18] [0]), 
            .I2(n67335), .I3(n6_adj_4856), .O(n62013));
    defparam i4_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_7_lut  (.I0(n75069), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n60223), .O(n28381)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4855), .S(n66665));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_7  (.CI(n60223), .I0(n28651), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n60224));
    SB_LUT4 i1_4_lut_adj_1148 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[22] [4]), 
            .I2(\data_out_frame[22] [3]), .I3(n62013), .O(n67274));
    defparam i1_4_lut_adj_1148.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30148));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_6_lut  (.I0(n75068), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n60222), .O(n28383)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_6  (.CI(n60222), .I0(n28651), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n60223));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_5_lut  (.I0(n75065), .I1(n28651), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n60221), .O(n28385)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_5  (.CI(n60221), .I0(n28651), .I1(\FRAME_MATCHER.i [3]), 
            .CO(n60222));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_4_lut  (.I0(n75064), .I1(n28651), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n60220), .O(n28387)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i59834_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75076));   // verilog/coms.v(158[12:15])
    defparam i59834_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_4  (.CI(n60220), .I0(n28651), .I1(\FRAME_MATCHER.i[2] ), 
            .CO(n60221));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_3_lut  (.I0(n75063), .I1(n28651), 
            .I2(\FRAME_MATCHER.i[1] ), .I3(n60219), .O(n28389)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_3  (.CI(n60219), .I0(n28651), .I1(\FRAME_MATCHER.i[1] ), 
            .CO(n60220));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i[0] ), 
            .CO(n60219));
    SB_LUT4 i59500_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75080));   // verilog/coms.v(158[12:15])
    defparam i59500_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i19832_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14]_c [3]), 
            .I3(deadband[19]), .O(n30077));   // verilog/coms.v(130[12] 305[6])
    defparam i19832_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1149 (.I0(\data_out_frame[20] [7]), .I1(n27096), 
            .I2(n61294), .I3(n62281), .O(n12_adj_4857));
    defparam i5_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1150 (.I0(\data_out_frame[21] [1]), .I1(n12_adj_4857), 
            .I2(n67280), .I3(n62302), .O(n62428));
    defparam i6_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i16092_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[11]_c [3]), .O(n30306));
    defparam i16092_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1151 (.I0(\data_out_frame[20] [6]), .I1(n25419), 
            .I2(\data_out_frame[20] [5]), .I3(GND_net), .O(n61312));
    defparam i2_3_lut_adj_1151.LUT_INIT = 16'h9696;
    SB_LUT4 i59534_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75081));   // verilog/coms.v(158[12:15])
    defparam i59534_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15862_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][4] ), 
            .I3(deadband[20]), .O(n30076));   // verilog/coms.v(130[12] 305[6])
    defparam i15862_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i59867_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75082));   // verilog/coms.v(158[12:15])
    defparam i59867_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26203));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i15529_3_lut (.I0(\data_in_frame[19]_c [1]), .I1(rx_data[1]), 
            .I2(n69075), .I3(GND_net), .O(n29743));   // verilog/coms.v(130[12] 305[6])
    defparam i15529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59541_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75083));   // verilog/coms.v(158[12:15])
    defparam i59541_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1153 (.I0(n62336), .I1(n67001), .I2(n44_adj_4793), 
            .I3(\data_out_frame[16] [2]), .O(n60995));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1153.LUT_INIT = 16'h9669;
    SB_LUT4 i15861_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][5] ), 
            .I3(deadband[21]), .O(n30075));   // verilog/coms.v(130[12] 305[6])
    defparam i15861_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i59542_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75084));   // verilog/coms.v(158[12:15])
    defparam i59542_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1154 (.I0(\data_out_frame[22] [6]), .I1(n69543), 
            .I2(GND_net), .I3(GND_net), .O(n67485));
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1155 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [0]), 
            .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4854));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1155.LUT_INIT = 16'ha088;
    SB_LUT4 i15860_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][6] ), 
            .I3(deadband[22]), .O(n30074));   // verilog/coms.v(130[12] 305[6])
    defparam i15860_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1156 (.I0(n61362), .I1(n62285), .I2(n61503), 
            .I3(\data_out_frame[21] [6]), .O(n67477));
    defparam i3_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1157 (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[21] [0]), 
            .I2(n67477), .I3(n67485), .O(n16_adj_4858));
    defparam i6_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1158 (.I0(n61312), .I1(n62428), .I2(\data_out_frame[22] [5]), 
            .I3(n67274), .O(n17));
    defparam i7_4_lut_adj_1158.LUT_INIT = 16'h9669;
    SB_LUT4 i59554_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75090));   // verilog/coms.v(158[12:15])
    defparam i59554_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15859_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][7] ), 
            .I3(deadband[23]), .O(n30073));   // verilog/coms.v(130[12] 305[6])
    defparam i15859_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i59740_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75092));   // verilog/coms.v(158[12:15])
    defparam i59740_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i9_4_lut_adj_1159 (.I0(n17), .I1(n67291), .I2(n16_adj_4858), 
            .I3(n67158), .O(n69880));
    defparam i9_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1160 (.I0(\data_out_frame[23] [7]), .I1(n67058), 
            .I2(n26232), .I3(\data_out_frame[24] [3]), .O(n21_adj_4859));
    defparam i8_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i15858_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n30072));   // verilog/coms.v(130[12] 305[6])
    defparam i15858_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15857_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13][2] ), 
            .I3(IntegralLimit[2]), .O(n30071));   // verilog/coms.v(130[12] 305[6])
    defparam i15857_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15856_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n30070));   // verilog/coms.v(130[12] 305[6])
    defparam i15856_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_3_lut (.I0(\data_out_frame[23] [5]), .I1(n67286), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n20_adj_4860));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut (.I0(n21_adj_4859), .I1(n17_adj_4861), .I2(n67132), 
            .I3(n69880), .O(n24_c));
    defparam i11_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut (.I0(n26607), .I1(n24_c), .I2(n20_adj_4860), .I3(\data_out_frame[24] [7]), 
            .O(n62273));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4850), .S(n66664));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i19636_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13][4] ), 
            .I3(IntegralLimit[4]), .O(n30069));   // verilog/coms.v(130[12] 305[6])
    defparam i19636_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30145));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_out_frame[22] [4]), .I1(n24023), 
            .I2(GND_net), .I3(GND_net), .O(n67161));
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(n67557), .I1(n24041), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4862));
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
           .D(n29980));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1163 (.I0(n67161), .I1(n67438), .I2(\data_out_frame[25] [7]), 
            .I3(n62273), .O(n12_adj_4863));
    defparam i5_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i15854_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13][5] ), 
            .I3(IntegralLimit[5]), .O(n30068));   // verilog/coms.v(130[12] 305[6])
    defparam i15854_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_209_i3_4_lut (.I0(n62332), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_4863), .I3(n8_adj_4862), .O(n3_adj_4864));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i15853_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13][6] ), 
            .I3(IntegralLimit[6]), .O(n30067));   // verilog/coms.v(130[12] 305[6])
    defparam i15853_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30141));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1164 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[10] [5]), 
            .I2(n67358), .I3(n6_adj_4865), .O(n26645));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1165 (.I0(\data_out_frame[17] [2]), .I1(n67429), 
            .I2(GND_net), .I3(GND_net), .O(n67305));
    defparam i1_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30138));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1166 (.I0(\data_out_frame[17] [3]), .I1(n67188), 
            .I2(n26645), .I3(n61327), .O(n61472));
    defparam i3_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67049));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1168 (.I0(n10_adj_4866), .I1(n67716), .I2(n8_adj_5), 
            .I3(GND_net), .O(n28692));
    defparam i2_3_lut_adj_1168.LUT_INIT = 16'hfbfb;
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30135));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1169 (.I0(n45), .I1(\data_out_frame[13] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(\data_out_frame[15] [1]), .O(n67429));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i15852_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13][7] ), 
            .I3(IntegralLimit[7]), .O(n30066));   // verilog/coms.v(130[12] 305[6])
    defparam i15852_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1170 (.I0(n27159), .I1(n67429), .I2(n67049), 
            .I3(n61384), .O(n61824));
    defparam i3_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63481 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n79372));
    defparam byte_transmit_counter_0__bdd_4_lut_63481.LUT_INIT = 16'he4aa;
    SB_LUT4 n79372_bdd_4_lut (.I0(n79372), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n79375));
    defparam n79372_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63467 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n79366));
    defparam byte_transmit_counter_0__bdd_4_lut_63467.LUT_INIT = 16'he4aa;
    SB_LUT4 n79366_bdd_4_lut (.I0(n79366), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n72550));
    defparam n79366_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63462 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n79360));
    defparam byte_transmit_counter_0__bdd_4_lut_63462.LUT_INIT = 16'he4aa;
    SB_LUT4 n79360_bdd_4_lut (.I0(n79360), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n79363));
    defparam n79360_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63581 (.I0(byte_transmit_counter_c[3]), 
            .I1(n77369), .I2(n75276), .I3(byte_transmit_counter_c[4]), 
            .O(n79354));
    defparam byte_transmit_counter_3__bdd_4_lut_63581.LUT_INIT = 16'he4aa;
    SB_LUT4 n79354_bdd_4_lut (.I0(n79354), .I1(n79177), .I2(n7_adj_4868), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[0]));
    defparam n79354_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63452 (.I0(byte_transmit_counter_c[3]), 
            .I1(n79231), .I2(n75267), .I3(byte_transmit_counter_c[4]), 
            .O(n79342));
    defparam byte_transmit_counter_3__bdd_4_lut_63452.LUT_INIT = 16'he4aa;
    SB_LUT4 n79342_bdd_4_lut (.I0(n79342), .I1(n79219), .I2(n7_adj_4815), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[7]));
    defparam n79342_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63457 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n79336));
    defparam byte_transmit_counter_0__bdd_4_lut_63457.LUT_INIT = 16'he4aa;
    SB_LUT4 n79336_bdd_4_lut (.I0(n79336), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n79339));
    defparam n79336_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1171 (.I0(\data_out_frame[19] [4]), .I1(n61472), 
            .I2(n67305), .I3(n27159), .O(n61503));
    defparam i1_4_lut_adj_1171.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n67503));
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1173 (.I0(n26064), .I1(n26060), .I2(n67536), 
            .I3(GND_net), .O(n67524));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1173.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26661));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1175 (.I0(n67347), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[7] [7]), .I3(n67524), .O(n10_adj_4869));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30132));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1176 (.I0(\data_out_frame[8] [4]), .I1(n10_adj_4869), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n61327));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1177 (.I0(n61327), .I1(n66961), .I2(\data_out_frame[16] [7]), 
            .I3(GND_net), .O(n61384));
    defparam i2_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63442 (.I0(byte_transmit_counter_c[3]), 
            .I1(n77345), .I2(n75277), .I3(byte_transmit_counter_c[4]), 
            .O(n79330));
    defparam byte_transmit_counter_3__bdd_4_lut_63442.LUT_INIT = 16'he4aa;
    SB_LUT4 i23518_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n23094), .I3(GND_net), .O(n30775));
    defparam i23518_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30129));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1178 (.I0(n27258), .I1(n61320), .I2(GND_net), 
            .I3(GND_net), .O(n62281));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n67344));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i15851_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n30065));   // verilog/coms.v(130[12] 305[6])
    defparam i15851_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1180 (.I0(n67593), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(n67599), .O(n10_adj_4870));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30126));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1181 (.I0(n67548), .I1(n10_adj_4870), .I2(\data_out_frame[9] [7]), 
            .I3(GND_net), .O(n66906));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1182 (.I0(n66906), .I1(n67344), .I2(\data_out_frame[14] [4]), 
            .I3(GND_net), .O(n27258));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1182.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30123));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30120));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1183 (.I0(n66935), .I1(n67361), .I2(\data_out_frame[12] [1]), 
            .I3(n26480), .O(n12_adj_4871));   // verilog/coms.v(77[16:27])
    defparam i5_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i23513_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n23094), .I3(GND_net), .O(n30777));
    defparam i23513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1184 (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[9] [4]), 
            .I2(n12_adj_4871), .I3(n8_adj_4872), .O(n61320));
    defparam i1_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i23517_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n23094), .I3(GND_net), .O(n30778));
    defparam i23517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15850_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n30064));   // verilog/coms.v(130[12] 305[6])
    defparam i15850_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67388));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i23519_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n23094), .I3(GND_net), .O(n37668));
    defparam i23519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22689_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12][2] ), 
            .I3(IntegralLimit[10]), .O(n30063));   // verilog/coms.v(130[12] 305[6])
    defparam i22689_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1186 (.I0(n67542), .I1(n67388), .I2(n67587), 
            .I3(n6_adj_4873), .O(n67271));
    defparam i4_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1187 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n36341));   // verilog/coms.v(100[12:26])
    defparam i5_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1188 (.I0(n67536), .I1(n66929), .I2(n36341), 
            .I3(n67551), .O(n10_adj_4874));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1189 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(n1130), .I3(\data_out_frame[13] [2]), .O(n67326));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4875));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 n79330_bdd_4_lut (.I0(n79330), .I1(n79189), .I2(n72454), .I3(byte_transmit_counter_c[4]), 
            .O(tx_data[3]));
    defparam n79330_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1191 (.I0(\data_out_frame[11] [2]), .I1(n4_adj_4876), 
            .I2(n67036), .I3(n6_adj_4875), .O(n67542));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i22645_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12][3] ), 
            .I3(IntegralLimit[11]), .O(n30062));   // verilog/coms.v(130[12] 305[6])
    defparam i22645_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_3_lut_adj_1192 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[8] [4]), 
            .I2(n67326), .I3(GND_net), .O(n14_adj_4877));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1193 (.I0(n67542), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[6] [3]), .I3(n67400), .O(n15_c));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1194 (.I0(n15_c), .I1(\data_out_frame[10] [6]), 
            .I2(n14_adj_4877), .I3(\data_out_frame[4] [2]), .O(n1720));   // verilog/coms.v(77[16:43])
    defparam i8_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_out_frame[13] [0]), .I1(n45), .I2(GND_net), 
            .I3(GND_net), .O(n61380));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
           .D(n30004));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
           .D(n30009));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
           .D(n30014));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_out_frame[7] [0]), .I1(n1168), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4876));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i8_2_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30097));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1197 (.I0(n27213), .I1(n67367), .I2(\data_out_frame[11] [4]), 
            .I3(n67379), .O(n10_adj_4878));
    defparam i4_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i15846_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12][5] ), 
            .I3(IntegralLimit[13]), .O(n30060));   // verilog/coms.v(130[12] 305[6])
    defparam i15846_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9_2_lut (.I0(PWMLimit[17]), .I1(n462), .I2(GND_net), .I3(GND_net), 
            .O(n36361));
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i22646_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12][4] ), 
            .I3(IntegralLimit[12]), .O(n30061));   // verilog/coms.v(130[12] 305[6])
    defparam i22646_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
           .D(n30017));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n30095), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n30094), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1198 (.I0(n67036), .I1(n27058), .I2(\data_out_frame[9] [2]), 
            .I3(n33), .O(n14_adj_4879));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1199 (.I0(\data_out_frame[13] [4]), .I1(n14_adj_4879), 
            .I2(n10_adj_4880), .I3(\data_out_frame[9] [0]), .O(n62080));   // verilog/coms.v(88[17:70])
    defparam i7_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n67036));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1201 (.I0(n105), .I1(n23), .I2(control_mode[0]), 
            .I3(control_update), .O(n24));
    defparam i3_4_lut_adj_1201.LUT_INIT = 16'hefff;
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n30093), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67367));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut (.I0(n1951), .I1(n4452), .I2(n1954), .I3(n1957), 
            .O(n68793));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1951), .I1(n4452), .I2(n71998), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n68593));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i4_4_lut_adj_1203 (.I0(n30), .I1(n66896), .I2(\data_out_frame[9] [4]), 
            .I3(n67102), .O(n10_adj_4883));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n30092), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1204 (.I0(\data_out_frame[6] [7]), .I1(n10_adj_4883), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n61164));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1204.LUT_INIT = 16'h9696;
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n30091), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n30090), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n30089), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n30088), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n30087), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66896));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n30086), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1206 (.I0(n66896), .I1(n66948), .I2(\data_out_frame[9] [1]), 
            .I3(n27006), .O(n12_adj_4884));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1207 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(n12_adj_4884), .I3(n8_adj_4885), .O(n27184));
    defparam i1_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n30085), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n30084), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56593_4_lut (.I0(\data_out_frame[0][4] ), .I1(\data_out_frame[3][4] ), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n72449));
    defparam i56593_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i56746_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72602));
    defparam i56746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56747_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72603));
    defparam i56747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56420_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72276));
    defparam i56420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56419_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72275));
    defparam i56419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56425_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72281));
    defparam i56425_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n30083), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n30082), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56426_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72282));
    defparam i56426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56444_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72300));
    defparam i56444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56443_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72299));
    defparam i56443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56599_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72455));
    defparam i56599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56600_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72456));
    defparam i56600_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n30081), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n30080), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n30079), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n30078), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n30077), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56726_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72582));
    defparam i56726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56725_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72581));
    defparam i56725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56668_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72524));
    defparam i56668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56669_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72525));
    defparam i56669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56720_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72576));
    defparam i56720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56719_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72575));
    defparam i56719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56695_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72551));
    defparam i56695_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n30076), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56696_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72552));
    defparam i56696_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n30075), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n30074), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n30073), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56639_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72495));
    defparam i56639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56638_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72494));
    defparam i56638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56698_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72554));
    defparam i56698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56699_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72555));
    defparam i56699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56612_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72468));
    defparam i56612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56611_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72467));
    defparam i56611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56707_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72563));
    defparam i56707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56708_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72564));
    defparam i56708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56714_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72570));
    defparam i56714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56713_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72569));
    defparam i56713_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n30072), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n30071), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n30070), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56743_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72599));
    defparam i56743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56744_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72600));
    defparam i56744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56750_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72606));
    defparam i56750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56749_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72605));
    defparam i56749_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n30069), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n30068), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n30067), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1208 (.I0(\data_out_frame[14] [5]), .I1(n1655), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n66961));
    defparam i2_3_lut_adj_1208.LUT_INIT = 16'h9696;
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n30066), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n30065), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n30064), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59647_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n75282));
    defparam i59647_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i56645_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72501));
    defparam i56645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56646_4_lut (.I0(n72501), .I1(n75282), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n72502));
    defparam i56646_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i56644_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72500));
    defparam i56644_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n30063), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59778_2_lut (.I0(n79429), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n75279));
    defparam i59778_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n30062), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i61577_3_lut (.I0(n79399), .I1(n79111), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n77433));
    defparam i61577_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n30061), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67188));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n30060), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n30059), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n30058), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n30057), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n30056), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4814), .S(n66663));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_4886));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59759_2_lut (.I0(\data_out_frame[3][3] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n75196));
    defparam i59759_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2874), .D(n6_adj_4813), .S(n66662));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4812), .S(n66661));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n30055), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4807), .S(n66660));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4806), .S(n66659));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n30054), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4805), .S(n66658));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4804), .S(n66657));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n30053), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n30052), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n30051), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n30050), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n30049), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4800), .S(n66656));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n30048), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n30047), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n30046), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n30045), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n30044), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4798), .S(n66655));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4796), .S(n66654));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1210 (.I0(n1193), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[14] [7]), .I3(n67397), .O(n10_adj_4887));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4792), .S(n66653));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4791), .S(n66652));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14187_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n28400));   // verilog/coms.v(109[34:55])
    defparam i14187_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4790), .S(n66651));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56651_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72507));
    defparam i56651_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n30043), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56652_4_lut (.I0(n72507), .I1(n28400), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n72508));
    defparam i56652_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i56650_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72506));
    defparam i56650_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n30042), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n30041), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2874), .D(n7), .S(n66650));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1211 (.I0(\data_out_frame[8] [1]), .I1(n10_adj_4887), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n67347));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_adj_1211.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4787), .S(n66649));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n30040), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n30039), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n30038), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4786), .S(n66648));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1212 (.I0(\data_out_frame[13] [1]), .I1(n27006), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n67530));
    defparam i2_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4785), .S(n66647));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4784), .S(n66646));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n30037), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n30036), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n30035), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n30034), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n30033), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n30032), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4782), .S(n66645));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4781), .S(n66644));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4780), .S(n66643));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4779), .S(n66642));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n30031), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n30030), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n67355));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4778), .S(n66641));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n30029), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27058));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n30028), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4775), .S(n66580));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4774), .S(n66581));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4773), .S(n66582));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n30027), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n30026), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n30025), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4771), .S(n66583));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n30024), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4767), .S(n66584));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4766), .S(n66585));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4763), .S(n66586));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n30023), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4760), .S(n66588));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n30873), .D(n2_adj_4759), .S(n29288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4758), .S(n66589));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4755), .S(n66590));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n30022), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n30021), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n30020), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4754), .S(n66591));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1215 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66935));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1215.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4753), .S(n66592));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4752), .S(n66593));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n67379));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4751), .S(n66594));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4750), .S(n66595));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4749), .S(n66596));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4747), .S(n66578));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n30883), .D(n2_adj_4745), .S(n29278));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1217 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n67533));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1217.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n67590));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n30007));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n30003));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59502_2_lut (.I0(n79423), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n75273));
    defparam i59502_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter_c[3]), 
            .I1(n77507), .I2(n75296), .I3(byte_transmit_counter_c[4]), 
            .O(n79642));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i61611_3_lut (.I0(n79339), .I1(n79165), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n77467));
    defparam i61611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n79642_bdd_4_lut (.I0(n79642), .I1(n79213), .I2(n7_adj_4888), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[6]));
    defparam n79642_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n66957));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n30002));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n30001));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n30000));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29999));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29998));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29997));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29996));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29995));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29994));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29993));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16086_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[11]_c [1]), .O(n30300));
    defparam i16086_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29992));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1220 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n67004));   // verilog/coms.v(74[16:62])
    defparam i2_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1221 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[4] [3]), .I3(GND_net), .O(n27006));
    defparam i2_3_lut_adj_1221.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1193));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63691 (.I0(byte_transmit_counter_c[3]), 
            .I1(n77811), .I2(n75275), .I3(byte_transmit_counter_c[4]), 
            .O(n79630));
    defparam byte_transmit_counter_3__bdd_4_lut_63691.LUT_INIT = 16'he4aa;
    SB_LUT4 i16082_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[11]_c [0]), .O(n30296));
    defparam i16082_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29991));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29990));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29989));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29988));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29987));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode_c[4]), .C(clk16MHz), .D(n29985));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(\control_mode[5] ), .C(clk16MHz), .D(n29984));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(\control_mode[6] ), .C(clk16MHz), .D(n29983));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(\control_mode[7] ), .C(clk16MHz), .D(n29979));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(\current_limit[1] ), .C(clk16MHz), .D(n29976));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(\current_limit[2] ), .C(clk16MHz), .D(n29975));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(\current_limit[3] ), .C(clk16MHz), .D(n29974));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(\current_limit[4] ), .C(clk16MHz), .D(n29973));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(\current_limit[5] ), .C(clk16MHz), .D(n29972));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_3_lut_3_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(reset), .I3(GND_net), .O(n23094));   // verilog/coms.v(130[12] 305[6])
    defparam i2_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29944), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(\current_limit[0] ), .C(clk16MHz), .D(n29943));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29942));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29941));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29940), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29939), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29938), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29935), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4889), .S(n66597));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n26197));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n67102));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4890), .S(n66598));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4891), .S(n66599));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4892), .S(n66600));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4893), .S(n66601));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4894), .S(n66602));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4895), .S(n29271));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_out_frame[6] [6]), .I1(n67587), 
            .I2(GND_net), .I3(GND_net), .O(n27213));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4896), .S(n66603));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4897), .S(n66604));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4898), .S(n66605));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4899), .S(n66606));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4900), .S(n66607));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4901), .S(n66576));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4902), .S(n66608));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4903), .S(n29263));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4904), .S(n66609));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4905), .S(n29261));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4906), .S(n66610));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4907), .S(n66611));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4908), .S(n66612));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4909), .S(n66613));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4910), .S(n66614));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4911), .S(n66615));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4912), .S(n66616));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4913), .S(n29253));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1225 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n26724));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1226 (.I0(n66878), .I1(\data_out_frame[8] [3]), 
            .I2(n26064), .I3(GND_net), .O(n67358));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1226.LUT_INIT = 16'h9696;
    SB_LUT4 n79630_bdd_4_lut (.I0(n79630), .I1(n79207), .I2(n7_adj_4914), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[5]));
    defparam n79630_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1227 (.I0(n67016), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n14_adj_4915));
    defparam i2_3_lut_adj_1227.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1228 (.I0(\data_out_frame[4] [6]), .I1(n67400), 
            .I2(\data_out_frame[4] [7]), .I3(\data_out_frame[5] [5]), .O(n20_adj_4916));
    defparam i8_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i6_2_lut (.I0(\data_out_frame[4] [4]), .I1(n27006), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4917));
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1229 (.I0(\data_out_frame[7] [1]), .I1(n20_adj_4916), 
            .I2(n14_adj_4915), .I3(\data_out_frame[6] [4]), .O(n22_c));
    defparam i10_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1230 (.I0(n26064), .I1(n22_c), .I2(n18_adj_4917), 
            .I3(\data_out_frame[4] [5]), .O(n69691));
    defparam i11_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1231 (.I0(\data_out_frame[7] [4]), .I1(n69691), 
            .I2(n67590), .I3(n67391), .O(n16_adj_4918));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1232 (.I0(\data_out_frame[8] [3]), .I1(n67545), 
            .I2(\data_out_frame[8] [1]), .I3(n67004), .O(n17_adj_4919));   // verilog/coms.v(77[16:43])
    defparam i7_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.i_2043__i0  (.Q(\FRAME_MATCHER.i[0] ), .C(clk16MHz), 
            .D(n28325), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(n28676), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n66088));
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1233 (.I0(n17_adj_4919), .I1(\data_out_frame[7] [2]), 
            .I2(n16_adj_4918), .I3(\data_out_frame[7] [3]), .O(n69308));   // verilog/coms.v(77[16:43])
    defparam i9_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1234 (.I0(n67533), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[9] [7]), .I3(n67379), .O(n15_adj_4920));
    defparam i6_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.i_2043__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n28327), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n28329), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n28331), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n28333), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n28337), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n28339), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n28341), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n28343), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n28345), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n28347), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n28349), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n28351), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n28353), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n28355), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n28357), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n28359), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n28361), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n28363), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n28365), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n28367), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n28369), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n28371), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n28373), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n28375), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n28377), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n28379), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n28381), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n28383), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n28385), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i2  (.Q(\FRAME_MATCHER.i[2] ), .C(clk16MHz), 
            .D(n28387), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i1  (.Q(\FRAME_MATCHER.i[1] ), .C(clk16MHz), 
            .D(n28389), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4921), .S(n66617));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4922), .S(n29251));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4923), .S(n66618));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1235 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [7]), 
            .I2(n27058), .I3(\data_out_frame[11] [4]), .O(n12_adj_4924));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1236 (.I0(n15_adj_4920), .I1(n69308), .I2(n14_adj_4925), 
            .I3(\data_out_frame[7] [5]), .O(n68705));
    defparam i8_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4926), .S(n66619));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4927), .S(n66620));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4928), .S(n66621));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1237 (.I0(n68705), .I1(n12_adj_4924), .I2(n8_adj_4929), 
            .I3(n26813), .O(n66926));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1238 (.I0(\data_out_frame[12] [2]), .I1(n66926), 
            .I2(\data_out_frame[11] [5]), .I3(n67358), .O(n10_adj_4930));   // verilog/coms.v(88[17:63])
    defparam i4_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1239 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n26190));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n26752));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4931), .S(n66743));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4932), .S(n66742));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4933), .S(n66741));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i19831_3_lut (.I0(n38), .I1(n460), .I2(n486), .I3(GND_net), 
            .O(n40));
    defparam i19831_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i13_4_lut (.I0(n67530), .I1(n67347), .I2(n27292), .I3(\data_out_frame[14] [4]), 
            .O(n34_c));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_4936), 
            .I2(n41637), .I3(reset), .O(n66852));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i22183_3_lut (.I0(n34), .I1(deadband[17]), .I2(n462), .I3(GND_net), 
            .O(n36));
    defparam i22183_3_lut.LUT_INIT = 16'hb2b2;
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4938), .S(n66740));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4939), .S(n66739));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(\current_limit[8] ), .C(clk16MHz), .D(n30786));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i17_4_lut_adj_1241 (.I0(n1699), .I1(n34_c), .I2(n24_adj_4940), 
            .I3(n67188), .O(n38_adj_4941));
    defparam i17_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n67313), .I1(n61380), .I2(\data_out_frame[6] [0]), 
            .I3(n1720), .O(n36_adj_4942));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1242 (.I0(n28676), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n66092));
    defparam i1_4_lut_4_lut_4_lut_adj_1242.LUT_INIT = 16'hfe10;
    SB_LUT4 i19_4_lut_adj_1243 (.I0(\data_out_frame[14] [1]), .I1(n38_adj_4941), 
            .I2(n32), .I3(n61320), .O(n40_adj_4943));
    defparam i19_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i31192_2_lut_3_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(GND_net), .O(n45283));
    defparam i31192_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i14_4_lut_adj_1244 (.I0(n26943), .I1(n67545), .I2(\data_out_frame[14] [6]), 
            .I3(n67355), .O(n35_adj_4944));
    defparam i14_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 i60444_2_lut (.I0(displacement[11]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n75232));   // verilog/TinyFPGA_B.v(246[14:26])
    defparam i60444_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i39039_3_lut (.I0(encoder0_position_scaled[11]), .I1(encoder1_position_scaled[11]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n60595));   // verilog/TinyFPGA_B.v(246[14:26])
    defparam i39039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1245 (.I0(n60595), .I1(n53108), .I2(n75232), 
            .I3(control_mode[1]), .O(n42994));   // verilog/coms.v(130[12] 305[6])
    defparam i1_4_lut_adj_1245.LUT_INIT = 16'hfcdd;
    SB_DFF current_limit_i0_i9 (.Q(\current_limit[9] ), .C(clk16MHz), .D(n30785));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(\current_limit[10] ), .C(clk16MHz), 
           .D(n30781));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n37668));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(\current_limit[12] ), .C(clk16MHz), 
           .D(n30779));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n30778));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n30777));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n65900));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n30775));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n30774), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n30773), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n30772), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n30770), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n65896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n30768), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n30766), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30763));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n65892));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n65888));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i30186_3_lut (.I0(encoder0_position_scaled[12]), .I1(\motor_state_23__N_91[12] ), 
            .I2(n15), .I3(GND_net), .O(n10));
    defparam i30186_3_lut.LUT_INIT = 16'h3535;
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29731));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n29734));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[7] [1]), .O(n10_adj_4880));   // verilog/coms.v(88[17:70])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30740));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n65884));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29740));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n30737), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n30736), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19]_c [1]), .C(clk16MHz), 
           .D(n29743));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n30734));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n30733), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n30732), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19][2] ), .C(clk16MHz), 
           .D(n29746));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n30730), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30727));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19][3] ), .C(clk16MHz), 
           .D(n29749));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n30725), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19][4] ), .C(clk16MHz), 
           .D(n29752));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n30723), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n30722), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n30699), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n30681), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19][5] ), .C(clk16MHz), 
           .D(n29756));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n30679), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n30678));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n30666));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n30665), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n30664));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n30663));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n30662));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n30661));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n30660));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n30659));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n30658));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n30657));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n30656));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n30655));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n30654));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n30653));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n30652));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n30651));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n30650));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n30649));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n30648));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n30647));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n30646));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n30645));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n30644));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n30643));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n30642));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n30641));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1246 (.I0(\data_out_frame[16] [0]), .I1(n35_adj_4944), 
            .I2(n40_adj_4943), .I3(n36_adj_4942), .O(n67249));
    defparam i1_4_lut_adj_1246.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4777), .S(n66738));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n30640));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n30639));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n30638));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n30637));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n30636));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n30635));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n30634));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n30633), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n30632));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n30631), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n30630), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n30249));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19][6] ), .C(clk16MHz), 
           .D(n29759));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n30252));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n30626), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n30255));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n30624), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19][7] ), .C(clk16MHz), 
           .D(n29763));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n30258));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n30261));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n30264));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n30619));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30616));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4762), .S(n66737));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20][0] ), .C(clk16MHz), 
           .D(n29766));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20][1] ), .C(clk16MHz), 
           .D(n29769));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20][2] ), .C(clk16MHz), 
           .D(n29772));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n29776));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n29779));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20][4] ), .C(clk16MHz), 
           .D(n29782));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n65834));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n29788));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n65838));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29794));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29797));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n30267));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n30603));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29800));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n29803));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
           .D(n30270));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
           .D(n30273));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1247 (.I0(n62080), .I1(n67271), .I2(GND_net), 
            .I3(GND_net), .O(n62277));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
           .D(n66088));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
           .D(n30280));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n66092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
           .D(n30286));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n30290));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30593));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n29806));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n30589));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n30588));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29809));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
           .D(n30293));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n30585));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29812));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29815));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11]_c [0]), .C(clk16MHz), 
           .D(n30296));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11]_c [1]), .C(clk16MHz), 
           .D(n30300));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11]_c [2]), .C(clk16MHz), 
           .D(n66022));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11]_c [3]), .C(clk16MHz), 
           .D(n30306));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11]_c [4]), .C(clk16MHz), 
           .D(n30310));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11]_c [5]), .C(clk16MHz), 
           .D(n66068));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11]_c [6]), .C(clk16MHz), 
           .D(n30316));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n30320));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n30323));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29818));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n30326));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12][2] ), .C(clk16MHz), 
           .D(n66112));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12][3] ), .C(clk16MHz), 
           .D(n66142));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12][4] ), .C(clk16MHz), 
           .D(n66144));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12][5] ), .C(clk16MHz), 
           .D(n30339));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12][6] ), .C(clk16MHz), 
           .D(n30342));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n30346));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13][0] ), .C(clk16MHz), 
           .D(n30349));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n30352));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13][2] ), .C(clk16MHz), 
           .D(n30355));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n30359));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13][4] ), .C(clk16MHz), 
           .D(n30362));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13][5] ), .C(clk16MHz), 
           .D(n30365));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13][6] ), .C(clk16MHz), 
           .D(n30368));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13][7] ), .C(clk16MHz), 
           .D(n30372));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n30375));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4947), .S(n66736));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4948), .S(n66735));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i114 (.Q(\data_in_frame[14]_c [1]), .C(clk16MHz), 
           .D(n30378));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i115 (.Q(\data_in_frame[14][2] ), .C(clk16MHz), 
           .D(n30382));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1248 (.I0(n62342), .I1(n62473), .I2(\data_in_frame[16] [3]), 
            .I3(n26551), .O(n61016));
    defparam i1_2_lut_3_lut_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i116 (.Q(\data_in_frame[14]_c [3]), .C(clk16MHz), 
           .D(n30385));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14][4] ), .C(clk16MHz), 
           .D(n30388));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i118 (.Q(\data_in_frame[14][5] ), .C(clk16MHz), 
           .D(n30392));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i119 (.Q(\data_in_frame[14][6] ), .C(clk16MHz), 
           .D(n30395));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1249 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25859), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n71998));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1249.LUT_INIT = 16'hfff4;
    SB_DFF data_in_frame_0___i120 (.Q(\data_in_frame[14][7] ), .C(clk16MHz), 
           .D(n30398));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n30402));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n30405));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n30408));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n30412));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n15_adj_4949));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15][5] ), .C(clk16MHz), 
           .D(n30418));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n30422));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n30425));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16][0] ), .C(clk16MHz), 
           .D(n65878));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n30432));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n65874));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n65870));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n65842));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16]_c [5]), .C(clk16MHz), 
           .D(n30445));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16]_c [6]), .C(clk16MHz), 
           .D(n30448));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16][7] ), .C(clk16MHz), 
           .D(n65866));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n65960));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n30458));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n65998));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n65994));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n65990));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n30517));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4950), .S(n66734));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29821));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n29824));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1250 (.I0(n26345), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[13][4] ), .I3(n67043), .O(n61494));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29827));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n29830));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29833));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29836));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n29839));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26053));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29842));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29845));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n66130));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
           .D(n66084));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n66132));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n65966));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n30469));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29863));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n65964));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n65962));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n29872));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n29876));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n29879));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
           .D(n66128));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1252 (.I0(\data_in_frame[10] [4]), .I1(n67111), 
            .I2(\data_in_frame[12][5] ), .I3(n26875), .O(n26418));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
           .D(n29885));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i10 (.Q(\data_in_frame[1][1] ), .C(clk16MHz), 
           .D(n29888));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1253 (.I0(n26687), .I1(n26848), .I2(\data_in_frame[9] [2]), 
            .I3(\data_in_frame[14]_c [1]), .O(n9_adj_4951));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i11 (.Q(\data_in_frame[1][2] ), .C(clk16MHz), 
           .D(n29891));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i12 (.Q(\data_in_frame[1][3] ), .C(clk16MHz), 
           .D(n29894));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n29897));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1][5] ), .C(clk16MHz), 
           .D(n29900));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1][6] ), .C(clk16MHz), 
           .D(n29903));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1][7] ), .C(clk16MHz), 
           .D(n29907));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
           .D(n29911));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
           .D(n29916));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1254 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n67548));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1254.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
           .D(n29919));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1255 (.I0(\data_out_frame[12] [3]), .I1(n67548), 
            .I2(n67013), .I3(\data_out_frame[10] [1]), .O(n10_adj_4952));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
           .D(n29922));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
           .D(n29925));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1256 (.I0(\data_out_frame[12] [4]), .I1(n66967), 
            .I2(n35_adj_4953), .I3(GND_net), .O(n1655));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1256.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4954), .S(n66733));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1257 (.I0(n28658), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n65834));
    defparam i1_4_lut_4_lut_4_lut_adj_1257.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4955), .S(n66732));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4956), .S(n66731));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4957), .S(n66730));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4958), .S(n66729));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1258 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[10] [1]), .O(n68795));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1259 (.I0(n68795), .I1(\data_out_frame[7] [6]), 
            .I2(n67599), .I3(\data_out_frame[14] [3]), .O(n67313));
    defparam i3_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
           .D(n29928));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
           .D(n29931));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4959), .S(n66728));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1260 (.I0(n28658), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n65838));
    defparam i1_4_lut_4_lut_4_lut_adj_1260.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4960), .S(n66727));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1261 (.I0(n61517), .I1(n67313), .I2(\data_out_frame[7] [7]), 
            .I3(\data_out_frame[12] [2]), .O(n62261));
    defparam i3_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1262 (.I0(n26592), .I1(n27292), .I2(n62261), 
            .I3(\data_out_frame[16] [6]), .O(n10_adj_4961));
    defparam i4_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n28131), 
            .D(n4932[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n28131), 
            .D(n4932[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n28131), 
            .D(n4932[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n28131), 
            .D(n4932[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n28131), 
            .D(n4932[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n28131), 
            .D(n4932[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n28131), 
            .D(n4932[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n28131), 
            .D(n4932[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n28131), 
            .D(n4932[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n28131), 
            .D(n4932[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n28131), 
            .D(n4932[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n28131), 
            .D(n4932[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n28131), 
            .D(n4932[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n28131), 
            .D(n4932[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n28131), 
            .D(n4932[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n28131), 
            .D(n4932[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n28131), 
            .D(n4932[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n28131), 
            .D(n4932[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n28131), 
            .D(n4932[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n28131), 
            .D(n4932[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n28131), 
            .D(n4932[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n28131), 
            .D(n4932[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n28131), 
            .D(n4932[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n79682), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n27429), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2048), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2049), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20639), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n65734), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2060), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n27432), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4962), .S(n66726));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1263 (.I0(\data_out_frame[16] [4]), .I1(n10_adj_4961), 
            .I2(n26311), .I3(GND_net), .O(n69868));
    defparam i5_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4963), .S(n66725));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4964), .S(n66724));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4965), .S(n66723));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26475));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4966), .S(n29387));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4967), .S(n66722));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4968), .S(n66721));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4969), .S(n66720));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4970), .S(n66719));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4971), .S(n66718));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4972), .S(n66717));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4973), .S(n66716));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4974), .S(n66715));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4975), .S(n66714));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4976), .S(n66713));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4977), .S(n66712));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1265 (.I0(\data_out_frame[18] [7]), .I1(n26592), 
            .I2(n69868), .I3(\data_out_frame[19] [1]), .O(n67572));
    defparam i3_4_lut_adj_1265.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67593));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n67551));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1268 (.I0(\data_in_frame[13][5] ), .I1(n26345), 
            .I2(n26364), .I3(\data_in_frame[17] [3]), .O(n71760));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i59537_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75099));   // verilog/coms.v(158[12:15])
    defparam i59537_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i59876_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75100));   // verilog/coms.v(158[12:15])
    defparam i59876_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1269 (.I0(\data_in_frame[13][5] ), .I1(n26345), 
            .I2(n26364), .I3(\data_in_frame[15] [6]), .O(n67581));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4849));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66922));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1271 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n67016));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1271.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1272 (.I0(\data_in_frame[2] [3]), .I1(n67129), 
            .I2(n67441), .I3(n26721), .O(n67456));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4848));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1273 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[8] [0]), .I3(\data_out_frame[8] [2]), .O(n67391));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4978), .S(n66711));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4979), .S(n29374));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59584_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75103));   // verilog/coms.v(158[12:15])
    defparam i59584_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4980), .S(n66710));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1274 (.I0(\data_out_frame[5] [4]), .I1(n67391), 
            .I2(n67016), .I3(n66922), .O(n35_adj_4953));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(n35_adj_4953), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4981));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(n67397), .I1(n67013), .I2(n67551), 
            .I3(n6_adj_4981), .O(n67094));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4982), .S(n66622));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4983), .S(n66623));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(\current_limit[6] ), .C(clk16MHz), .D(n29755));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n31022), .D(n2_adj_4984), .S(n29244));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n31023), .D(n2_adj_4985), .S(n29243));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4986), .S(n66624));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4987), .S(n66625));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4988), .S(n66626));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1277 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_767), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[3] [0]), .O(n26986));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4989), .S(n66627));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4990), .S(n66628));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4991), .S(n66629));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4992), .S(n29236));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n31031), .D(n2_adj_4993), .S(n29235));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4994), .S(n66587));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4995), .S(n66630));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n31034), .D(n2_adj_4996), .S(n29232));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59670_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75124));   // verilog/coms.v(158[12:15])
    defparam i59670_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4997), .S(n66709));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i60416_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75127));   // verilog/coms.v(158[12:15])
    defparam i60416_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4847));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59652_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75131));   // verilog/coms.v(158[12:15])
    defparam i59652_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1278 (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i[0] ), 
            .I2(n44662), .I3(n82), .O(n28703));
    defparam i1_2_lut_3_lut_4_lut_adj_1278.LUT_INIT = 16'h4000;
    SB_LUT4 select_787_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4846));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4845));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1279 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[6] [5]), .I3(n67456), .O(Kp_23__N_993));
    defparam i1_2_lut_3_lut_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4844));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1280 (.I0(n28672), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[12][2] ), .O(n66112));
    defparam i1_4_lut_4_lut_4_lut_adj_1280.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1281 (.I0(n67572), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[16] [1]), .I3(n26475), .O(n67229));
    defparam i3_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4843));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4998), .S(n66708));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\data_out_frame[17] [0]), .I1(n27159), 
            .I2(GND_net), .I3(GND_net), .O(n27298));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4999), .S(n66707));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n31038), .D(n2_adj_5000), .S(n29369));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n31039), .D(n2_adj_5001), .S(n29231));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1283 (.I0(n26311), .I1(n67249), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5002));
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5003), .S(n66631));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5004), .S(n66632));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5005), .S(n66633));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5006), .S(n66634));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5007), .S(n66635));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5008), .S(n66636));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n31046), .D(n2_adj_5009), .S(n29224));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5010), .S(n66579));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5011), .S(n66637));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5012), .S(n66638));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5013), .S(n66639));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5014), .S(n66640));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5015), .S(n66761));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4864), .S(n66762));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4772), .S(n66763));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4769), .S(n66764));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4768), .S(n66760));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4765), .S(n66765));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5016), .S(n66766));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1284 (.I0(n62281), .I1(n69868), .I2(n67207), 
            .I3(n6_adj_5002), .O(n61795));
    defparam i4_4_lut_adj_1284.LUT_INIT = 16'h9669;
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2874), .D(n5_c), 
            .S(n29211));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4757), .S(n66767));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_4748), .S(n66706));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2874), .D(n27318), 
            .S(n29201));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2874), .D(n1_c), .S(n29195));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4744), .S(n66768));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4743), .S(n66769));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4740), .S(n66770));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4738), .S(n66758));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4737), .S(n66759));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5017), .S(n66771));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_4736), .S(n66772));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2874), .D(n3), .S(n66773));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n2874), .D(n1_adj_5018), .S(n66751));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5019), .S(n66752));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n31088), .D(n2), .S(n29367));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(\current_limit[7] ), .C(clk16MHz), .D(n29727));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n31093), .D(n2_adj_5020), .S(n29366));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4842));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5021), .S(n66753));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1285 (.I0(\data_out_frame[23] [5]), .I1(n61447), 
            .I2(n61577), .I3(\data_out_frame[25] [0]), .O(n67061));
    defparam i1_2_lut_3_lut_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4841));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1286 (.I0(\data_out_frame[23] [5]), .I1(n61447), 
            .I2(n61577), .I3(n62464), .O(n67126));
    defparam i1_2_lut_3_lut_4_lut_adj_1286.LUT_INIT = 16'h9669;
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), 
            .C(clk16MHz), .E(n2874), .D(n1_adj_5022), .S(n66754));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5023), .S(n66749));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), 
            .C(clk16MHz), .E(n2874), .D(n1_adj_5024), .S(n66755));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n2874), .D(n1_adj_5025), .S(n66756));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5026), .S(n66705));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5027), .S(n66704));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n2874), .D(n1_adj_5028), .S(n66750));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5029), .S(n66702));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4840));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5030), .S(n66701));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1287 (.I0(control_mode[0]), .I1(n53108), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_6));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1287.LUT_INIT = 16'hefef;
    SB_LUT4 select_787_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4839));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1288 (.I0(n27298), .I1(\data_out_frame[19] [0]), 
            .I2(n67229), .I3(n6_adj_5032), .O(n27164));
    defparam i4_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1289 (.I0(\data_out_frame[21] [3]), .I1(n67216), 
            .I2(n61384), .I3(\data_out_frame[17] [1]), .O(n61577));
    defparam i3_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 i16420_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n30634));   // verilog/coms.v(130[12] 305[6])
    defparam i16420_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4838));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(\data_out_frame[21] [2]), .I1(n27164), 
            .I2(GND_net), .I3(GND_net), .O(n61294));
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1291 (.I0(n67503), .I1(\data_out_frame[19] [3]), 
            .I2(n61503), .I3(n61824), .O(n67286));
    defparam i3_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i16450_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n30664));   // verilog/coms.v(130[12] 305[6])
    defparam i16450_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4837));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15737_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29951));   // verilog/coms.v(130[12] 305[6])
    defparam i15737_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4836));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16449_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n30663));   // verilog/coms.v(130[12] 305[6])
    defparam i16449_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4835));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16448_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n30662));   // verilog/coms.v(130[12] 305[6])
    defparam i16448_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4834));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16447_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n30661));   // verilog/coms.v(130[12] 305[6])
    defparam i16447_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4833));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16446_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n30660));   // verilog/coms.v(130[12] 305[6])
    defparam i16446_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4832));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59629_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75132));   // verilog/coms.v(158[12:15])
    defparam i59629_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(\data_out_frame[21] [4]), .I1(\data_out_frame[19] [3]), 
            .I2(n67139), .I3(n6_adj_5033), .O(n61447));   // verilog/coms.v(79[16:43])
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n67435));
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i16445_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n30659));   // verilog/coms.v(130[12] 305[6])
    defparam i16445_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_208_i3_4_lut (.I0(n62268), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5034), .I3(n67286), .O(n3_adj_5015));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i16444_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n30658));   // verilog/coms.v(130[12] 305[6])
    defparam i16444_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_207_i2_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5014));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_207_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59656_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75133));   // verilog/coms.v(158[12:15])
    defparam i59656_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5013));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16443_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n30657));   // verilog/coms.v(130[12] 305[6])
    defparam i16443_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5012));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59678_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75144));   // verilog/coms.v(158[12:15])
    defparam i59678_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16441_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n30655));   // verilog/coms.v(130[12] 305[6])
    defparam i16441_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i59681_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75145));   // verilog/coms.v(158[12:15])
    defparam i59681_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i28798_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_7), .I3(n15_adj_6), .O(\motor_state_23__N_91[8] ));
    defparam i28798_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_787_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5011));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16440_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n30654));   // verilog/coms.v(130[12] 305[6])
    defparam i16440_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1294 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [3]), 
            .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5010));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1294.LUT_INIT = 16'ha088;
    SB_LUT4 i16439_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n30653));   // verilog/coms.v(130[12] 305[6])
    defparam i16439_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16438_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n30652));   // verilog/coms.v(130[12] 305[6])
    defparam i16438_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1295 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [2]), 
            .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5009));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1295.LUT_INIT = 16'ha088;
    SB_LUT4 i16437_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n30651));   // verilog/coms.v(130[12] 305[6])
    defparam i16437_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5008));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16436_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n30650));   // verilog/coms.v(130[12] 305[6])
    defparam i16436_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5007));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16435_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n30649));   // verilog/coms.v(130[12] 305[6])
    defparam i16435_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5006));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16434_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n30648));   // verilog/coms.v(130[12] 305[6])
    defparam i16434_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i59711_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75167));   // verilog/coms.v(158[12:15])
    defparam i59711_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16433_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n30647));   // verilog/coms.v(130[12] 305[6])
    defparam i16433_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5005));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16432_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n30646));   // verilog/coms.v(130[12] 305[6])
    defparam i16432_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4831));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5004));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16431_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n30645));   // verilog/coms.v(130[12] 305[6])
    defparam i16431_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5030));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16430_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n30644));   // verilog/coms.v(130[12] 305[6])
    defparam i16430_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16429_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n30643));   // verilog/coms.v(130[12] 305[6])
    defparam i16429_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16428_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n30642));   // verilog/coms.v(130[12] 305[6])
    defparam i16428_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16427_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n30641));   // verilog/coms.v(130[12] 305[6])
    defparam i16427_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_1194_9_lut (.I0(n66748), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n59006), .O(n66751)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16426_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n30640));   // verilog/coms.v(130[12] 305[6])
    defparam i16426_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16425_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n30639));   // verilog/coms.v(130[12] 305[6])
    defparam i16425_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5003));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16424_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n30638));   // verilog/coms.v(130[12] 305[6])
    defparam i16424_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4830));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1194_8_lut (.I0(n66748), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n59005), .O(n66750)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16423_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n30637));   // verilog/coms.v(130[12] 305[6])
    defparam i16423_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_1194_8 (.CI(n59005), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n59006));
    SB_LUT4 add_1194_7_lut (.I0(n66748), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n59004), .O(n66756)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16422_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n30636));   // verilog/coms.v(130[12] 305[6])
    defparam i16422_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16421_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n30635));   // verilog/coms.v(130[12] 305[6])
    defparam i16421_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_1194_7 (.CI(n59004), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n59005));
    SB_LUT4 add_1194_6_lut (.I0(n66748), .I1(byte_transmit_counter_c[4]), 
            .I2(GND_net), .I3(n59003), .O(n66755)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16442_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n30656));   // verilog/coms.v(130[12] 305[6])
    defparam i16442_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_1194_6 (.CI(n59003), .I0(byte_transmit_counter_c[4]), .I1(GND_net), 
            .CO(n59004));
    SB_LUT4 add_1194_5_lut (.I0(n66748), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(n59002), .O(n66754)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_5 (.CI(n59002), .I0(byte_transmit_counter_c[3]), .I1(GND_net), 
            .CO(n59003));
    SB_LUT4 add_1194_4_lut (.I0(n66748), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n59001), .O(n66753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_4 (.CI(n59001), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n59002));
    SB_LUT4 add_1194_3_lut (.I0(n66748), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n59000), .O(n66752)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_787_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5029));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY add_1194_3 (.CI(n59000), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n59001));
    SB_LUT4 add_1194_2_lut (.I0(n66748), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n66749)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[20] [5]), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[18] [4]), .I3(\data_in_frame[22] [6]), .O(n6_adj_5036));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1296 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [3]), 
            .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5001));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1296.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(n62342), .I1(\data_in_frame[14][2] ), 
            .I2(n62356), .I3(GND_net), .O(n25590));
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[3] [5]), .O(n71704));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_1194_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3416), 
            .CO(n59000));
    SB_LUT4 i1_4_lut_adj_1298 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[10] [3]), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4829));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1298.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1299 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [4]), .O(n27052));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[0] [3]), .I1(n67067), .I2(\data_in_frame[2] [3]), 
            .I3(n67129), .O(Kp_23__N_799));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1300 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n41637), .O(n28658));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1300.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1301 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n66860), .O(n66867));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1301.LUT_INIT = 16'hffef;
    SB_LUT4 select_787_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5027));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1302 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1][1] ), 
            .I2(n67338), .I3(\data_in_frame[1] [4]), .O(Kp_23__N_767));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5026));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4828));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1303 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n66868), .O(n66869));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1303.LUT_INIT = 16'hffbf;
    SB_LUT4 select_787_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5000));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1304 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n66860), .O(n66862));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1304.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_4_lut_adj_1305 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[7] [4]), 
            .I2(encoder0_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5020));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1305.LUT_INIT = 16'ha088;
    SB_LUT4 i16132_3_lut_4_lut (.I0(n28672), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n30346));
    defparam i16132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1306 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(n67067), .I3(n26752), .O(n26721));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4999));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4998));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n66761));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_adj_1307 (.I0(n27258), .I1(\data_out_frame[16] [6]), 
            .I2(n61795), .I3(GND_net), .O(n6_adj_5032));
    defparam i1_2_lut_3_lut_adj_1307.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1308 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n66762));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1308.LUT_INIT = 16'h5100;
    SB_LUT4 i2_3_lut_4_lut_adj_1309 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[14] [6]), .I3(n67094), .O(n27159));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4827));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1310 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [2]), 
            .O(n66763));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1310.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1311 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n66764));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1311.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_adj_1312 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[10] [0]), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4826));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1312.LUT_INIT = 16'ha088;
    SB_LUT4 i2_3_lut_4_lut_adj_1313 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[12] [1]), .I3(n36341), .O(n67474));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1314 (.I0(n26687), .I1(n26848), .I2(n67412), 
            .I3(GND_net), .O(n67554));
    defparam i1_2_lut_3_lut_adj_1314.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4825));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1315 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n66760));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1315.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4824));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1316 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n66765));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1316.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4997));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1317 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n66766));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1317.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4823));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1318 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[7] [7]), 
            .I2(n67105), .I3(\data_in_frame[1][5] ), .O(n67462));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1319 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [4]), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4822));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1319.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1320 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n66767));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1320.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_adj_1321 (.I0(n27048), .I1(n26585), .I2(n10_adj_5037), 
            .I3(\data_in_frame[7] [4]), .O(n24270));
    defparam i1_2_lut_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i16128_3_lut_4_lut (.I0(n28672), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[12][6] ), .O(n30342));
    defparam i16128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4821));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1322 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [2]), 
            .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4996));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1322.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4995));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(\data_in_frame[11]_c [6]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n67560));
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4820));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1324 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[10] [3]), .O(n67397));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4994));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1325 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n26060));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1326 (.I0(n28672), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[12][4] ), .O(n66144));
    defparam i1_4_lut_4_lut_4_lut_adj_1326.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1327 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n66768));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1327.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_adj_1328 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [7]), 
            .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4993));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1328.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1329 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n66769));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1329.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4992));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1330 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [2]), 
            .O(n66770));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1330.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4991));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1331 (.I0(\data_in_frame[11]_c [3]), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[9] [2]), .I3(\data_in_frame[8] [7]), .O(n67406));
    defparam i2_3_lut_4_lut_adj_1331.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4990));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1332 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n66758));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1332.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4989));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1333 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n66759));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1333.LUT_INIT = 16'h5100;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63681 (.I0(byte_transmit_counter_c[3]), 
            .I1(n77467), .I2(n75273), .I3(byte_transmit_counter_c[4]), 
            .O(n79528));
    defparam byte_transmit_counter_3__bdd_4_lut_63681.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4819));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4988));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4818));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4817));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1334 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n66771));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1334.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4987));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1335 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n66772));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1335.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_adj_1336 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [6]), 
            .I2(encoder0_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4816));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1336.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4986));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1337 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n66773));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1337.LUT_INIT = 16'h5100;
    SB_LUT4 i59722_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75168));   // verilog/coms.v(158[12:15])
    defparam i59722_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4985));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4984));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1338 (.I0(n26818), .I1(n26317), .I2(n27225), 
            .I3(\data_in_frame[8] [2]), .O(n67111));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i59724_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75171));   // verilog/coms.v(158[12:15])
    defparam i59724_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n67361));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4983));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[7] [5]), .I3(n10_adj_4952), .O(n66967));   // verilog/coms.v(78[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1340 (.I0(\data_in_frame[15] [2]), .I1(n26246), 
            .I2(n26331), .I3(\data_in_frame[10] [6]), .O(n67584));
    defparam i1_2_lut_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1341 (.I0(\data_in_frame[11]_c [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n26776));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1341.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4982));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59726_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75181));   // verilog/coms.v(158[12:15])
    defparam i59726_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n79528_bdd_4_lut (.I0(n79528), .I1(n79159), .I2(n7_adj_5038), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[1]));
    defparam n79528_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [5]), .I3(n67167), .O(n24_adj_4940));   // verilog/coms.v(79[16:43])
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4980));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1342 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [5]), .I3(n62080), .O(n67332));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1343 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [5]), .I3(n67425), .O(n6_adj_4856));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1344 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[8] [5]), .I3(n66957), .O(n26813));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1345 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n26064));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1346 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[6] [4]), 
            .I2(encoder0_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4979));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1346.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1347 (.I0(n28692), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n66130));
    defparam i1_4_lut_4_lut_4_lut_adj_1347.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4978));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n67545));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1349 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n66929));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1349.LUT_INIT = 16'h9696;
    SB_LUT4 LessThan_26_i38_3_lut_3_lut (.I0(deadband[19]), .I1(n460), .I2(n461), 
            .I3(GND_net), .O(n38_adj_8));
    defparam LessThan_26_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_3_lut_adj_1350 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n6_adj_5040));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1350.LUT_INIT = 16'h9696;
    SB_LUT4 i59959_3_lut_4_lut (.I0(deadband[19]), .I1(n460), .I2(n461), 
            .I3(deadband[18]), .O(n75815));
    defparam i59959_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(n26480), .I3(GND_net), .O(n6));
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1352 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11]_c [2]), 
            .I2(n67468), .I3(n26687), .O(n26959));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n67468));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1354 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(n26813), .I3(\data_out_frame[9] [1]), .O(n14_adj_4925));
    defparam i5_3_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1355 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(n26053), .I3(n67004), .O(n1168));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n67536));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 i60411_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75189));   // verilog/coms.v(158[12:15])
    defparam i60411_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(n69576), .I1(\data_in_frame[15][5] ), 
            .I2(n24167), .I3(GND_net), .O(n67284));
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'h6969;
    SB_LUT4 i59729_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n75190));   // verilog/coms.v(158[12:15])
    defparam i59729_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4977));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14438_1_lut (.I0(n3476), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n28651));   // verilog/coms.v(148[4] 304[11])
    defparam i14438_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1358 (.I0(n28692), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n66128));
    defparam i1_4_lut_4_lut_4_lut_adj_1358.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4808));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_301_i7_2_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4936));   // verilog/coms.v(157[7:23])
    defparam equal_301_i7_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 select_787_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4976));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4975));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1359 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [7]), 
            .I2(\control_mode[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4974));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1359.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(n26818), .I1(\data_in_frame[10] [5]), 
            .I2(n26331), .I3(GND_net), .O(n67385));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1361 (.I0(n69576), .I1(n67539), .I2(\data_in_frame[17] [7]), 
            .I3(\data_in_frame[17] [6]), .O(n67149));
    defparam i2_3_lut_4_lut_adj_1361.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1362 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [6]), 
            .I2(\control_mode[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4973));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1362.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4972));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1363 (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[13][5] ), 
            .I2(n67329), .I3(\data_in_frame[15] [6]), .O(n66945));
    defparam i1_2_lut_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4971));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(\data_in_frame[20] [5]), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[18] [4]), .I3(GND_net), .O(n67262));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4970));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_3_lut_4_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(n66961), .I3(n61378), .O(n32));   // verilog/coms.v(74[16:27])
    defparam i11_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4969));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4968));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1365 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [0]), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4967));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1365.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [4]), .I2(\data_out_frame[7] [4]), .I3(byte_transmit_counter[1]), 
            .O(n79522));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4966));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4965));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4964));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4963));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[13][0] ), 
            .I2(\data_in_frame[13][2] ), .I3(GND_net), .O(n6_adj_5042));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 n79522_bdd_4_lut (.I0(n79522), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(byte_transmit_counter[1]), 
            .O(n72450));
    defparam n79522_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1366 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [3]), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4962));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1366.LUT_INIT = 16'ha088;
    SB_LUT4 i61605_3_lut (.I0(n79417), .I1(n79243), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n77461));
    defparam i61605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61606_4_lut (.I0(n77461), .I1(n79411), .I2(byte_transmit_counter_c[3]), 
            .I3(byte_transmit_counter[2]), .O(n77462));
    defparam i61606_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i56436_3_lut (.I0(n79147), .I1(n77462), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(tx_data[4]));
    defparam i56436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n1), .I2(n5), .I3(byte_transmit_counter[2]), .O(n79516));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1367 (.I0(\data_out_frame[11] [5]), .I1(n61164), 
            .I2(n26783), .I3(GND_net), .O(n67259));
    defparam i1_2_lut_3_lut_adj_1367.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1368 (.I0(\data_out_frame[11] [5]), .I1(n61164), 
            .I2(n27184), .I3(n27089), .O(n61378));
    defparam i2_3_lut_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i6772_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1951), 
            .I2(n68793), .I3(n4452), .O(n20634));   // verilog/coms.v(148[4] 304[11])
    defparam i6772_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1369 (.I0(n20634), .I1(n1951), .I2(n23017), .I3(n71998), 
            .O(n27432));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1369.LUT_INIT = 16'hbbba;
    SB_LUT4 i460_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2060));   // verilog/coms.v(148[4] 304[11])
    defparam i460_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_787_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4799));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1370 (.I0(n62383), .I1(n69522), .I2(\data_in_frame[20] [6]), 
            .I3(\data_in_frame[21] [0]), .O(n71754));
    defparam i1_4_lut_adj_1370.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1371 (.I0(n25590), .I1(n67341), .I2(n67497), 
            .I3(n71754), .O(n61755));
    defparam i1_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1372 (.I0(n61016), .I1(\data_in_frame[20] [6]), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n67373));
    defparam i2_3_lut_adj_1372.LUT_INIT = 16'h9696;
    SB_LUT4 i56159_4_lut (.I0(n1951), .I1(n1954), .I2(n3303), .I3(n1957), 
            .O(n72001));   // verilog/coms.v(139[4] 141[7])
    defparam i56159_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n71620));
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1374 (.I0(n69485), .I1(n69866), .I2(n27045), 
            .I3(n71620), .O(n67341));
    defparam i1_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1375 (.I0(\data_in_frame[18] [7]), .I1(n62404), 
            .I2(\data_in_frame[20] [7]), .I3(\data_in_frame[18] [4]), .O(n69568));
    defparam i3_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1376 (.I0(\data_in_frame[11]_c [6]), .I1(n67301), 
            .I2(n67170), .I3(n71938), .O(n71942));
    defparam i1_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1377 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[20][0] ), .I3(GND_net), .O(n71836));
    defparam i1_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1378 (.I0(n71836), .I1(n66932), .I2(\data_in_frame[19][7] ), 
            .I3(\data_in_frame[18] [6]), .O(n71840));
    defparam i1_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1379 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1954), 
            .I2(n72001), .I3(n68593), .O(n65734));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1379.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1_4_lut_adj_1380 (.I0(n62406), .I1(n67539), .I2(n67262), 
            .I3(n71840), .O(n71846));
    defparam i1_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1381 (.I0(n67316), .I1(n67283), .I2(n62365), 
            .I3(n71846), .O(n71852));
    defparam i1_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1382 (.I0(n61366), .I1(n67373), .I2(n67382), 
            .I3(n71852), .O(n71858));
    defparam i1_4_lut_adj_1382.LUT_INIT = 16'h9669;
    SB_LUT4 i6777_4_lut (.I0(n1955), .I1(\FRAME_MATCHER.state[3] ), .I2(n1957), 
            .I3(n25859), .O(n20639));   // verilog/coms.v(148[4] 304[11])
    defparam i6777_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_adj_1383 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[21] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66893));
    defparam i1_2_lut_adj_1383.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1384 (.I0(n61424), .I1(n67298), .I2(n71858), 
            .I3(n67152), .O(n71864));
    defparam i1_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1385 (.I0(n67191), .I1(n67064), .I2(n66893), 
            .I3(\data_in_frame[21] [7]), .O(n69350));
    defparam i1_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1386 (.I0(n69350), .I1(n71864), .I2(n24227), 
            .I3(n69224), .O(n66970));
    defparam i1_4_lut_adj_1386.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1387 (.I0(\data_in_frame[16]_c [6]), .I1(n67194), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5045));
    defparam i1_2_lut_adj_1387.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1388 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[19]_c [1]), 
            .I2(n69042), .I3(n6_adj_5045), .O(n62365));
    defparam i4_4_lut_adj_1388.LUT_INIT = 16'h9669;
    SB_LUT4 i449_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2049));   // verilog/coms.v(148[4] 304[11])
    defparam i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1389 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[21] [4]), 
            .I2(n62365), .I3(GND_net), .O(n67191));
    defparam i2_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 i448_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2048));   // verilog/coms.v(148[4] 304[11])
    defparam i448_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1390 (.I0(\data_in_frame[16]_c [5]), .I1(n6_adj_9), 
            .I2(n66889), .I3(n67310), .O(n67194));
    defparam i1_4_lut_adj_1390.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1391 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16][0] ), 
            .I2(n67246), .I3(n6_adj_5047), .O(n69065));
    defparam i4_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1392 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16));
    defparam i2_2_lut_adj_1392.LUT_INIT = 16'h6666;
    SB_LUT4 n79516_bdd_4_lut (.I0(n79516), .I1(n75196), .I2(n1_adj_4886), 
            .I3(byte_transmit_counter[2]), .O(n72454));
    defparam n79516_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i30728_4_lut (.I0(n5_adj_5049), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i30728_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(\FRAME_MATCHER.i [4]), .I1(n25879), .I2(GND_net), 
            .I3(GND_net), .O(n25749));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'heeee;
    SB_LUT4 i30732_4_lut (.I0(n8_adj_5), .I1(\FRAME_MATCHER.i [31]), .I2(n25749), 
            .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i30732_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_2_lut_adj_1394 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n23017));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1394.LUT_INIT = 16'h4444;
    SB_LUT4 i3_2_lut (.I0(n25859), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n27994));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1395 (.I0(n69522), .I1(n69485), .I2(n67232), 
            .I3(GND_net), .O(n69866));
    defparam i1_3_lut_adj_1395.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1396 (.I0(n4452), .I1(n27994), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n23017), .O(n69098));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1396.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_4_lut_adj_1397 (.I0(n67364), .I1(n6_adj_9), .I2(\data_in_frame[12][6] ), 
            .I3(\data_in_frame[15] [7]), .O(n71812));
    defparam i1_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1398 (.I0(n25868), .I1(n1957), .I2(n1955), .I3(n69098), 
            .O(n27429));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1398.LUT_INIT = 16'hbaaa;
    SB_LUT4 i1_4_lut_adj_1399 (.I0(n67581), .I1(n26872), .I2(n66985), 
            .I3(n71812), .O(n71818));
    defparam i1_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1400 (.I0(n62266), .I1(n62313), .I2(n66889), 
            .I3(n71818), .O(n71824));
    defparam i1_4_lut_adj_1400.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1401 (.I0(n67284), .I1(n67500), .I2(n69062), 
            .I3(n71824), .O(n69224));
    defparam i1_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27045));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1403 (.I0(n26796), .I1(n27045), .I2(n26292), 
            .I3(\data_in_frame[18] [5]), .O(n67232));
    defparam i3_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1404 (.I0(n61016), .I1(n25493), .I2(n62473), 
            .I3(n71892), .O(n71898));
    defparam i1_4_lut_adj_1404.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1405 (.I0(n69224), .I1(n69866), .I2(n71898), 
            .I3(n61366), .O(n67471));
    defparam i1_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1406 (.I0(\data_in_frame[17] [1]), .I1(n69479), 
            .I2(GND_net), .I3(GND_net), .O(n67135));
    defparam i1_2_lut_adj_1406.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(\data_in_frame[21] [6]), .I1(\data_in_frame[21] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n71920));
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1408 (.I0(n71920), .I1(n69235), .I2(n68596), 
            .I3(\data_in_frame[19][5] ), .O(n67064));
    defparam i1_4_lut_adj_1408.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(\data_in_frame[20][1] ), .I1(n69235), 
            .I2(GND_net), .I3(GND_net), .O(n67382));
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1410 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5050));
    defparam i4_4_lut_adj_1410.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1411 (.I0(\data_in[2] [7]), .I1(n10_adj_5050), 
            .I2(\data_in[3] [4]), .I3(GND_net), .O(n25915));
    defparam i5_3_lut_adj_1411.LUT_INIT = 16'hdfdf;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63596 (.I0(byte_transmit_counter_c[3]), 
            .I1(n77433), .I2(n75279), .I3(byte_transmit_counter_c[4]), 
            .O(n79510));
    defparam byte_transmit_counter_3__bdd_4_lut_63596.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_1412 (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5051));
    defparam i6_4_lut_adj_1412.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1413 (.I0(\data_in[1] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [3]), .O(n17_adj_5052));
    defparam i7_4_lut_adj_1413.LUT_INIT = 16'hfffd;
    SB_LUT4 i6_4_lut_adj_1414 (.I0(n67569), .I1(\data_in_frame[11]_c [5]), 
            .I2(n67422), .I3(\data_in_frame[13][7] ), .O(n14_adj_5053));
    defparam i6_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1415 (.I0(\data_out_frame[4] [2]), .I1(n66957), 
            .I2(\data_out_frame[6] [0]), .I3(n10_adj_4874), .O(n45));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1416 (.I0(n9_adj_4951), .I1(n14_adj_5053), .I2(n67468), 
            .I3(n62400), .O(n62342));
    defparam i7_4_lut_adj_1416.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1417 (.I0(n17_adj_5052), .I1(\data_in[3] [7]), 
            .I2(n16_adj_5051), .I3(\data_in[2] [6]), .O(n25956));
    defparam i9_4_lut_adj_1417.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_1418 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67246));
    defparam i1_2_lut_adj_1418.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1419 (.I0(\data_in_frame[11]_c [5]), .I1(n62392), 
            .I2(n26675), .I3(\data_in_frame[9] [3]), .O(n10_adj_5054));
    defparam i4_4_lut_adj_1419.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1420 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5055));
    defparam i2_2_lut_adj_1420.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1421 (.I0(n62348), .I1(n67246), .I2(n62342), 
            .I3(n61494), .O(n25493));
    defparam i3_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1422 (.I0(n62348), .I1(\data_in_frame[16][0] ), 
            .I2(\data_in_frame[17] [7]), .I3(n67043), .O(n10_adj_5056));
    defparam i4_4_lut_adj_1422.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1423 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5057));
    defparam i6_4_lut_adj_1423.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1424 (.I0(n26875), .I1(n69463), .I2(\data_in_frame[12][4] ), 
            .I3(n26418), .O(n62313));
    defparam i2_3_lut_4_lut_adj_1424.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1425 (.I0(\data_in[3] [6]), .I1(n14_adj_5057), 
            .I2(n10_adj_5055), .I3(\data_in[2] [1]), .O(n25909));
    defparam i7_4_lut_adj_1425.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1426 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n25909), .I3(\data_in[0] [5]), .O(n20_adj_5058));
    defparam i8_4_lut_adj_1426.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1427 (.I0(n25779), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_5059));
    defparam i7_4_lut_adj_1427.LUT_INIT = 16'hfeff;
    SB_LUT4 i56329_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [3]), .I2(\data_in[1] [2]), 
            .I3(\data_in[3] [2]), .O(n72176));
    defparam i56329_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_1428 (.I0(n72176), .I1(n19_adj_5059), .I2(n20_adj_5058), 
            .I3(GND_net), .O(n1951));
    defparam i11_3_lut_adj_1428.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_4_lut_adj_1429 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n26551), .I3(n62383), .O(n62404));
    defparam i1_2_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1430 (.I0(\data_in_frame[18] [3]), .I1(n25493), 
            .I2(GND_net), .I3(GND_net), .O(n61300));
    defparam i1_2_lut_adj_1430.LUT_INIT = 16'h6666;
    SB_LUT4 i56213_2_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n72057));
    defparam i56213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1431 (.I0(\data_in[3] [0]), .I1(\data_in[1] [5]), 
            .I2(n25915), .I3(n25909), .O(n18_adj_5060));
    defparam i7_4_lut_adj_1431.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1432 (.I0(\data_in_frame[20][4] ), .I1(\data_in_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5061));
    defparam i2_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1433 (.I0(n61300), .I1(\data_in_frame[18] [1]), 
            .I2(n6_adj_5061), .I3(n62329), .O(n67152));
    defparam i1_4_lut_adj_1433.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(\data_in_frame[14][6] ), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67364));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1435 (.I0(n62003), .I1(n67488), .I2(n67329), 
            .I3(n67519), .O(n68666));
    defparam i1_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1436 (.I0(n62307), .I1(n66942), .I2(n67416), 
            .I3(n67364), .O(n71738));
    defparam i1_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1437 (.I0(n71738), .I1(n71668), .I2(n62327), 
            .I3(n68666), .O(n69479));
    defparam i1_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1438 (.I0(n25956), .I1(\data_in[0] [3]), .I2(\data_in[1] [0]), 
            .I3(\data_in[2] [2]), .O(n19_adj_5062));
    defparam i8_4_lut_adj_1438.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1439 (.I0(n19_adj_5062), .I1(\data_in[0] [6]), 
            .I2(n18_adj_5060), .I3(n72057), .O(n1954));
    defparam i10_4_lut_adj_1439.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_adj_1440 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_5063));
    defparam i5_3_lut_adj_1440.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1441 (.I0(\data_in[0] [6]), .I1(n25915), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_5064));
    defparam i6_4_lut_adj_1441.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_3_lut_adj_1442 (.I0(n68596), .I1(n69479), .I2(\data_in_frame[19][4] ), 
            .I3(GND_net), .O(n69302));
    defparam i1_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1443 (.I0(n15_adj_5064), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5063), .I3(\data_in[0] [3]), .O(n25779));
    defparam i8_4_lut_adj_1443.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1444 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n25779), .O(n16_adj_5065));
    defparam i6_4_lut_adj_1444.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1445 (.I0(n25956), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5066));
    defparam i7_4_lut_adj_1445.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1446 (.I0(n17_adj_5066), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5065), .I3(\data_in[3] [3]), .O(n1957));
    defparam i9_4_lut_adj_1446.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1447 (.I0(n61404), .I1(n27243), .I2(\data_in_frame[14]_c [3]), 
            .I3(n67301), .O(n10_adj_5067));
    defparam i4_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i366_2_lut (.I0(n1954), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n1955));   // verilog/coms.v(142[4] 144[7])
    defparam i366_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_adj_1448 (.I0(\data_in_frame[9] [6]), .I1(n10_adj_5067), 
            .I2(n61345), .I3(GND_net), .O(n69042));
    defparam i5_3_lut_adj_1448.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1449 (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(GND_net), .I3(GND_net), .O(n66854));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1450 (.I0(\data_in_frame[14][2] ), .I1(n62356), 
            .I2(GND_net), .I3(GND_net), .O(n62473));
    defparam i1_2_lut_adj_1450.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5068));   // verilog/coms.v(217[11:56])
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1452 (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_5069));
    defparam i1_4_lut_adj_1452.LUT_INIT = 16'ha8a0;
    SB_LUT4 i31299_4_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4_adj_5069), .I3(n4_adj_5068), .O(n45392));
    defparam i31299_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i2_4_lut_adj_1453 (.I0(n66854), .I1(n1955), .I2(n1957), .I3(\FRAME_MATCHER.i_31__N_2507 ), 
            .O(n6_adj_5070));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1453.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_4_lut_adj_1454 (.I0(n33), .I1(n26813), .I2(\data_out_frame[10] [7]), 
            .I3(\data_out_frame[15] [5]), .O(n6_adj_4873));
    defparam i1_2_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1455 (.I0(n26760), .I1(n61396), .I2(GND_net), 
            .I3(GND_net), .O(n66889));
    defparam i1_2_lut_adj_1455.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1456 (.I0(n69824), .I1(n6_adj_5070), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n79682));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1456.LUT_INIT = 16'hefee;
    SB_LUT4 n79510_bdd_4_lut (.I0(n79510), .I1(n79183), .I2(n7_adj_5071), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[2]));
    defparam n79510_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(\data_in_frame[16]_c [6]), .I1(n26760), 
            .I2(n61396), .I3(GND_net), .O(n62383));
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1458 (.I0(n33), .I1(n26813), .I2(\data_out_frame[10] [7]), 
            .I3(n67530), .O(n6_adj_4865));
    defparam i1_2_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1459 (.I0(n26551), .I1(n62383), .I2(GND_net), 
            .I3(GND_net), .O(n67316));
    defparam i1_2_lut_adj_1459.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1460 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26292));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1460.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1461 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[12][4] ), 
            .I2(\data_in_frame[14][7] ), .I3(n67385), .O(n67416));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1462 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[9] [7]), 
            .I2(n67265), .I3(GND_net), .O(n27243));
    defparam i1_3_lut_adj_1462.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1463 (.I0(n27243), .I1(n67416), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5072));
    defparam i1_2_lut_adj_1463.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1464 (.I0(\data_in_frame[19][6] ), .I1(n68596), 
            .I2(n69479), .I3(\data_in_frame[19][4] ), .O(n67298));
    defparam i1_2_lut_4_lut_adj_1464.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1465 (.I0(\data_in_frame[16][7] ), .I1(\data_in_frame[14][5] ), 
            .I2(n67028), .I3(n6_adj_5072), .O(n25507));
    defparam i4_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\data_in_frame[14][6] ), .I1(\data_in_frame[16][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5073));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1467 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[16]_c [6]), 
            .I2(n62313), .I3(n6_adj_5073), .O(n67310));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[19][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66932));
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1469 (.I0(n26760), .I1(n67310), .I2(n25507), 
            .I3(\data_in_frame[17] [1]), .O(n62406));
    defparam i3_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1470 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n71966));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1470.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1471 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[6] [3]), .I3(\data_in_frame[8] [4]), .O(n71970));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1471.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1472 (.I0(\data_in_frame[1][7] ), .I1(n71970), 
            .I2(n71966), .I3(\data_in_frame[1][6] ), .O(n71974));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1473 (.I0(n26261), .I1(n67563), .I2(n71974), 
            .I3(n67566), .O(n71980));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1474 (.I0(n67079), .I1(n61427), .I2(n71980), 
            .I3(n67179), .O(n67569));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1474.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1475 (.I0(n61404), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n67268));
    defparam i1_2_lut_adj_1475.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1476 (.I0(n67117), .I1(\data_in_frame[14] [0]), 
            .I2(n26364), .I3(GND_net), .O(n67238));
    defparam i2_3_lut_adj_1476.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1477 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[7] [1]), .I3(\data_in_frame[5] [0]), .O(n71938));
    defparam i1_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1478 (.I0(n27073), .I1(n67091), .I2(n71942), 
            .I3(n67441), .O(n71948));
    defparam i1_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1479 (.I0(n67268), .I1(n67322), .I2(n67114), 
            .I3(n71948), .O(n71954));
    defparam i1_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1480 (.I0(n71766), .I1(n67569), .I2(n67596), 
            .I3(n71954), .O(n62356));
    defparam i1_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63591 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n79504));
    defparam byte_transmit_counter_0__bdd_4_lut_63591.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1481 (.I0(\data_in_frame[13][7] ), .I1(n67459), 
            .I2(GND_net), .I3(GND_net), .O(n67043));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1481.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1482 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[13][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n67235));
    defparam i1_2_lut_adj_1482.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1483 (.I0(\data_in_frame[13] [1]), .I1(n62034), 
            .I2(n6_adj_5042), .I3(n26418), .O(n67459));
    defparam i1_4_lut_adj_1483.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1484 (.I0(\data_in_frame[11]_c [6]), .I1(n24270), 
            .I2(n26100), .I3(n26848), .O(n67117));
    defparam i3_4_lut_adj_1484.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1485 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[16][0] ), .I3(\data_in_frame[16] [1]), .O(n18_adj_5074));
    defparam i7_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1486 (.I0(\data_in_frame[13][5] ), .I1(\data_in_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5075));
    defparam i5_2_lut_adj_1486.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1487 (.I0(n61494), .I1(n18_adj_5074), .I2(n30_adj_5076), 
            .I3(n67459), .O(n20_adj_5077));
    defparam i9_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1488 (.I0(\FRAME_MATCHER.i [5]), .I1(n89), 
            .I2(n8_adj_5078), .I3(n66835), .O(n69075));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1488.LUT_INIT = 16'hfffb;
    SB_LUT4 i10_4_lut_adj_1489 (.I0(n67117), .I1(n20_adj_5077), .I2(n16_adj_5075), 
            .I3(\data_in_frame[13][6] ), .O(n69589));
    defparam i10_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 n79504_bdd_4_lut (.I0(n79504), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n79507));
    defparam n79504_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1490 (.I0(n7_adj_5079), .I1(\data_in_frame[14][2] ), 
            .I2(n62356), .I3(n67238), .O(n67497));
    defparam i4_4_lut_adj_1490.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1491 (.I0(\FRAME_MATCHER.i [5]), .I1(n89), 
            .I2(n3476), .I3(GND_net), .O(n41637));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1491.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_adj_1492 (.I0(n67497), .I1(\data_in_frame[16] [3]), 
            .I2(n69589), .I3(GND_net), .O(n61366));
    defparam i2_3_lut_adj_1492.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1493 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26796));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1493.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1494 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[8] [6]), .O(n33));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1495 (.I0(n62392), .I1(n26345), .I2(n26959), 
            .I3(\data_in_frame[17] [2]), .O(n71668));
    defparam i1_3_lut_4_lut_adj_1495.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1496 (.I0(control_mode[1]), .I1(control_mode[0]), 
            .I2(n53108), .I3(n105), .O(n4));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_adj_1496.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_adj_1497 (.I0(n26345), .I1(n26959), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_5076));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1497.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1498 (.I0(\data_in_frame[20][2] ), .I1(n30_adj_5076), 
            .I2(n66945), .I3(\data_in_frame[13][4] ), .O(n67539));
    defparam i3_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1499 (.I0(control_mode[1]), .I1(control_mode[0]), 
            .I2(n53108), .I3(control_update), .O(n25921));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_adj_1499.LUT_INIT = 16'h08ff;
    SB_LUT4 i5_3_lut_4_lut_adj_1500 (.I0(\data_in_frame[13][0] ), .I1(n26418), 
            .I2(n10_adj_5054), .I3(n67268), .O(n62348));
    defparam i5_3_lut_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1501 (.I0(n26246), .I1(n26776), .I2(n67225), 
            .I3(n67385), .O(n67519));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1502 (.I0(\data_in_frame[19][3] ), .I1(n25507), 
            .I2(\data_in_frame[17] [1]), .I3(n69479), .O(n61424));
    defparam i1_3_lut_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1503 (.I0(n67519), .I1(n67294), .I2(\data_in_frame[13] [1]), 
            .I3(\data_in_frame[15] [3]), .O(n69062));
    defparam i1_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1504 (.I0(\data_in_frame[15] [3]), .I1(n62321), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n69235));
    defparam i1_3_lut_adj_1504.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(\data_in_frame[15][5] ), .I1(n24167), 
            .I2(GND_net), .I3(GND_net), .O(n67283));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1506 (.I0(n67294), .I1(n62327), .I2(\data_in_frame[15] [4]), 
            .I3(\data_in_frame[13] [3]), .O(n69576));
    defparam i1_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i15665_3_lut_4_lut (.I0(n28692), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29879));
    defparam i15665_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4960));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1507 (.I0(n26345), .I1(n26364), .I2(GND_net), 
            .I3(GND_net), .O(n67329));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1507.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(GND_net), .I3(GND_net), .O(n27073));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4959));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1509 (.I0(n26323), .I1(n67456), .I2(n67409), 
            .I3(n67406), .O(n26345));
    defparam i3_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4958));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4939));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_787_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4938));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15662_3_lut_4_lut (.I0(n28692), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n29876));
    defparam i15662_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16125_3_lut_4_lut (.I0(n28672), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[12][5] ), .O(n30339));
    defparam i16125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4957));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i62419_3_lut_4_lut (.I0(n28692), .I1(reset), .I2(\data_in_frame[0] [4]), 
            .I3(rx_data[4]), .O(n66132));
    defparam i62419_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i2_2_lut_adj_1510 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5081));
    defparam i2_2_lut_adj_1510.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1511 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26100));
    defparam i1_2_lut_adj_1511.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1512 (.I0(\data_in_frame[9] [6]), .I1(n26655), 
            .I2(\data_in_frame[9] [7]), .I3(n6_adj_5040), .O(n67032));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4956));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i62418_3_lut_4_lut (.I0(n28692), .I1(reset), .I2(\data_in_frame[0] [3]), 
            .I3(rx_data[3]), .O(n66084));
    defparam i62418_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n71990));   // verilog/coms.v(74[16:69])
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1514 (.I0(Kp_23__N_767), .I1(n26190), .I2(n71990), 
            .I3(\data_in_frame[0] [7]), .O(n71996));   // verilog/coms.v(74[16:69])
    defparam i1_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i15562_3_lut_4_lut (.I0(n28692), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29776));
    defparam i15562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1515 (.I0(n67019), .I1(n71996), .I2(n67403), 
            .I3(n26585), .O(n61404));   // verilog/coms.v(88[17:70])
    defparam i1_4_lut_adj_1515.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(Kp_23__N_993), .I1(n61404), .I2(GND_net), 
            .I3(GND_net), .O(n67422));
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(n61345), .I1(n67032), .I2(GND_net), 
            .I3(GND_net), .O(n71766));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4933));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1518 (.I0(n71766), .I1(n26246), .I2(n25469), 
            .I3(\data_in_frame[9] [0]), .O(n61427));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1519 (.I0(n67111), .I1(n26675), .I2(n71776), 
            .I3(n7_adj_5082), .O(n71782));
    defparam i1_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4932));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16549_3_lut_4_lut (.I0(n28692), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n30763));
    defparam i16549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1520 (.I0(n67422), .I1(n67554), .I2(n24270), 
            .I3(n71782), .O(n25469));
    defparam i1_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1521 (.I0(n25469), .I1(n61427), .I2(n61345), 
            .I3(GND_net), .O(n69556));
    defparam i1_3_lut_adj_1521.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4955));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_4_lut_adj_1522 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n25879), .I3(\FRAME_MATCHER.i[1] ), .O(n5_adj_5049));
    defparam i1_3_lut_4_lut_adj_1522.LUT_INIT = 16'hfefc;
    SB_LUT4 select_787_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4931));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1523 (.I0(n7_adj_5081), .I1(n69556), .I2(n67032), 
            .I3(\data_in_frame[11]_c [1]), .O(n67419));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1523.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1524 (.I0(n26776), .I1(n67419), .I2(n26331), 
            .I3(\data_in_frame[10] [6]), .O(n62003));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1525 (.I0(\data_in_frame[19] [0]), .I1(n62365), 
            .I2(n26292), .I3(n67316), .O(n24227));
    defparam i2_3_lut_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4954));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_in_frame[13][2] ), .I1(n62003), 
            .I2(GND_net), .I3(GND_net), .O(n67294));
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1527 (.I0(n26317), .I1(n27225), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n4_adj_5083));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1527.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1528 (.I0(\data_in_frame[12][5] ), .I1(n26875), 
            .I2(GND_net), .I3(GND_net), .O(n66985));
    defparam i1_2_lut_adj_1528.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4928));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1529 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5084));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1529.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4927));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4926));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1530 (.I0(\data_in_frame[13][5] ), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n71658));
    defparam i1_2_lut_adj_1530.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1531 (.I0(n27_adj_5084), .I1(n62266), .I2(n71658), 
            .I3(\data_in_frame[13][2] ), .O(n62392));
    defparam i1_4_lut_adj_1531.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1532 (.I0(\data_in_frame[13][0] ), .I1(n26418), 
            .I2(GND_net), .I3(GND_net), .O(n26872));
    defparam i1_2_lut_adj_1532.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1533 (.I0(n26779), .I1(n67198), .I2(n66918), 
            .I3(\data_in_frame[1] [4]), .O(n27225));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4923));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1534 (.I0(\data_in_frame[8] [5]), .I1(n67099), 
            .I2(n44_adj_5085), .I3(\data_in_frame[6] [3]), .O(n26246));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1535 (.I0(\data_in_frame[8] [3]), .I1(n35_adj_5086), 
            .I2(\data_in_frame[6] [2]), .I3(n26317), .O(n26818));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(n26818), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n66991));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4921));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1537 (.I0(n26282), .I1(n27225), .I2(n61345), 
            .I3(GND_net), .O(n67265));
    defparam i2_3_lut_adj_1537.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1538 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26655));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1538.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1539 (.I0(\data_in_frame[12][3] ), .I1(\data_in_frame[12][5] ), 
            .I2(\data_in_frame[12][6] ), .I3(GND_net), .O(n67028));
    defparam i2_3_lut_adj_1539.LUT_INIT = 16'h9696;
    SB_LUT4 i56202_3_lut_4_lut (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [6]), .I3(n26724), .O(n72045));
    defparam i56202_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i1_2_lut_adj_1540 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67301));
    defparam i1_2_lut_adj_1540.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1541 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(Kp_23__N_767), .I3(\data_in_frame[1] [0]), .O(n26585));
    defparam i1_2_lut_3_lut_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i16008_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n30222));
    defparam i16008_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16011_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n30225));
    defparam i16011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16014_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n30228));
    defparam i16014_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16017_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n30231));
    defparam i16017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16020_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n30234));
    defparam i16020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1542 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n67225));
    defparam i1_2_lut_adj_1542.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1543 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n67179));
    defparam i1_2_lut_adj_1543.LUT_INIT = 16'h6666;
    SB_LUT4 i16023_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n30237));
    defparam i16023_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1544 (.I0(n26687), .I1(n26848), .I2(GND_net), 
            .I3(GND_net), .O(n27117));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1544.LUT_INIT = 16'h6666;
    SB_LUT4 i16026_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n30240));
    defparam i16026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1545 (.I0(n26986), .I1(\data_in_frame[5] [2]), 
            .I2(\data_in_frame[5] [3]), .I3(n67173), .O(n10_adj_5037));
    defparam i4_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1546 (.I0(n26585), .I1(n10_adj_5037), .I2(\data_in_frame[7] [4]), 
            .I3(GND_net), .O(n67114));
    defparam i5_3_lut_adj_1546.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1547 (.I0(n24270), .I1(\data_in_frame[9] [7]), 
            .I2(n24274), .I3(GND_net), .O(n67079));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1547.LUT_INIT = 16'h9696;
    SB_LUT4 i16029_3_lut_4_lut (.I0(n8_adj_5), .I1(n66868), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n30243));
    defparam i16029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1548 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n67566));
    defparam i1_2_lut_adj_1548.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1549 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[16] [0]), .I3(\data_out_frame[13] [6]), 
            .O(n6_adj_4795));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 equal_304_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_10));   // verilog/coms.v(157[7:23])
    defparam equal_304_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1550 (.I0(\data_in_frame[5] [5]), .I1(n26299), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5088));
    defparam i1_2_lut_adj_1550.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1551 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [3]), 
            .I2(n26286), .I3(n6_adj_5088), .O(n67105));
    defparam i4_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1552 (.I0(\data_in_frame[7] [7]), .I1(n67105), 
            .I2(\data_in_frame[1][5] ), .I3(GND_net), .O(n26261));
    defparam i2_3_lut_adj_1552.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1553 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26779));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1553.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_adj_1554 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5));   // verilog/coms.v(157[7:23])
    defparam i2_2_lut_3_lut_adj_1554.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1555 (.I0(n26139), .I1(\data_in_frame[7] [6]), 
            .I2(n26299), .I3(GND_net), .O(n24274));
    defparam i2_3_lut_adj_1555.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1556 (.I0(n161), .I1(n66835), .I2(n10_adj_4866), 
            .I3(GND_net), .O(n66860));
    defparam i1_2_lut_3_lut_adj_1556.LUT_INIT = 16'hfdfd;
    SB_LUT4 i3_4_lut_adj_1557 (.I0(\data_in_frame[8] [0]), .I1(n67462), 
            .I2(n67142), .I3(n26779), .O(n26282));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1557.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1558 (.I0(n26282), .I1(n69356), .I2(n24274), 
            .I3(\data_in_frame[8] [1]), .O(n67412));
    defparam i1_4_lut_adj_1558.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1559 (.I0(n161), .I1(n66835), .I2(n10_adj_5089), 
            .I3(GND_net), .O(n66868));
    defparam i1_2_lut_3_lut_adj_1559.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1560 (.I0(n67105), .I1(n62400), .I2(GND_net), 
            .I3(GND_net), .O(n62438));
    defparam i1_2_lut_adj_1560.LUT_INIT = 16'h6666;
    SB_LUT4 i15983_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n30197));
    defparam i15983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1561 (.I0(n62438), .I1(n67412), .I2(\data_in_frame[7] [7]), 
            .I3(\data_in_frame[10] [2]), .O(n69463));
    defparam i1_4_lut_adj_1561.LUT_INIT = 16'h9669;
    SB_LUT4 i15986_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n30200));
    defparam i15986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(n67352), .I1(n67566), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5090));
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1563 (.I0(\data_in_frame[10] [3]), .I1(n67198), 
            .I2(n67462), .I3(n6_adj_5090), .O(n26875));
    defparam i4_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 i15989_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n30203));
    defparam i15989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(n26875), .I1(n69463), .I2(GND_net), 
            .I3(GND_net), .O(n62307));
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h9999;
    SB_LUT4 i15992_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n30206));
    defparam i15992_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15995_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n30209));
    defparam i15995_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15998_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n30212));
    defparam i15998_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16001_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n30215));
    defparam i16001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11]_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n67146));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1566 (.I0(\data_in_frame[11]_c [1]), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[11]_c [4]), .I3(\data_in_frame[11]_c [0]), 
            .O(n71590));
    defparam i1_4_lut_adj_1566.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1567 (.I0(n71590), .I1(n67146), .I2(\data_in_frame[9] [0]), 
            .I3(\data_in_frame[10] [4]), .O(n71596));
    defparam i1_4_lut_adj_1567.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1568 (.I0(n67560), .I1(n71596), .I2(n67179), 
            .I3(n67225), .O(n71600));
    defparam i1_4_lut_adj_1568.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(n67578), .I1(n67406), .I2(GND_net), 
            .I3(GND_net), .O(n71602));
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1570 (.I0(Kp_23__N_993), .I1(Kp_23__N_974), .I2(n71602), 
            .I3(n71600), .O(n71608));
    defparam i1_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 i16005_3_lut_4_lut (.I0(n45283), .I1(n66860), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n30219));
    defparam i16005_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15717_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29931));
    defparam i15717_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15714_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29928));
    defparam i15714_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1571 (.I0(n67265), .I1(n67515), .I2(n71608), 
            .I3(n66991), .O(n71614));
    defparam i1_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i15711_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29925));
    defparam i15711_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1572 (.I0(n67554), .I1(n62307), .I2(n67243), 
            .I3(n71614), .O(n62034));
    defparam i1_4_lut_adj_1572.LUT_INIT = 16'h9669;
    SB_LUT4 i15708_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29922));
    defparam i15708_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15705_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29919));
    defparam i15705_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15702_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29916));
    defparam i15702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1573 (.I0(\data_in_frame[13][0] ), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n71796));
    defparam i1_2_lut_adj_1573.LUT_INIT = 16'h6666;
    SB_LUT4 i15697_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29911));
    defparam i15697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1574 (.I0(n67001), .I1(n67453), .I2(\data_out_frame[18] [4]), 
            .I3(GND_net), .O(n61406));
    defparam i1_2_lut_3_lut_adj_1574.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1575 (.I0(n67584), .I1(n67294), .I2(n66942), 
            .I3(n71796), .O(n62321));
    defparam i1_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1576 (.I0(n62266), .I1(n24167), .I2(\data_in_frame[15] [1]), 
            .I3(GND_net), .O(n67213));
    defparam i1_3_lut_adj_1576.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1577 (.I0(\data_in_frame[14][7] ), .I1(n26872), 
            .I2(n62392), .I3(n26364), .O(n67488));
    defparam i1_4_lut_adj_1577.LUT_INIT = 16'h9669;
    SB_LUT4 i15739_3_lut_4_lut (.I0(n8_adj_11), .I1(n66860), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29953));
    defparam i15739_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1578 (.I0(n67001), .I1(n67453), .I2(n26203), 
            .I3(n60995), .O(n69543));
    defparam i2_3_lut_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1579 (.I0(\FRAME_MATCHER.i [5]), .I1(n8_adj_10), 
            .I2(n82), .I3(GND_net), .O(n28715));
    defparam i1_2_lut_3_lut_adj_1579.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut_adj_1580 (.I0(n67488), .I1(n67213), .I2(n62321), 
            .I3(n71760), .O(n68596));
    defparam i1_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(n69235), .I1(n69576), .I2(n69062), 
            .I3(\data_in_frame[17] [5]), .O(n68717));
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'h9669;
    SB_LUT4 i59849_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n8_adj_10), 
            .I2(n89), .I3(n3476), .O(n75246));
    defparam i59849_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 equal_311_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_11));   // verilog/coms.v(157[7:23])
    defparam equal_311_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_310_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5078));   // verilog/coms.v(157[7:23])
    defparam equal_310_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_3_lut_adj_1582 (.I0(n67284), .I1(\data_in_frame[17] [6]), 
            .I2(\data_in_frame[20][0] ), .I3(GND_net), .O(n66988));
    defparam i2_3_lut_adj_1582.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1583 (.I0(n68717), .I1(n68596), .I2(GND_net), 
            .I3(GND_net), .O(n27203));
    defparam i1_2_lut_adj_1583.LUT_INIT = 16'h6666;
    SB_LUT4 i15803_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n30017));
    defparam i15803_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15883_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n30097));
    defparam i15883_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1584 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[4] [6]), .I3(GND_net), .O(n67170));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1584.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1585 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[1] [4]), .O(n69802));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1585.LUT_INIT = 16'h6996;
    SB_LUT4 i15800_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n30014));
    defparam i15800_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15795_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n30009));
    defparam i15795_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1586 (.I0(n26296), .I1(n44_adj_5085), .I2(n35_adj_5086), 
            .I3(\data_in_frame[8] [4]), .O(n26331));
    defparam i3_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(n26585), .I1(n67338), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5092));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1588 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[5] [4]), 
            .I2(n66964), .I3(n6_adj_5092), .O(n61345));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1588.LUT_INIT = 16'h6996;
    SB_LUT4 i15790_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n30004));
    defparam i15790_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15906_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n30120));
    defparam i15906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1589 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n14_adj_5093));
    defparam i5_3_lut_adj_1589.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1590 (.I0(n67067), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[2] [5]), .I3(n66974), .O(n15_adj_5094));
    defparam i6_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1591 (.I0(n15_adj_5094), .I1(\data_in_frame[2] [7]), 
            .I2(n14_adj_5093), .I3(\data_in_frame[4] [6]), .O(n26848));
    defparam i8_4_lut_adj_1591.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1592 (.I0(n26721), .I1(n67170), .I2(n26724), 
            .I3(n27052), .O(n26687));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1592.LUT_INIT = 16'h6996;
    SB_LUT4 i15766_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29980));
    defparam i15766_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15748_3_lut_4_lut (.I0(n8_adj_5078), .I1(n66860), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29962));
    defparam i15748_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1593 (.I0(\data_in_frame[1][5] ), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n66918));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1593.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1594 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26323));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_adj_1594.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1595 (.I0(\data_in_frame[6] [0]), .I1(n67465), 
            .I2(GND_net), .I3(GND_net), .O(n67091));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1595.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1596 (.I0(\FRAME_MATCHER.i[0] ), .I1(n44662), 
            .I2(n41637), .I3(reset), .O(n66853));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1596.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_adj_1597 (.I0(\data_in_frame[4] [5]), .I1(n61339), 
            .I2(GND_net), .I3(GND_net), .O(n67322));
    defparam i1_2_lut_adj_1597.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1598 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67070));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1598.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1599 (.I0(\data_in_frame[1][7] ), .I1(n67070), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[4] [4]), .O(n67441));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1599.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1600 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[2] [0]), 
            .I2(n67185), .I3(n26752), .O(n67099));   // verilog/coms.v(76[16:42])
    defparam i3_4_lut_adj_1600.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1601 (.I0(\data_in_frame[4] [7]), .I1(n27048), 
            .I2(GND_net), .I3(GND_net), .O(n67019));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1601.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1602 (.I0(\data_in_frame[7] [1]), .I1(n67019), 
            .I2(n27052), .I3(n26718), .O(n67409));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1602.LUT_INIT = 16'h6996;
    SB_LUT4 equal_306_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_5089));   // verilog/coms.v(158[12:15])
    defparam equal_306_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1603 (.I0(Kp_23__N_799), .I1(n67322), .I2(n67091), 
            .I3(n26323), .O(n62400));   // verilog/coms.v(88[17:28])
    defparam i1_4_lut_adj_1603.LUT_INIT = 16'h6996;
    SB_LUT4 equal_314_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4866));   // verilog/coms.v(158[12:15])
    defparam equal_314_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1604 (.I0(\data_in_frame[4] [5]), .I1(n67409), 
            .I2(GND_net), .I3(GND_net), .O(n26675));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1604.LUT_INIT = 16'h6666;
    SB_LUT4 equal_2036_i7_2_lut (.I0(Kp_23__N_974), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5082));   // verilog/coms.v(239[9:81])
    defparam equal_2036_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1605 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26296));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1605.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1606 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n26286));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1606.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1607 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[3] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66974));
    defparam i1_2_lut_adj_1607.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1608 (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_4936), 
            .I2(n67716), .I3(n10_adj_5089), .O(n28672));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1608.LUT_INIT = 16'hffef;
    SB_LUT4 i14112_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n133[0]), .I2(n3476), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n28325));   // verilog/coms.v(158[12:15])
    defparam i14112_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_4_lut_adj_1609 (.I0(\data_in_frame[1][1] ), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[3] [2]), .O(n67173));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1609.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1610 (.I0(\data_in_frame[5] [4]), .I1(n67173), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n26139));
    defparam i1_3_lut_adj_1610.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1611 (.I0(\data_in_frame[5] [0]), .I1(Kp_23__N_799), 
            .I2(GND_net), .I3(GND_net), .O(n26718));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1611.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1612 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1][3] ), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n26299));   // verilog/coms.v(79[16:43])
    defparam i1_3_lut_adj_1612.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1613 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n66848), .I3(LED_c), .O(n27770));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1613.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_1614 (.I0(\data_in_frame[5] [6]), .I1(n26299), 
            .I2(GND_net), .I3(GND_net), .O(n67198));
    defparam i1_2_lut_adj_1614.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1615 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3476));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1615.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1616 (.I0(\data_in_frame[1][5] ), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n67182));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1616.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1617 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67403));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1617.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1618 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[5] [3]), .O(n66964));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n72502), .I3(n72500), .O(n7_adj_5071));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1619 (.I0(\data_in_frame[1][3] ), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n67142));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1619.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1620 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[4] [4]), .I3(\data_in_frame[4] [0]), .O(n71682));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1620.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n72508), .I3(n72506), .O(n7_adj_5038));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_4_lut_adj_1621 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(\data_in_frame[4] [6]), .I3(\data_in_frame[4] [7]), .O(n71684));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1621.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1622 (.I0(n71684), .I1(Kp_23__N_753), .I2(n71682), 
            .I3(GND_net), .O(n71690));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_adj_1622.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1623 (.I0(n26190), .I1(n71690), .I2(n67182), 
            .I3(n66982), .O(n71694));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1623.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1624 (.I0(n67185), .I1(n67198), .I2(n71706), 
            .I3(n71704), .O(n71712));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1624.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1625 (.I0(n26718), .I1(n26139), .I2(n71694), 
            .I3(n26724), .O(n71700));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1626 (.I0(n26986), .I1(n71700), .I2(n71712), 
            .I3(n26585), .O(n61339));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1626.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n72487), .I3(n72485), .O(n7_adj_4914));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n72466), .I3(n72464), .O(n7_adj_4868));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i3_4_lut_adj_1627 (.I0(\data_in_frame[6] [1]), .I1(n26296), 
            .I2(\data_in_frame[6] [7]), .I3(\data_in_frame[6] [4]), .O(n67465));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1627.LUT_INIT = 16'h6996;
    SB_LUT4 i56630_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72486));
    defparam i56630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1628 (.I0(n67465), .I1(n61339), .I2(\data_in_frame[3] [6]), 
            .I3(n67142), .O(n15_adj_5095));   // verilog/coms.v(73[16:69])
    defparam i6_4_lut_adj_1628.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1629 (.I0(n15_adj_5095), .I1(n66918), .I2(n14_adj_5096), 
            .I3(n26724), .O(n69633));   // verilog/coms.v(73[16:69])
    defparam i8_4_lut_adj_1629.LUT_INIT = 16'h6996;
    SB_LUT4 i56631_4_lut (.I0(n72486), .I1(n28443), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][5] ), .O(n72487));
    defparam i56631_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i56629_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n72485));
    defparam i56629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1630 (.I0(n7_adj_5082), .I1(n26675), .I2(n69356), 
            .I3(\data_in_frame[8] [0]), .O(n69451));
    defparam i2_4_lut_adj_1630.LUT_INIT = 16'h1001;
    SB_LUT4 i56345_4_lut (.I0(n26687), .I1(n26848), .I2(n61345), .I3(n26331), 
            .O(n72192));
    defparam i56345_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1631 (.I0(n24274), .I1(n69633), .I2(n69421), 
            .I3(n24270), .O(n24_adj_5097));
    defparam i9_4_lut_adj_1631.LUT_INIT = 16'h0200;
    SB_LUT4 i10_4_lut_adj_1632 (.I0(n69451), .I1(n7_adj_5081), .I2(n26246), 
            .I3(n26818), .O(n25));
    defparam i10_4_lut_adj_1632.LUT_INIT = 16'h0002;
    SB_LUT4 i8_4_lut_adj_1633 (.I0(n4_adj_5083), .I1(n61404), .I2(n62438), 
            .I3(\data_in_frame[7] [7]), .O(n23_adj_5098));
    defparam i8_4_lut_adj_1633.LUT_INIT = 16'h0440;
    SB_LUT4 i14_4_lut_adj_1634 (.I0(n23_adj_5098), .I1(n25), .I2(n24_adj_5097), 
            .I3(n72192), .O(LED_N_3408));
    defparam i14_4_lut_adj_1634.LUT_INIT = 16'h0080;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n72478), .I3(n72476), .O(n7_adj_4888));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i16211_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n30425));
    defparam i16211_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16208_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n30422));
    defparam i16208_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1635 (.I0(n27203), .I1(\data_in_frame[22] [1]), 
            .I2(\data_in_frame[21] [7]), .I3(n66988), .O(n10_adj_5099));
    defparam i4_4_lut_adj_1635.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1636 (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[18] [2]), 
            .I2(n67149), .I3(GND_net), .O(n8_adj_5100));
    defparam i3_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i16204_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(rx_data[5]), 
            .I3(\data_in_frame[15][5] ), .O(n30418));
    defparam i16204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i23_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(\data_in_frame[15] [4]), 
            .I3(rx_data[4]), .O(n15_adj_4949));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i16198_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n30412));
    defparam i16198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1637 (.I0(\data_in_frame[20][4] ), .I1(n69421), 
            .I2(n6_adj_5036), .I3(n61366), .O(n71628));
    defparam i1_4_lut_adj_1637.LUT_INIT = 16'h2112;
    SB_LUT4 i16194_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n30408));
    defparam i16194_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16191_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n30405));
    defparam i16191_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1638 (.I0(n62406), .I1(\data_in_frame[21] [3]), 
            .I2(\data_in_frame[23] [4]), .I3(n66932), .O(n10_adj_5101));
    defparam i4_4_lut_adj_1638.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1639 (.I0(n69589), .I1(n71628), .I2(n8_adj_5100), 
            .I3(\data_in_frame[22] [4]), .O(n71630));
    defparam i1_4_lut_adj_1639.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut_adj_1640 (.I0(n62404), .I1(n71630), .I2(n10_adj_5101), 
            .I3(\data_in_frame[21] [2]), .O(n71632));
    defparam i1_4_lut_adj_1640.LUT_INIT = 16'h4884;
    SB_LUT4 i5_3_lut_adj_1641 (.I0(\data_in_frame[19][7] ), .I1(n10_adj_5099), 
            .I2(\data_in_frame[19][5] ), .I3(GND_net), .O(n69188));
    defparam i5_3_lut_adj_1641.LUT_INIT = 16'h9696;
    SB_LUT4 i16188_3_lut_4_lut (.I0(n45283), .I1(n66868), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n30402));
    defparam i16188_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_3_lut_adj_1642 (.I0(\data_in_frame[21] [7]), .I1(n68717), 
            .I2(n67298), .I3(GND_net), .O(n8_adj_5102));
    defparam i3_3_lut_adj_1642.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1643 (.I0(n69188), .I1(\data_in_frame[22] [5]), 
            .I2(n71632), .I3(n67152), .O(n71636));
    defparam i1_4_lut_adj_1643.LUT_INIT = 16'h4010;
    SB_LUT4 i4_4_lut_adj_1644 (.I0(\data_in_frame[19][2] ), .I1(n69302), 
            .I2(\data_in_frame[23] [6]), .I3(\data_in_frame[21] [5]), .O(n10_adj_5103));
    defparam i4_4_lut_adj_1644.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(\data_in_frame[22] [0]), .I1(n71636), 
            .I2(n8_adj_5102), .I3(\data_in_frame[21] [6]), .O(n71638));
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n71638), .I1(\data_in_frame[21] [4]), 
            .I2(n10_adj_5103), .I3(n62406), .O(n71640));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(n61424), .I1(n71640), .I2(n67064), 
            .I3(\data_in_frame[23] [7]), .O(n71642));
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut_adj_1648 (.I0(n67382), .I1(n62329), .I2(\data_in_frame[19][6] ), 
            .I3(\data_in_frame[22] [2]), .O(n71908));
    defparam i1_4_lut_adj_1648.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1649 (.I0(n71642), .I1(\data_in_frame[23] [5]), 
            .I2(n67191), .I3(n61424), .O(n71644));
    defparam i1_4_lut_adj_1649.LUT_INIT = 16'h2882;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[20][1] ), 
            .I2(\data_in_frame[19][7] ), .I3(\data_in_frame[22] [3]), .O(n71916));
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n66988), .I1(n71644), .I2(n67471), 
            .I3(n71908), .O(n71646));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1652 (.I0(n71646), .I1(n67149), .I2(n67471), 
            .I3(n71916), .O(n71648));
    defparam i1_4_lut_adj_1652.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(n24227), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[23] [3]), .I3(\data_in_frame[21] [2]), .O(n71886));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1654 (.I0(n66970), .I1(n71648), .I2(Kp_23__N_1607), 
            .I3(\data_in_frame[23] [1]), .O(n71650));
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'h8448;
    SB_LUT4 i1_3_lut_adj_1655 (.I0(\data_in_frame[21] [1]), .I1(n61755), 
            .I2(\data_in_frame[23] [2]), .I3(GND_net), .O(n69696));
    defparam i1_3_lut_adj_1655.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4912));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4911));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1656 (.I0(n69696), .I1(n71650), .I2(n71886), 
            .I3(Kp_23__N_1607), .O(n71654));
    defparam i1_4_lut_adj_1656.LUT_INIT = 16'h0880;
    SB_LUT4 select_787_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4910));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1657 (.I0(n67373), .I1(n61300), .I2(\data_in_frame[20] [5]), 
            .I3(\data_in_frame[22] [7]), .O(n71568));
    defparam i1_4_lut_adj_1657.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4909));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1658 (.I0(\data_in_frame[23] [0]), .I1(n71654), 
            .I2(n61755), .I3(n66970), .O(n71656));
    defparam i1_4_lut_adj_1658.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(n71656), .I1(n71568), .I2(n61755), 
            .I3(n66970), .O(Kp_23__N_612));
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'h2882;
    SB_LUT4 select_787_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4908));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1660 (.I0(n26783), .I1(n27089), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[13] [6]), .O(n67001));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1660.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4907));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1661 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(n61294), .I3(n67075), .O(n61412));
    defparam i2_3_lut_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4906));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(\data_out_frame[24] [6]), .I3(GND_net), .O(n17_adj_4861));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1662 (.I0(\data_out_frame[20] [2]), .I1(n61333), 
            .I2(\data_out_frame[20] [3]), .I3(n69502), .O(n24023));
    defparam i1_2_lut_3_lut_4_lut_adj_1662.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1663 (.I0(\data_out_frame[20] [2]), .I1(n61333), 
            .I2(n68641), .I3(\data_out_frame[22] [3]), .O(n25458));
    defparam i2_3_lut_4_lut_adj_1663.LUT_INIT = 16'h9669;
    SB_LUT4 i62466_4_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_612), 
            .I2(LED_N_3408), .I3(Kp_23__N_1748), .O(n28131));
    defparam i62466_4_lut.LUT_INIT = 16'hc4a0;
    SB_LUT4 i18_4_lut_adj_1664 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_5104));   // verilog/coms.v(157[7:23])
    defparam i18_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 select_787_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4905));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4904));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16_4_lut_adj_1665 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_5105));   // verilog/coms.v(157[7:23])
    defparam i16_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1666 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_5106));   // verilog/coms.v(157[7:23])
    defparam i17_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1667 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_5107));   // verilog/coms.v(157[7:23])
    defparam i15_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1668 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_5108));   // verilog/coms.v(157[7:23])
    defparam i14_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(157[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41_adj_5107), .I1(n43_adj_5106), .I2(n42_adj_5105), 
            .I3(n44_adj_5104), .O(n50));   // verilog/coms.v(157[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1669 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45_adj_5109));   // verilog/coms.v(157[7:23])
    defparam i19_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45_adj_5109), .I1(n50), .I2(n39), .I3(n40_adj_5108), 
            .O(n25879));   // verilog/coms.v(157[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30733_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25879), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i30733_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i468_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2068));   // verilog/coms.v(148[4] 304[11])
    defparam i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [3]), 
            .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4903));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4902));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4901));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4900));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4899));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1671 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [6]), 
            .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4898));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1671.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4897));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4896));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1672 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [3]), 
            .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4895));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1672.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4894));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4893));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4892));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [7]), 
            .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4891));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4890));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4889));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(\control_mode[6] ), .I1(\control_mode[5] ), 
            .I2(control_mode_c[4]), .I3(\control_mode[7] ), .O(n71502));
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1676 (.I0(n71502), .I1(control_mode[2]), .I2(control_mode[3]), 
            .I3(GND_net), .O(n53108));
    defparam i1_3_lut_adj_1676.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1677 (.I0(n53108), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n23));
    defparam i1_2_lut_adj_1677.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1678 (.I0(n27258), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[16] [7]), .I3(\data_out_frame[19] [2]), 
            .O(n67139));
    defparam i1_2_lut_3_lut_4_lut_adj_1678.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1679 (.I0(n53108), .I1(control_mode[1]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15_adj_7));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1679.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1680 (.I0(n53108), .I1(control_mode[1]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1680.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1681 (.I0(n10_adj_5089), .I1(n67716), .I2(n8_adj_5078), 
            .I3(GND_net), .O(n28674));
    defparam i1_2_lut_3_lut_adj_1681.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1682 (.I0(n10_adj_5089), .I1(n67716), .I2(n8_adj_11), 
            .I3(GND_net), .O(n28676));
    defparam i1_2_lut_3_lut_adj_1682.LUT_INIT = 16'hfbfb;
    SB_LUT4 i14517_3_lut_4_lut (.I0(n10_adj_5089), .I1(n67716), .I2(reset), 
            .I3(n8_adj_10), .O(n28730));
    defparam i14517_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_3_lut_4_lut_adj_1683 (.I0(\data_out_frame[23] [5]), .I1(n67291), 
            .I2(\data_out_frame[24] [0]), .I3(n62273), .O(n67557));
    defparam i2_3_lut_4_lut_adj_1683.LUT_INIT = 16'h9669;
    SB_LUT4 i39074_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n23094), .I3(GND_net), .O(n29942));
    defparam i39074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\current[15] ), 
            .I2(\data_out_frame[21] [7]), .I3(\FRAME_MATCHER.i_31__N_2509 ), 
            .O(n2_adj_4922));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hd800;
    SB_LUT4 i1_4_lut_4_lut_adj_1684 (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I1(\current[15] ), .I2(\data_out_frame[21] [5]), .I3(\FRAME_MATCHER.i_31__N_2509 ), 
            .O(n2_adj_4913));
    defparam i1_4_lut_4_lut_adj_1684.LUT_INIT = 16'hd800;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [3]), 
            .I2(encoder0_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4797));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4950));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i5_3_lut_4_lut_adj_1686 (.I0(\data_in_frame[4] [5]), .I1(n26323), 
            .I2(n26197), .I3(\data_in_frame[8] [1]), .O(n14_adj_5096));
    defparam i5_3_lut_4_lut_adj_1686.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1687 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[4] [2]), .I3(n67070), .O(n67563));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1687.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1688 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [7]), 
            .I2(n61447), .I3(GND_net), .O(n6_adj_5034));
    defparam i2_2_lut_3_lut_adj_1688.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1689 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[17] [2]), 
            .I2(n67429), .I3(GND_net), .O(n6_adj_5033));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1689.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1690 (.I0(\data_out_frame[21] [2]), .I1(n27164), 
            .I2(n61577), .I3(\data_out_frame[23] [4]), .O(n62268));
    defparam i2_3_lut_4_lut_adj_1690.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1691 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(n66964), .I3(GND_net), .O(n71706));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1691.LUT_INIT = 16'h9696;
    SB_LUT4 i59848_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n45283), 
            .I2(n89), .I3(n3476), .O(n75250));
    defparam i59848_2_lut_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1692 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(\data_in_frame[1][3] ), .I3(\data_in_frame[1][5] ), .O(n67338));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1692.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1693 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(n67563), .I3(\data_in_frame[1][5] ), .O(n44_adj_5085));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1693.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1694 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[4] [2]), .O(n67185));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut_adj_1694.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1695 (.I0(\data_in_frame[1] [4]), .I1(n67142), 
            .I2(n62400), .I3(n67198), .O(n69356));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut_adj_1695.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1696 (.I0(\data_in_frame[1] [4]), .I1(n67142), 
            .I2(n67352), .I3(n66918), .O(n26317));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1696.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1697 (.I0(n26724), .I1(n67441), .I2(\data_in_frame[6] [5]), 
            .I3(n67099), .O(Kp_23__N_974));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_4_lut_adj_1697.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1698 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[6] [1]), .O(n67352));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1698.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1699 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[4] [0]), 
            .I2(n69802), .I3(n67182), .O(n35_adj_5086));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1699.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1700 (.I0(\data_in_frame[13][7] ), .I1(\data_in_frame[13][6] ), 
            .I2(\data_in_frame[16] [2]), .I3(GND_net), .O(n7_adj_5079));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_3_lut_adj_1700.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1701 (.I0(\data_in_frame[13][7] ), .I1(\data_in_frame[13][6] ), 
            .I2(n62034), .I3(GND_net), .O(n62266));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1701.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63576 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n79456));
    defparam byte_transmit_counter_0__bdd_4_lut_63576.LUT_INIT = 16'he4aa;
    SB_LUT4 i15574_3_lut_4_lut (.I0(n28658), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n29788));
    defparam i15574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16234_3_lut (.I0(\data_in_frame[16]_c [6]), .I1(rx_data[6]), 
            .I2(n28717), .I3(GND_net), .O(n30448));   // verilog/coms.v(130[12] 305[6])
    defparam i16234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16231_3_lut (.I0(\data_in_frame[16]_c [5]), .I1(rx_data[5]), 
            .I2(n28717), .I3(GND_net), .O(n30445));   // verilog/coms.v(130[12] 305[6])
    defparam i16231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1702 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[8] [1]), .I3(GND_net), .O(n67013));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1702.LUT_INIT = 16'h9696;
    SB_LUT4 i15568_3_lut_4_lut (.I0(n28658), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[20][4] ), .O(n29782));
    defparam i15568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1703 (.I0(n62080), .I1(n67271), .I2(n67249), 
            .I3(GND_net), .O(n26592));
    defparam i1_2_lut_3_lut_adj_1703.LUT_INIT = 16'h9696;
    SB_LUT4 i15565_3_lut_4_lut (.I0(n28658), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29779));
    defparam i15565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1704 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n66967), .I3(n35_adj_4953), .O(n27292));
    defparam i1_2_lut_4_lut_adj_1704.LUT_INIT = 16'h6996;
    SB_LUT4 i15693_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[7]), 
            .I3(\data_in_frame[1][7] ), .O(n29907));
    defparam i15693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15558_3_lut_4_lut (.I0(n28658), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[20][2] ), .O(n29772));
    defparam i15558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1705 (.I0(\data_out_frame[12] [1]), .I1(n30), 
            .I2(n10_adj_12), .I3(\data_out_frame[11] [7]), .O(n61517));
    defparam i1_2_lut_4_lut_adj_1705.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n66748));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15689_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[6]), 
            .I3(\data_in_frame[1][6] ), .O(n29903));
    defparam i15689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1706 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[4] [7]), .O(n30));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1706.LUT_INIT = 16'h6996;
    SB_LUT4 i15686_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[5]), 
            .I3(\data_in_frame[1][5] ), .O(n29900));
    defparam i15686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15683_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29897));
    defparam i15683_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15555_3_lut_4_lut (.I0(n28658), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[20][1] ), .O(n29769));
    defparam i15555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15680_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[3]), 
            .I3(\data_in_frame[1][3] ), .O(n29894));
    defparam i15680_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15677_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[2]), 
            .I3(\data_in_frame[1][2] ), .O(n29891));
    defparam i15677_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15674_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[1]), 
            .I3(\data_in_frame[1][1] ), .O(n29888));
    defparam i15674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15671_3_lut_4_lut (.I0(n8_adj_10), .I1(n66860), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29885));
    defparam i15671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1707 (.I0(n67079), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[10] [0]), .I3(\data_in_frame[11] [7]), .O(n67596));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1707.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1708 (.I0(n67079), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[10] [0]), .I3(\data_in_frame[12][2] ), .O(n67243));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1708.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1709 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n66868), .O(n66872));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1709.LUT_INIT = 16'hffdf;
    SB_LUT4 i39075_3_lut (.I0(control_mode_c[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n23094), .I3(GND_net), .O(n29985));
    defparam i39075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1710 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n66860), .O(n66866));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1710.LUT_INIT = 16'hffdf;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63353 (.I0(byte_transmit_counter[1]), 
            .I1(n72605), .I2(n72606), .I3(byte_transmit_counter[2]), .O(n79228));
    defparam byte_transmit_counter_1__bdd_4_lut_63353.LUT_INIT = 16'he4aa;
    SB_LUT4 n79228_bdd_4_lut (.I0(n79228), .I1(n72600), .I2(n72599), .I3(byte_transmit_counter[2]), 
            .O(n79231));
    defparam n79228_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1711 (.I0(n26246), .I1(n26331), .I2(\data_in_frame[10] [6]), 
            .I3(GND_net), .O(n67515));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1711.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63348 (.I0(byte_transmit_counter[1]), 
            .I1(n72569), .I2(n72570), .I3(byte_transmit_counter[2]), .O(n79216));
    defparam byte_transmit_counter_1__bdd_4_lut_63348.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1712 (.I0(n26246), .I1(n26331), .I2(\data_in_frame[8] [7]), 
            .I3(GND_net), .O(n71776));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1712.LUT_INIT = 16'h9696;
    SB_LUT4 n79456_bdd_4_lut (.I0(n79456), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n79459));
    defparam n79456_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1713 (.I0(n27117), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11]_c [4]), .I3(\data_in_frame[9] [3]), .O(n26364));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1713.LUT_INIT = 16'h6996;
    SB_LUT4 i15552_3_lut_4_lut (.I0(n28658), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[20][0] ), .O(n29766));
    defparam i15552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_789_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5028));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[5]), 
            .I3(GND_net), .O(n1_adj_5025));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i5_3_lut_4_lut_adj_1714 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [4]), 
            .I2(n10_adj_4930), .I3(n67527), .O(n67167));   // verilog/coms.v(88[17:63])
    defparam i5_3_lut_4_lut_adj_1714.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1715 (.I0(\data_in_frame[10] [4]), .I1(n67111), 
            .I2(\data_in_frame[12][6] ), .I3(GND_net), .O(n66942));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1715.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(n1_adj_5024));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1716 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n8_adj_4929));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1716.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1717 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [6]), 
            .I2(n67587), .I3(GND_net), .O(n67400));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1717.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5023));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_3_lut_4_lut_adj_1718 (.I0(n26345), .I1(n27_adj_5084), .I2(n26959), 
            .I3(n62327), .O(n24167));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_4_lut_adj_1718.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1719 (.I0(\data_in_frame[10] [7]), .I1(n67419), 
            .I2(\data_in_frame[15][5] ), .I3(n10_adj_5056), .O(n62329));   // verilog/coms.v(88[17:63])
    defparam i5_3_lut_4_lut_adj_1719.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n1_adj_5022));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1720 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[6] [7]), .I3(n1168), .O(n67587));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1720.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1721 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[8] [4]), .O(n66878));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1721.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1722 (.I0(\data_in_frame[10] [7]), .I1(n67419), 
            .I2(n26959), .I3(GND_net), .O(n62327));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1722.LUT_INIT = 16'h9696;
    SB_LUT4 n79216_bdd_4_lut (.I0(n79216), .I1(n72564), .I2(n72563), .I3(byte_transmit_counter[2]), 
            .O(n79219));
    defparam n79216_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_789_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n1_adj_5021));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1723 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [2]), .I3(\data_out_frame[10] [6]), 
            .O(n67527));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1723.LUT_INIT = 16'h6996;
    SB_LUT4 i61955_3_lut (.I0(n79441), .I1(n79237), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n77811));
    defparam i61955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63536 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n79450));
    defparam byte_transmit_counter_0__bdd_4_lut_63536.LUT_INIT = 16'he4aa;
    SB_LUT4 i63185_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n45392), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i63185_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_3_lut_4_lut_adj_1724 (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n45392), .I3(\FRAME_MATCHER.i_31__N_2511 ), .O(n25859));
    defparam i1_3_lut_4_lut_adj_1724.LUT_INIT = 16'hef00;
    SB_LUT4 n79450_bdd_4_lut (.I0(n79450), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n79453));
    defparam n79450_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1725 (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(\FRAME_MATCHER.i_31__N_2511 ), .I3(n45392), .O(n69824));
    defparam i2_3_lut_4_lut_adj_1725.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_1726 (.I0(n6_adj_9), .I1(n69042), .I2(n26760), 
            .I3(\data_in_frame[16]_c [5]), .O(n69522));
    defparam i2_3_lut_4_lut_adj_1726.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1727 (.I0(n6_adj_9), .I1(n69042), .I2(\data_in_frame[16] [4]), 
            .I3(n62473), .O(n26551));
    defparam i2_3_lut_4_lut_adj_1727.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1728 (.I0(reset), .I1(n3476), .I2(GND_net), .I3(GND_net), 
            .O(n66835));
    defparam i1_2_lut_adj_1728.LUT_INIT = 16'hbbbb;
    SB_LUT4 i16171_3_lut (.I0(\data_in_frame[14]_c [3]), .I1(rx_data[3]), 
            .I2(n66869), .I3(GND_net), .O(n30385));   // verilog/coms.v(130[12] 305[6])
    defparam i16171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_4_lut_adj_1729 (.I0(\data_in_frame[16]_c [5]), .I1(\data_in_frame[16] [4]), 
            .I2(n67232), .I3(n26760), .O(n71892));
    defparam i1_3_lut_4_lut_adj_1729.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1_adj_5019));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1730 (.I0(\data_in_frame[16]_c [5]), .I1(\data_in_frame[16] [4]), 
            .I2(n61396), .I3(GND_net), .O(n6_adj_5047));
    defparam i1_2_lut_3_lut_adj_1730.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1731 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n66848));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1731.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut_adj_1732 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1951), .I3(n1954), .O(n25868));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1732.LUT_INIT = 16'h4000;
    SB_LUT4 i30428_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n23025), .I3(GND_net), .O(n29992));
    defparam i30428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5018));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_3_lut_4_lut_adj_1733 (.I0(n25590), .I1(\data_in_frame[16] [3]), 
            .I2(n67341), .I3(n69568), .O(Kp_23__N_1607));
    defparam i1_3_lut_4_lut_adj_1733.LUT_INIT = 16'h9669;
    SB_LUT4 i16164_3_lut (.I0(\data_in_frame[14]_c [1]), .I1(rx_data[1]), 
            .I2(n66869), .I3(GND_net), .O(n30378));   // verilog/coms.v(130[12] 305[6])
    defparam i16164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16112_3_lut_4_lut (.I0(n28672), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n30326));
    defparam i16112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1734 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[11] [3]), .I3(GND_net), .O(n8_adj_4885));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1734.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1735 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n66948));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1735.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4948));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_1087_i2_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19]_c [1]), .O(n4932[1]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i2_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i3_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19][2] ), .O(n4932[2]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i4_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19][3] ), .O(n4932[3]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1736 (.I0(n28674), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[11]_c [2]), .O(n66022));
    defparam i1_4_lut_4_lut_4_lut_adj_1736.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1087_i5_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19][4] ), .O(n4932[4]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i5_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_4_lut_adj_1737 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n26480));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1737.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i6_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19][5] ), .O(n4932[5]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i7_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19][6] ), .O(n4932[6]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i8_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19][7] ), .O(n4932[7]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i8_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63531 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n79444));
    defparam byte_transmit_counter_0__bdd_4_lut_63531.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63339 (.I0(byte_transmit_counter[1]), 
            .I1(n72467), .I2(n72468), .I3(byte_transmit_counter[2]), .O(n79210));
    defparam byte_transmit_counter_1__bdd_4_lut_63339.LUT_INIT = 16'he4aa;
    SB_LUT4 n79210_bdd_4_lut (.I0(n79210), .I1(n72555), .I2(n72554), .I3(byte_transmit_counter[2]), 
            .O(n79213));
    defparam n79210_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1087_i9_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n4932[8]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i10_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n4932[9]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63334 (.I0(byte_transmit_counter[1]), 
            .I1(n72494), .I2(n72495), .I3(byte_transmit_counter[2]), .O(n79204));
    defparam byte_transmit_counter_1__bdd_4_lut_63334.LUT_INIT = 16'he4aa;
    SB_LUT4 n79204_bdd_4_lut (.I0(n79204), .I1(n72552), .I2(n72551), .I3(byte_transmit_counter[2]), 
            .O(n79207));
    defparam n79204_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1087_i11_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n4932[10]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i12_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n4932[11]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63358 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n79198));
    defparam byte_transmit_counter_0__bdd_4_lut_63358.LUT_INIT = 16'he4aa;
    SB_LUT4 n79198_bdd_4_lut (.I0(n79198), .I1(\data_out_frame[21] [3]), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n79201));
    defparam n79198_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1738 (.I0(n62080), .I1(\data_out_frame[11] [5]), 
            .I2(n61164), .I3(n26783), .O(n26943));
    defparam i1_2_lut_4_lut_adj_1738.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4947));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i5_3_lut_4_lut_adj_1739 (.I0(\data_out_frame[7] [0]), .I1(n1168), 
            .I2(n10_adj_4878), .I3(n1130), .O(n26783));
    defparam i5_3_lut_4_lut_adj_1739.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i13_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n4932[12]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i14_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n4932[13]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63329 (.I0(byte_transmit_counter[1]), 
            .I1(n72575), .I2(n72576), .I3(byte_transmit_counter[2]), .O(n79186));
    defparam byte_transmit_counter_1__bdd_4_lut_63329.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1087_i15_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n4932[14]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i15_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i16_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n4932[15]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i16_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i21095_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[1] [0]), 
            .I3(\data_in_frame[17] [0]), .O(n4932[16]));   // verilog/coms.v(130[12] 305[6])
    defparam i21095_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i18_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][1] ), .I3(\data_in_frame[17] [1]), .O(n4932[17]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i18_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i19_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][2] ), .I3(\data_in_frame[17] [2]), .O(n4932[18]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i19_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i20_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][3] ), .I3(\data_in_frame[17] [3]), .O(n4932[19]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i21_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n4932[20]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i16079_3_lut_4_lut (.I0(n28676), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n30293));
    defparam i16079_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n79186_bdd_4_lut (.I0(n79186), .I1(n72525), .I2(n72524), .I3(byte_transmit_counter[2]), 
            .O(n79189));
    defparam n79186_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1087_i22_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][5] ), .I3(\data_in_frame[17] [5]), .O(n4932[21]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i23_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][6] ), .I3(\data_in_frame[17] [6]), .O(n4932[22]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i24_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][7] ), .I3(\data_in_frame[17] [7]), .O(n4932[23]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_1087_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i16410_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [7]), 
            .I3(PWMLimit[23]), .O(n30624));   // verilog/coms.v(130[12] 305[6])
    defparam i16410_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16412_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n30626));   // verilog/coms.v(130[12] 305[6])
    defparam i16412_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n79444_bdd_4_lut (.I0(n79444), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n79447));
    defparam n79444_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16416_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [5]), 
            .I3(PWMLimit[21]), .O(n30630));   // verilog/coms.v(130[12] 305[6])
    defparam i16416_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16417_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n30631));   // verilog/coms.v(130[12] 305[6])
    defparam i16417_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16076_3_lut_4_lut (.I0(n28676), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n30290));
    defparam i16076_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16419_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [3]), 
            .I3(PWMLimit[19]), .O(n30633));   // verilog/coms.v(130[12] 305[6])
    defparam i16419_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16451_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n30665));   // verilog/coms.v(130[12] 305[6])
    defparam i16451_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16465_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n30679));   // verilog/coms.v(130[12] 305[6])
    defparam i16465_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16145_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n66872), .I3(GND_net), .O(n30359));   // verilog/coms.v(130[12] 305[6])
    defparam i16145_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1740 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[12] [0]), .O(n8_adj_4872));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1740.LUT_INIT = 16'h6996;
    SB_LUT4 i16467_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n30681));   // verilog/coms.v(130[12] 305[6])
    defparam i16467_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1741 (.I0(\FRAME_MATCHER.i [4]), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(\FRAME_MATCHER.i [3]), 
            .O(n89));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1741.LUT_INIT = 16'h0008;
    SB_LUT4 i2_3_lut_4_lut_adj_1742 (.I0(n62080), .I1(n67271), .I2(\data_out_frame[18] [6]), 
            .I3(\data_out_frame[18] [7]), .O(n67207));
    defparam i2_3_lut_4_lut_adj_1742.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1743 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(n67229), .I3(GND_net), .O(n67216));
    defparam i1_2_lut_3_lut_adj_1743.LUT_INIT = 16'h9696;
    SB_LUT4 i30573_2_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n44662));
    defparam i30573_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51909_2_lut_3_lut (.I0(n3476), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n67716));
    defparam i51909_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i16485_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n30699));   // verilog/coms.v(130[12] 305[6])
    defparam i16485_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16508_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n30722));   // verilog/coms.v(130[12] 305[6])
    defparam i16508_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63315 (.I0(byte_transmit_counter[1]), 
            .I1(n72581), .I2(n72582), .I3(byte_transmit_counter[2]), .O(n79180));
    defparam byte_transmit_counter_1__bdd_4_lut_63315.LUT_INIT = 16'he4aa;
    SB_LUT4 i16072_3_lut_4_lut (.I0(n28676), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n30286));
    defparam i16072_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n79180_bdd_4_lut (.I0(n79180), .I1(n72456), .I2(n72455), .I3(byte_transmit_counter[2]), 
            .O(n79183));
    defparam n79180_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1744 (.I0(n69502), .I1(\data_out_frame[20] [3]), 
            .I2(n67274), .I3(n25458), .O(n67438));
    defparam i1_2_lut_4_lut_adj_1744.LUT_INIT = 16'h9669;
    SB_LUT4 i16509_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n30723));   // verilog/coms.v(130[12] 305[6])
    defparam i16509_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63310 (.I0(byte_transmit_counter[1]), 
            .I1(n72299), .I2(n72300), .I3(byte_transmit_counter[2]), .O(n79174));
    defparam byte_transmit_counter_1__bdd_4_lut_63310.LUT_INIT = 16'he4aa;
    SB_LUT4 i16511_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n30725));   // verilog/coms.v(130[12] 305[6])
    defparam i16511_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1745 (.I0(n61320), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n67453));
    defparam i1_2_lut_3_lut_adj_1745.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1746 (.I0(n67548), .I1(n10_adj_4870), .I2(\data_out_frame[9] [7]), 
            .I3(\data_out_frame[14] [1]), .O(n4_c));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1746.LUT_INIT = 16'h6996;
    SB_LUT4 i16516_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n30730));   // verilog/coms.v(130[12] 305[6])
    defparam i16516_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1747 (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[16] [1]), 
            .I2(n61445), .I3(GND_net), .O(n67222));
    defparam i1_2_lut_3_lut_adj_1747.LUT_INIT = 16'h9696;
    SB_LUT4 n79174_bdd_4_lut (.I0(n79174), .I1(n72282), .I2(n72281), .I3(byte_transmit_counter[2]), 
            .O(n79177));
    defparam n79174_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i23688_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n30732));   // verilog/coms.v(130[12] 305[6])
    defparam i23688_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16519_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n30733));   // verilog/coms.v(130[12] 305[6])
    defparam i16519_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i20487_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n30736));   // verilog/coms.v(130[12] 305[6])
    defparam i20487_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16523_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n30737));   // verilog/coms.v(130[12] 305[6])
    defparam i16523_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63526 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n79438));
    defparam byte_transmit_counter_0__bdd_4_lut_63526.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_3_lut_adj_1748 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[15] [4]), 
            .I2(n1720), .I3(GND_net), .O(n8_adj_4803));
    defparam i2_2_lut_3_lut_adj_1748.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1749 (.I0(n28674), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[11]_c [5]), .O(n66068));
    defparam i1_4_lut_4_lut_4_lut_adj_1749.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1750 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(\data_out_frame[18] [3]), .I3(\data_out_frame[18] [4]), 
            .O(n26));
    defparam i2_2_lut_4_lut_adj_1750.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_out_frame[14] [4]), .I1(n67332), .I2(\data_out_frame[17] [5]), 
            .I3(n26645), .O(n30_c));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i16138_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n66872), .I3(GND_net), .O(n30352));   // verilog/coms.v(130[12] 305[6])
    defparam i16138_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut_adj_1751 (.I0(\data_out_frame[13] [0]), .I1(n45), 
            .I2(\data_out_frame[17] [4]), .I3(\data_out_frame[15] [2]), 
            .O(n67010));
    defparam i2_3_lut_4_lut_adj_1751.LUT_INIT = 16'h6996;
    SB_LUT4 i23301_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n30766));   // verilog/coms.v(130[12] 305[6])
    defparam i23301_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16554_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n30768));   // verilog/coms.v(130[12] 305[6])
    defparam i16554_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16066_3_lut_4_lut (.I0(n28676), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n30280));
    defparam i16066_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n79438_bdd_4_lut (.I0(n79438), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n79441));
    defparam n79438_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16109_3_lut_4_lut (.I0(n28672), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n30323));
    defparam i16109_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1752 (.I0(\data_out_frame[20] [4]), .I1(n26517), 
            .I2(n67203), .I3(GND_net), .O(n26232));
    defparam i1_2_lut_3_lut_adj_1752.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [2]), 
            .I2(encoder0_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4735));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1754 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66982));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1754.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1755 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [1]), 
            .I2(ID[6]), .I3(ID[1]), .O(n12_adj_5111));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut_adj_1755.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1756 (.I0(ID[7]), .I1(ID[2]), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[0] [2]), .O(n10_adj_5112));   // verilog/coms.v(99[12:25])
    defparam i2_4_lut_adj_1756.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1757 (.I0(\data_in_frame[0] [5]), .I1(ID[3]), .I2(ID[5]), 
            .I3(\data_in_frame[0] [3]), .O(n11));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1757.LUT_INIT = 16'h7bde;
    SB_LUT4 i23384_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n30770));   // verilog/coms.v(130[12] 305[6])
    defparam i23384_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63521 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n79432));
    defparam byte_transmit_counter_0__bdd_4_lut_63521.LUT_INIT = 16'he4aa;
    SB_LUT4 n79432_bdd_4_lut (.I0(n79432), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n79435));
    defparam n79432_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(ID[4]), .I1(\data_in_frame[0] [0]), .I2(\data_in_frame[0] [4]), 
            .I3(ID[0]), .O(n9_adj_5113));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'h7bde;
    SB_LUT4 i16558_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n30772));   // verilog/coms.v(130[12] 305[6])
    defparam i16558_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut_adj_1759 (.I0(n9_adj_5113), .I1(n11), .I2(n10_adj_5112), 
            .I3(n12_adj_5111), .O(n69421));   // verilog/coms.v(99[12:25])
    defparam i7_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1760 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_748), 
            .I2(GND_net), .I3(GND_net), .O(n67025));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1760.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1761 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n67067));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1761.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63324 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(byte_transmit_counter[1]), .O(n79162));
    defparam byte_transmit_counter_0__bdd_4_lut_63324.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1762 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n66998));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1762.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1763 (.I0(n61681), .I1(n67001), .I2(n67453), 
            .I3(\data_out_frame[18] [4]), .O(n67277));
    defparam i1_2_lut_4_lut_adj_1763.LUT_INIT = 16'h6996;
    SB_LUT4 i23406_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n30773));   // verilog/coms.v(130[12] 305[6])
    defparam i23406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1764 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n67129));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1764.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_0__7__I_0_4044_2_lut (.I0(\data_in_frame[0] [7]), 
            .I1(\data_in_frame[0] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_753));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_0__7__I_0_4044_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1765 (.I0(Kp_23__N_753), .I1(n67129), .I2(n66998), 
            .I3(\data_in_frame[0] [5]), .O(Kp_23__N_748));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1765.LUT_INIT = 16'h6996;
    SB_LUT4 i23418_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n30774));   // verilog/coms.v(130[12] 305[6])
    defparam i23418_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1766 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n27048));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1766.LUT_INIT = 16'h9696;
    SB_LUT4 equal_2035_i10_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5114));   // verilog/coms.v(169[9:87])
    defparam equal_2035_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n79162_bdd_4_lut (.I0(n79162), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(byte_transmit_counter[1]), 
            .O(n79165));
    defparam n79162_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15721_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16][0] ), 
            .I3(deadband[0]), .O(n29935));   // verilog/coms.v(130[12] 305[6])
    defparam i15721_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1767 (.I0(n27048), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[0] [6]), .O(n23_adj_5115));
    defparam i6_4_lut_adj_1767.LUT_INIT = 16'h4114;
    SB_LUT4 i5_3_lut_adj_1768 (.I0(n26197), .I1(Kp_23__N_748), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n22_adj_5116));
    defparam i5_3_lut_adj_1768.LUT_INIT = 16'h1414;
    SB_LUT4 i10_4_lut_adj_1769 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1][3] ), 
            .I2(\data_in_frame[1][2] ), .I3(\data_in_frame[1][6] ), .O(n27_adj_5117));
    defparam i10_4_lut_adj_1769.LUT_INIT = 16'h8000;
    SB_LUT4 i15724_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13][0] ), 
            .I3(IntegralLimit[0]), .O(n29938));   // verilog/coms.v(130[12] 305[6])
    defparam i15724_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1770 (.I0(current_limit[14]), .I1(\current_limit[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n71866));   // verilog/TinyFPGA_B.v(251[22:35])
    defparam i1_2_lut_adj_1770.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_63305 (.I0(byte_transmit_counter[1]), 
            .I1(n72275), .I2(n72276), .I3(byte_transmit_counter[2]), .O(n79156));
    defparam byte_transmit_counter_1__bdd_4_lut_63305.LUT_INIT = 16'he4aa;
    SB_LUT4 n79156_bdd_4_lut (.I0(n79156), .I1(n72603), .I2(n72602), .I3(byte_transmit_counter[2]), 
            .O(n79159));
    defparam n79156_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(n72550), .I2(n72529), .I3(byte_transmit_counter_c[3]), 
            .O(n79144));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n79144_bdd_4_lut (.I0(n79144), .I1(n72450), .I2(n72449), .I3(byte_transmit_counter_c[3]), 
            .O(n79147));
    defparam n79144_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63296 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(byte_transmit_counter[1]), .O(n79138));
    defparam byte_transmit_counter_0__bdd_4_lut_63296.LUT_INIT = 16'he4aa;
    SB_LUT4 n79138_bdd_4_lut (.I0(n79138), .I1(\data_out_frame[21] [0]), 
            .I2(\data_out_frame[20] [0]), .I3(byte_transmit_counter[1]), 
            .O(n79141));
    defparam n79138_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1771 (.I0(\data_in_frame[2] [0]), .I1(n10_adj_5114), 
            .I2(n67025), .I3(\data_in_frame[1][5] ), .O(n26_adj_5118));
    defparam i9_4_lut_adj_1771.LUT_INIT = 16'h2100;
    SB_LUT4 i15725_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [0]), 
            .I3(\Kp[0] ), .O(n29939));   // verilog/coms.v(130[12] 305[6])
    defparam i15725_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63278 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(byte_transmit_counter[1]), .O(n79132));
    defparam byte_transmit_counter_0__bdd_4_lut_63278.LUT_INIT = 16'he4aa;
    SB_LUT4 n79132_bdd_4_lut (.I0(n79132), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(byte_transmit_counter[1]), 
            .O(n79135));
    defparam n79132_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15726_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n29940));   // verilog/coms.v(130[12] 305[6])
    defparam i15726_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(current_limit[15]), .I1(n71866), .I2(n65), 
            .I3(current_limit[13]), .O(n51));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'h5554;
    SB_LUT4 i12_4_lut_adj_1773 (.I0(n23_adj_5115), .I1(\data_in_frame[1][7] ), 
            .I2(n26190), .I3(n67025), .O(n29));
    defparam i12_4_lut_adj_1773.LUT_INIT = 16'h0208;
    SB_LUT4 i65_3_lut (.I0(n22), .I1(\current[11] ), .I2(current_limit[11]), 
            .I3(GND_net), .O(n65));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i65_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i14_4_lut_adj_1774 (.I0(n27_adj_5117), .I1(n69421), .I2(n22_adj_5116), 
            .I3(n26752), .O(n31));
    defparam i14_4_lut_adj_1774.LUT_INIT = 16'h0020;
    SB_LUT4 i59626_4_lut (.I0(current_limit[14]), .I1(n65), .I2(current_limit[13]), 
            .I3(\current_limit[12] ), .O(n75118));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i59626_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i23436_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n29944));   // verilog/coms.v(130[12] 305[6])
    defparam i23436_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23502_4_lut (.I0(n51), .I1(n75118), .I2(\current[15] ), .I3(current_limit[15]), 
            .O(n260));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i23502_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i16059_3_lut_4_lut (.I0(n28676), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n30273));
    defparam i16059_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1775 (.I0(n31), .I1(n29), .I2(n72045), .I3(n26_adj_5118), 
            .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut_adj_1775.LUT_INIT = 16'h0800;
    SB_LUT4 i15806_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n30020));   // verilog/coms.v(130[12] 305[6])
    defparam i15806_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15807_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n30021));   // verilog/coms.v(130[12] 305[6])
    defparam i15807_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15808_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n30022));   // verilog/coms.v(130[12] 305[6])
    defparam i15808_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16056_3_lut_4_lut (.I0(n28676), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n30270));
    defparam i16056_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_214_i3_3_lut_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\data_out_frame[24] [4]), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(n67438), .O(n3_adj_5016));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_214_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i2_2_lut_4_lut_adj_1776 (.I0(\data_out_frame[23] [5]), .I1(n67291), 
            .I2(\data_out_frame[25] [0]), .I3(\data_out_frame[24] [5]), 
            .O(n6_adj_4756));
    defparam i2_2_lut_4_lut_adj_1776.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [1]), 
            .I2(encoder0_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4734));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'ha088;
    SB_LUT4 i15809_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n30023));   // verilog/coms.v(130[12] 305[6])
    defparam i15809_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_3_lut_adj_1778 (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(\FRAME_MATCHER.i_31__N_2512 ), .I3(GND_net), .O(n6_adj_4746));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_3_lut_adj_1778.LUT_INIT = 16'hfefe;
    SB_LUT4 i14987_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n29201));   // verilog/coms.v(130[12] 305[6])
    defparam i14987_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15810_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n30024));   // verilog/coms.v(130[12] 305[6])
    defparam i15810_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14981_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n29195));   // verilog/coms.v(130[12] 305[6])
    defparam i14981_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15811_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n30025));   // verilog/coms.v(130[12] 305[6])
    defparam i15811_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15812_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n30026));   // verilog/coms.v(130[12] 305[6])
    defparam i15812_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15813_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n30027));   // verilog/coms.v(130[12] 305[6])
    defparam i15813_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1779 (.I0(\data_out_frame[22] [4]), .I1(n24023), 
            .I2(\data_out_frame[24] [6]), .I3(n26232), .O(n67432));
    defparam i2_3_lut_4_lut_adj_1779.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_3_lut (.I0(LED_N_3408), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(reset), .I3(GND_net), .O(n23025));   // verilog/coms.v(130[12] 305[6])
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i15814_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n30028));   // verilog/coms.v(130[12] 305[6])
    defparam i15814_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15815_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n30029));   // verilog/coms.v(130[12] 305[6])
    defparam i15815_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15816_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n30030));   // verilog/coms.v(130[12] 305[6])
    defparam i15816_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_3_lut_4_lut_adj_1780 (.I0(\data_out_frame[23] [0]), .I1(n61954), 
            .I2(n10_adj_4741), .I3(\data_out_frame[24] [7]), .O(n61789));
    defparam i5_3_lut_4_lut_adj_1780.LUT_INIT = 16'h6996;
    SB_LUT4 i15817_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n30031));   // verilog/coms.v(130[12] 305[6])
    defparam i15817_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15818_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n30032));   // verilog/coms.v(130[12] 305[6])
    defparam i15818_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_3_lut_adj_1781 (.I0(\data_out_frame[25] [4]), .I1(n61412), 
            .I2(n62268), .I3(GND_net), .O(n6_c));
    defparam i2_2_lut_3_lut_adj_1781.LUT_INIT = 16'h6969;
    SB_LUT4 i15819_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n30033));   // verilog/coms.v(130[12] 305[6])
    defparam i15819_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15820_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n30034));   // verilog/coms.v(130[12] 305[6])
    defparam i15820_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15821_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n30035));   // verilog/coms.v(130[12] 305[6])
    defparam i15821_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [0]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n16_c));
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15822_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n30036));   // verilog/coms.v(130[12] 305[6])
    defparam i15822_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i20913_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[13] ), .O(n30037));   // verilog/coms.v(130[12] 305[6])
    defparam i20913_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_3_lut_adj_1782 (.I0(n61681), .I1(n26517), .I2(n27164), 
            .I3(GND_net), .O(n10_c));
    defparam i2_2_lut_3_lut_adj_1782.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1783 (.I0(n67161), .I1(\data_out_frame[24] [6]), 
            .I2(n26232), .I3(\data_out_frame[25] [0]), .O(n6_adj_4739));
    defparam i2_2_lut_4_lut_adj_1783.LUT_INIT = 16'h6996;
    SB_LUT4 i15824_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[12] ), .O(n30038));   // verilog/coms.v(130[12] 305[6])
    defparam i15824_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15825_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[11] ), .O(n30039));   // verilog/coms.v(130[12] 305[6])
    defparam i15825_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_221_i3_3_lut_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(n61412), .I2(\FRAME_MATCHER.state[3] ), .I3(n62476), .O(n3_adj_5017));
    defparam select_787_Select_221_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i1_2_lut_4_lut_adj_1784 (.I0(\data_out_frame[25] [3]), .I1(n21), 
            .I2(n19), .I3(n20_adj_4742), .O(n62476));
    defparam i1_2_lut_4_lut_adj_1784.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63273 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter[1]), .O(n79108));
    defparam byte_transmit_counter_0__bdd_4_lut_63273.LUT_INIT = 16'he4aa;
    SB_LUT4 i20938_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[10] ), .O(n30040));   // verilog/coms.v(130[12] 305[6])
    defparam i20938_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n79108_bdd_4_lut (.I0(n79108), .I1(\data_out_frame[21] [2]), 
            .I2(\data_out_frame[20] [2]), .I3(byte_transmit_counter[1]), 
            .O(n79111));
    defparam n79108_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15827_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[9] ), .O(n30041));   // verilog/coms.v(130[12] 305[6])
    defparam i15827_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15828_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[8] ), .O(n30042));   // verilog/coms.v(130[12] 305[6])
    defparam i15828_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15829_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [7]), 
            .I3(\Kp[7] ), .O(n30043));   // verilog/coms.v(130[12] 305[6])
    defparam i15829_3_lut_4_lut.LUT_INIT = 16'hf780;
    uart_tx tx (.clk16MHz(clk16MHz), .tx_o(tx_o), .tx_data({tx_data}), 
            .r_SM_Main({r_SM_Main}), .GND_net(GND_net), .n29956(n29956), 
            .tx_active(tx_active), .r_Clock_Count({r_Clock_Count}), .VCC_net(VCC_net), 
            .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n5220(n5220), .n29(n29_adj_5120), .n23(n23_adj_5121), .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), 
            .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), .n27(n27_adj_13), 
            .n67730(n67730), .n68353(n68353), .n6(n6_adj_14), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.GND_net(GND_net), .r_Clock_Count({r_Clock_Count_adj_26}), 
            .VCC_net(VCC_net), .baudrate({baudrate}), .n28240(n28240), 
            .clk16MHz(clk16MHz), .n67800(n67800), .\r_SM_Main[2] (\r_SM_Main[2]_adj_23 ), 
            .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), 
            .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), .n5217(n5217), .n66790(n66790), 
            .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), .n29(n29_adj_5120), 
            .n23(n23_adj_5121), .\r_SM_Main[1] (\r_SM_Main[1]_adj_24 ), 
            .n27(n27_adj_13), .n28117(n28117), .n70292(n70292), .n29937(n29937), 
            .rx_data({rx_data}), .n29936(n29936), .n29934(n29934), .n29915(n29915), 
            .n29914(n29914), .n29910(n29910), .n29906(n29906), .n30762(n30762), 
            .n62510(n62510), .rx_data_ready(rx_data_ready), .n30758(n30758), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n70662(n70662), .n34(n34_adj_25), 
            .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), 
            .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), 
            .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), 
            .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), 
            .n70340(n70340), .n5220(n5220), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
            .n70356(n70356), .n70276(n70276), .n70324(n70324), .n70308(n70308), 
            .n70388(n70388), .n70372(n70372), .\r_SM_Main[0] (r_SM_Main[0]), 
            .n68353(n68353)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk16MHz, tx_o, tx_data, r_SM_Main, GND_net, n29956, 
            tx_active, r_Clock_Count, VCC_net, \r_SM_Main_2__N_3536[1] , 
            \r_SM_Main_2__N_3545[0] , n5220, n29, n23, \o_Rx_DV_N_3488[12] , 
            \o_Rx_DV_N_3488[24] , n27, n67730, n68353, n6, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output tx_o;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    input GND_net;
    input n29956;
    output tx_active;
    output [8:0]r_Clock_Count;
    input VCC_net;
    input \r_SM_Main_2__N_3536[1] ;
    input \r_SM_Main_2__N_3545[0] ;
    input n5220;
    input n29;
    input n23;
    input \o_Rx_DV_N_3488[12] ;
    input \o_Rx_DV_N_3488[24] ;
    input n27;
    input n67730;
    input n68353;
    output n6;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n460;
    
    wire n67828;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n29498, n3, n40346, n25370;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n62542, n75129, n67611, n62540, n72293, n72294, n72297, 
        n72296, n79648;
    wire [8:0]n41;
    
    wire n40318, n3_adj_4733, n60328, n60327, n60326, n60325, n60324, 
        n60323, n60322, n60321, n70220, n70226, n66774, n75111, 
        n75108, n9, n79171, n14, n15, n79168;
    
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n67828), 
            .D(n460[1]), .R(n29498));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n67828), 
            .D(n460[2]), .R(n29498));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n40346), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n62542), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i12_4_lut (.I0(n75129), .I1(n67828), .I2(r_Bit_Index[0]), 
            .I3(n67611), .O(n62540));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i56437_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n72293));
    defparam i56437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56438_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n72294));
    defparam i56438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56441_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n72297));
    defparam i56441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56440_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n72296));
    defparam i56440_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n79648));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n29956));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Clock_Count_2056__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n40346), .D(n41[0]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n40346), .D(n41[1]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n40346), .D(n41[2]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n40346), .D(n41[3]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n40346), .D(n41[4]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n40346), .D(n41[5]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n40346), .D(n41[6]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n40346), .D(n41[7]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n40346), .D(n41[8]), .R(n40318));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n62540));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_4733), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n25370), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i63234_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n67828));
    defparam i63234_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n25370));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 r_Clock_Count_2056_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n60328), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2056_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n60327), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_9 (.CI(n60327), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n60328));
    SB_LUT4 r_Clock_Count_2056_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n60326), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_8 (.CI(n60326), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n60327));
    SB_LUT4 r_Clock_Count_2056_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n60325), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_7 (.CI(n60325), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n60326));
    SB_LUT4 r_Clock_Count_2056_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n60324), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_6 (.CI(n60324), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n60325));
    SB_LUT4 r_Clock_Count_2056_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n60323), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_5 (.CI(n60323), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n60324));
    SB_LUT4 r_Clock_Count_2056_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n60322), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_4 (.CI(n60322), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n60323));
    SB_LUT4 r_Clock_Count_2056_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n60321), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_3 (.CI(n60321), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n60322));
    SB_LUT4 r_Clock_Count_2056_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n60321));
    SB_LUT4 i1_2_lut (.I0(n5220), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n70220));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), .I3(n70220), 
            .O(n70226));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i10_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(r_SM_Main[1]), .I2(n27), 
            .I3(n70226), .O(n3_adj_4733));   // verilog/uart_tx.v(32[16:25])
    defparam i10_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i63182_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n40318));
    defparam i63182_4_lut.LUT_INIT = 16'h1113;
    SB_LUT4 i60370_3_lut (.I0(n66774), .I1(\o_Rx_DV_N_3488[12] ), .I2(n5220), 
            .I3(GND_net), .O(n75111));   // verilog/uart_tx.v(32[16:25])
    defparam i60370_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i60366_4_lut (.I0(n75111), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n75108));   // verilog/uart_tx.v(32[16:25])
    defparam i60366_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i23_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n75108), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n9));   // verilog/uart_tx.v(32[16:25])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_3_lut (.I0(n9), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n62542));   // verilog/uart_tx.v(32[16:25])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40346));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(n79171), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i26200_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(34[16:27])
    defparam i26200_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n66774));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i51811_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n67611));
    defparam i51811_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1077 (.I0(n67730), .I1(n67611), .I2(r_SM_Main[1]), 
            .I3(n66774), .O(n29498));
    defparam i1_4_lut_adj_1077.LUT_INIT = 16'h1101;
    SB_LUT4 i16_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n68353), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5220), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n40346), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n79648));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i60412_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n75129));   // verilog/uart_tx.v(32[16:25])
    defparam i60412_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(n72296), 
            .I2(n72297), .I3(r_Bit_Index[1]), .O(n79168));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n79168_bdd_4_lut (.I0(n79168), .I1(n72294), .I2(n72293), .I3(r_Bit_Index[1]), 
            .O(n79171));
    defparam n79168_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, r_Clock_Count, VCC_net, baudrate, n28240, 
            clk16MHz, n67800, \r_SM_Main[2] , r_Rx_Data, RX_N_2, \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[12] , n5217, n66790, \o_Rx_DV_N_3488[24] , 
            n29, n23, \r_SM_Main[1] , n27, n28117, n70292, n29937, 
            rx_data, n29936, n29934, n29915, n29914, n29910, n29906, 
            n30762, n62510, rx_data_ready, n30758, \r_Bit_Index[0] , 
            n70662, n34, \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , n70340, n5220, 
            \r_SM_Main_2__N_3536[1] , n70356, n70276, n70324, n70308, 
            n70388, n70372, \r_SM_Main[0] , n68353) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [7:0]r_Clock_Count;
    input VCC_net;
    input [31:0]baudrate;
    output n28240;
    input clk16MHz;
    output n67800;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[12] ;
    input n5217;
    input n66790;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    output \r_SM_Main[1] ;
    output n27;
    output n28117;
    output n70292;
    input n29937;
    output [7:0]rx_data;
    input n29936;
    input n29934;
    input n29915;
    input n29914;
    input n29910;
    input n29906;
    input n30762;
    input n62510;
    output rx_data_ready;
    input n30758;
    output \r_Bit_Index[0] ;
    output n70662;
    output n34;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n70340;
    input n5220;
    output \r_SM_Main_2__N_3536[1] ;
    output n70356;
    output n70276;
    output n70324;
    output n70308;
    output n70388;
    output n70372;
    input \r_SM_Main[0] ;
    output n68353;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]n1;
    
    wire n60285, n60286, n60284, n60283, n1742, n3060;
    wire [23:0]n8683;
    wire [23:0]n294;
    
    wire n3165, n1879, n3059, n3164, n2013, n3058, n3163, n2144, 
        n3057, n3162, n2272, n3056, n3161, n2397, n3055, n3160;
    wire [2:0]n479;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n2519, n3054, n3159, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire r_Rx_Data_R, n75177, n75174, n70280, n70286, n2638, n3053, 
        n3158, n2754, n3052, n3157, n2867, n3051, n3156, n2977, 
        n3050, n3155, n3084, n3049, n3154, n3188, n3048, n3153, 
        n3082, n3047, n3152, n2951;
    wire [23:0]n8657;
    
    wire n2939, n2940, n2941, n2944, n35, n2942, n39, n2945, 
        n33, n2943, n37, n2947, n2948, n27_adj_4455, n29_adj_4456, 
        n2949, n2950, n23_adj_4457, n25, n2956, n3064, n2957, 
        n3065, n11, n2952, n2946, n2954, n3062, n2953, n3061, 
        n15, n17, n19, n31, n2955, n3063, n13, n21, n75913, 
        n76885, n77381, n72184, n77377, n75917, n72228, n72230, 
        n3066, n8, n77581, n77582, n16, n34_c, n78173, n1831, 
        n70074, n1977, n75906, n14, n75902, n77870, n76641, n10, 
        n77583, n77584, n75928, n76865, n12, n20, n76639, n77761, 
        n78233, n77670, n72232, n78259, n78260, n77884, n77885, 
        n2829;
    wire [23:0]n8631;
    
    wire n2828, n77243, n1408, n72242, n2832, n37_adj_4458, n2830, 
        n41, n2833, n35_adj_4459, n2831, n39_adj_4460, n2835, n2836, 
        n29_adj_4461, n31_adj_4462, n2837, n2839, n2838, n23_adj_4463, 
        n25_adj_4464, n27_adj_4465, n70072, n1560, n2843, n2844, 
        n2845, n13_adj_4466, n15_adj_4467, n2840, n2834, n2713;
    wire [23:0]n8605;
    
    wire n2827, n2714, n2717, n39_adj_4468, n2718, n37_adj_4469, 
        n2715, n43_adj_4470, n2716, n41_adj_4471, n2722, n2724, 
        n2723, n25_adj_4472, n27_adj_4473, n29_adj_4474, n2728, n2842, 
        n2729, n2730, n71350;
    wire [23:0]n8371;
    
    wire n48, n1702, n15_adj_4475, n17_adj_4476, n2720, n2721, n31_adj_4477, 
        n33_adj_4478, n2719, n35_adj_4479, n2601;
    wire [23:0]n8579;
    
    wire n2596, n2599, n41_adj_4480, n2597, n45_adj_4481, n2600, 
        n39_adj_4482, n79649, n2598, n43_adj_4483, n2604, n2606, 
        n2605, n27_adj_4484, n29_adj_4485, n31_adj_4486, n2602, n2603, 
        n33_adj_4487, n35_adj_4488, n2610, n2727, n2611, n2612, 
        n17_adj_4489, n19_adj_4490, n1413, n1414, n75472, n2607, 
        n2726, n21_adj_4491, n2725, n23_adj_4492, n25_adj_4493, n37_adj_4494, 
        n28161, n29423, n76092, n77037, n77459, n77457, n76094, 
        n14_adj_4497, n77601, n77602, n22, n40_adj_4498, n76082, 
        n20_adj_4499, n76078, n77664, n36, n76617, n18, n26, n16_adj_4500, 
        n76108, n78093, n78094, n77873, n77795, n78105;
    wire [23:0]n8709;
    
    wire n3151, n3186, n60147, n60146, n60145, n76615, n78107, 
        n2608, n60144, n60143, n60142, n2476;
    wire [23:0]n8553;
    
    wire n2477, n60141, n60140, n2481, n60139, n60138, n37_adj_4501, 
        n60137, n2478, n60136, n60135, n60134, n43_adj_4502, n2479, 
        n60133, n67928, n3166, n1602, n60132, n3167, n1459, n60131, 
        n41_adj_4503, n2480, n3168, n1460, n60130, n3169, n1011, 
        n60129, n3170, n856, n60128, n39_adj_4504, n3171, n698, 
        n60127, n3172, n858, n60126, n70092, n538, n60125, n67874, 
        n2486, n2485, n27_adj_4505, n29_adj_4506, n3046, n60124, 
        n72246, n60123, n2491, n60122, n60121, n2482, n2483, n48_adj_4507, 
        n2484, n60120, n31_adj_4508, n33_adj_4509, n60119, n35_adj_4510, 
        n60118, n60117, n41_adj_4511, n39_adj_4512, n2490, n29_adj_4513, 
        n19_adj_4514, n31_adj_4515, n37_adj_4516, n23_adj_4517, n25_adj_4518, 
        n7, n45_adj_4519, n9, n2609, n21_adj_4520, n17_adj_4521, 
        n2353;
    wire [23:0]n8527;
    
    wire n60116, n2363, n2357, n21_adj_4522, n19_adj_4523, n43_adj_4524, 
        n33_adj_4525, n39_adj_4526, n35_adj_4527, n11_adj_4528, n13_adj_4529, 
        n15_adj_4530, n27_adj_4531, n2354, n75819, n60115, n45_adj_4532, 
        n60114, n2355, n12_adj_4533, n75811, n10_adj_4534, n60113, 
        n43_adj_4535, n30, n60112, n60111, n60110, n2356, n60109, 
        n75827, n16_adj_4536, n41_adj_4537, n60108, n75799, n2358, 
        n60107, n60106, n8_adj_4538, n2360, n24, n60105, n3274, 
        n75837, n60104, n76789, n70090, n67878, n2938, n60103, 
        n76783, n60102, n2359, n77956, n33_adj_4539, n60101, n35_adj_4540, 
        n37_adj_4541, n77319, n78120, n60100, n6, n60099, n60098, 
        n77545, n60097, n77546, n48_adj_4542, n4, n60096, n2361, 
        n77543, n60095, n60094, n60093, n2362, n77544, n75813, 
        n78004, n60092, n1265, n38_adj_4543, n1266, n75495, n72256, 
        n76666, n78211, n78212, n78144, n60091, n60090, n60089, 
        n75801, n60088, n77678, n29_adj_4544, n60087, n76664, n75803, 
        n31_adj_4545, n78108, n60086, n70554, n2365, n2488, n76672, 
        n2366, n2489, n3253, n60085, n21_adj_4546, n23_adj_4547, 
        n78110, n2227;
    wire [23:0]n8501;
    
    wire n60084, n2228, n70088, n67882, n70018, n69091, n60083, 
        n60082, n60081, n3_adj_4548, n33_adj_4549, n31_adj_4550, n60080, 
        n60079, n37_adj_4551, n35_adj_4552, n21_adj_4553, n23_adj_4554, 
        n25_adj_4555, n27_adj_4556, n9_adj_4557, n72260, n11_adj_4558, 
        n19_adj_4559, n2229, n2230, n60078, n13_adj_4560, n15_adj_4561, 
        n17_adj_4562, n60077, n29_adj_4563, n60076, n41_adj_4564, 
        n75866, n76835, n77355, n77353, n75868, n6_adj_4565, n77573, 
        n2232, n60075, n37_adj_4566, n60074, n14_adj_4567, n32, 
        n60073, n77574, n75855, n12_adj_4568, n75853, n77982, n76652, 
        n8_adj_4569, n77674, n77675, n75876, n76821, n10_adj_4570, 
        n77676, n76650, n77755, n78207, n60072, n77835, n2231, 
        n78271, n78272, n78264, n60071, n78036, n78037, n60070, 
        n2841, n60069, n39_adj_4571, n2233, n35_adj_4572, n60068, 
        n60067, n60066, n2234, n60065, n2236, n2235, n70086, n67886, 
        n29_adj_4573, n31_adj_4574, n33_adj_4575, n2237, n60064, n60063, 
        n60062, n71354, n60061, n60060, n60059, n71352, n70588, 
        n71474, n71468, n71470, n60058, n60057, n2239, n60056, 
        n2238, n2364, n71472, n9_adj_4576, n14_adj_4577, n71480, 
        n60055, n71478, n26019, n44852, n60054, n42_adj_4578, n21181, 
        n68370, n70654, n28, n60053, n60052, n60051, n60050, n60049, 
        n60048, n60047, n23_adj_4580, n70084, n67890, n77656, n1111, 
        n25_adj_4581, n60046, n27_adj_4582, n2098;
    wire [23:0]n8475;
    
    wire n60045, n60044, n2099, n72264, n60043, n67932, n60042, 
        n60041, n1968;
    wire [23:0]n8449;
    
    wire n2100, n43_adj_4583, n60040, n60039, n2101, n4_adj_4584, 
        n41_adj_4585, n2102, n39_adj_4586, n60038, n2103, n37_adj_4587, 
        n60037, n60036, n60035, n60034, n60033, n60032, n60031, 
        n2104, n60030, n2106, n2105, n31_adj_4588, n70082, n67894, 
        n67924, n60029, n33_adj_4589, n35_adj_4590, n60028, n2107, 
        n60027, n60026, n60025, n60024, n60023, n2108, n2109, 
        n60022, n60021, n60020, n25_adj_4591, n27_adj_4592, n60019, 
        n2487, n60018, n70068, n1267, n60017, n60016, n60015, 
        n60014, n70080, n67898, n1114, n40_adj_4593, n29_adj_4594, 
        n60013, n60012, n1966, n60011, n60010, n60009, n60008, 
        n1967, n60007, n59030, n60006, n60005, n67906, n59029, 
        n70030, n1971, n1972, n59028, n70132, n60004, n35_adj_4595, 
        n60003, n60002, n60001, n60000, n2367, n59999, n70078, 
        n67902, n59998, n37_adj_4596, n59997, n59996, n1969, n41_adj_4597, 
        n59995, n1970, n59994, n59993, n59992, n1115, n75510, 
        n59991, n59027;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n59990, n59989, n59988, n39_adj_4598, n59026, n70130, n59987, 
        n59986, n2240, n59985, n1973, n70076, n59984, n59025, 
        n70128, n59983, n59982, n59981, n59980, n59979, n42_adj_4599, 
        n21191, n68354, n59978, n59024, n59023, n70126, n59977, 
        n1975, n59976, n59975, n59974, n1974, n59973, n59022, 
        n70124, n2110, n29_adj_4600, n31_adj_4601, n33_adj_4602, n59972, 
        n59971, n59021, n70028;
    wire [23:0]n8423;
    
    wire n59970, n59969, n59968, n59967, n59966, n59020, n70122, 
        n59965, n59964, n59963, n1976, n59962, n1832, n1833, n59019, 
        n59961, n59960, n59959, n59018, n59958, n1834, n59957, 
        n1835, n59956, n1836, n59955, n1837, n59954, n1838, n59953, 
        n1558, n1559, n75463, n1839, n59952, n1840, n59951, n41_adj_4603, 
        n1841, n59950, n67915;
    wire [23:0]n8397;
    
    wire n1693, n59949, n1694, n59948, n1695, n59947, n1696, n59946, 
        n59017, n1697, n59945, n37_adj_4604, n1698, n59944, n1699, 
        n59943, n1700, n59942, n35_adj_4605, n59016, n1701, n59941, 
        n1552, n59940, n1553, n59939, n39_adj_4606, n1554, n59938, 
        n1555, n59937, n34_adj_4607, n1556, n59936, n1557, n59935, 
        n59934, n59933, n59932, n59015;
    wire [23:0]n8345;
    
    wire n59931, n1409, n59930, n1410, n59929, n1411, n59928, 
        n1412, n59927, n59926, n59925, n1415, n59924;
    wire [23:0]n8319;
    
    wire n1261, n59923, n1262, n59922, n1263, n59921, n59014, 
        n1264, n59920, n59919, n59918, n59917, n59013, n39_adj_4608, 
        n70070;
    wire [23:0]n8293;
    
    wire n59916, n1112, n59915, n1113, n59914, n59913, n59912, 
        n1116, n59911, n59012, n37_adj_4609, n43_adj_4610, n26029, 
        n48_adj_4611, n59011, n59010, n41_adj_4612, n59009, n75446, 
        n34_adj_4613, n43_adj_4614, n59008, n59007, n37_adj_4615, 
        n41_adj_4616, n71486, n39_adj_4617, n71488, n71416, n71418, 
        n70620, n67918, n32_adj_4618, n77906, n77907, n76392;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n77247, n77632, n77904, n77905, n71358, n71364, n43_adj_4619, 
        n37_adj_4620, n41_adj_4621, n39_adj_4622, n25967, n32_adj_4623, 
        n71362, n70602, n77645, n77646, n76408, n77245, n77628, 
        n77639, n77640, n45_adj_4624, n39_adj_4625, n43_adj_4626, 
        n41_adj_4627, n41_adj_4628, n959, n44_adj_4629, n46, n67645, 
        n960, n11692, n21189, n961, n40_adj_4630, n962, n43_adj_4631, 
        n26035, n48_adj_4632, n38_adj_4633, n42_adj_4634, n77655, 
        n803, n44_adj_4635, n46_adj_4636, n67643, n60289, n60288, 
        n60287, n804, n21179, n25970, n805, n25991, n48_adj_4637, 
        n44854, n68378, n644, n44_adj_4638, n46_adj_4639, n67641, 
        n75551, n48_adj_4640, n26022, n25988, n48_adj_4641, n68402, 
        n5, n72202, n71360, n70512, n25937, n70444, n72206, n72190, 
        n72116, n70486, n72118, n72216, n72218, n45376, n75548, 
        n70552, n70556, n75234, n46_adj_4642, n42_adj_4643, n77666, 
        n77667, n48_adj_4644, n25976, n67935, n42_adj_4645, n77662, 
        n77663, n36_adj_4646, n40_adj_4647, n78153, n78154, n12_adj_4648, 
        n78090, n75994, n14_adj_4649, n34_adj_4650, n77896, n77897, 
        n76414, n38_adj_4651, n44_adj_4652, n16_adj_4653, n75968, 
        n18_adj_4654, n31_adj_4655, n75205, n33_adj_4656, n35_adj_4657, 
        n66553, n75211, n75202, n29_adj_4658, n75208, n75428, n32_adj_4659, 
        n40_adj_4660, n28_adj_4661, n77900, n77901, n75422, n30_adj_4662, 
        n75416, n77898, n77636, n78172, n71490, n71438, n71442, 
        n29_adj_4663, n31_adj_4664, n33_adj_4665, n27_adj_4666, n75386, 
        n30_adj_4667, n38_adj_4668, n26_adj_4669, n77892, n77893, 
        n75382, n28_adj_4670, n75379, n78155, n77642, n78253, n78254, 
        n78228, n48_adj_4671, n26010, n27_adj_4672, n75368, n30_adj_4673, 
        n38_adj_4674, n67909, n26_adj_4675, n77888, n77889, n75362, 
        n28_adj_4676, n75359, n78159, n77648, n78255, n78256, n78226, 
        n48_adj_4677, n72224, n72196, n23_adj_4678, n75348, n75344, 
        n22_adj_4679, n28_adj_4680, n30_adj_4681, n26_adj_4682, n34_adj_4683, 
        n24_adj_4684, n75338, n78073, n78074, n77925, n77521, n75346, 
        n78081, n76583, n78165, n78166, n14_adj_4685, n71462, n26016, 
        n21_adj_4686, n76293, n76285, n20_adj_4687, n26_adj_4688, 
        n28_adj_4689, n24_adj_4690, n32_adj_4691, n22_adj_4692, n76283, 
        n78075, n78076, n77923, n77813, n76289, n78077, n76587, 
        n78149, n78150, n78113, n76054, n16_adj_4693, n18_adj_4694, 
        n25_adj_4695, n27_adj_4696, n19_adj_4697, n76239, n76227, 
        n76022, n77807, n18_adj_4698, n77613, n77614, n76234, n77085, 
        n24_adj_4699, n26_adj_4700, n76599, n22_adj_4701, n30_adj_4702, 
        n20_adj_4703, n76215, n78087, n78088, n77903, n77087, n77657, 
        n76597, n77659, n20_adj_4704, n23_adj_4705, n25_adj_4706, 
        n17_adj_4707, n76175, n76167, n77803, n16_adj_4708, n77607, 
        n77608, n76171, n77043, n22_adj_4709, n77660, n76607, n71436, 
        n20_adj_4710, n28_adj_4711, n18_adj_4712, n76160, n78091, 
        n78092, n77881, n77045, n77876, n76605, n78170, n78171, 
        n19_adj_4713, n21_adj_4714, n23_adj_4715, n76036, n76999, 
        n77441, n77437, n76040, n12_adj_4716, n77597, n38_adj_4717, 
        n77598, n76028, n78079, n76623, n24_adj_4718, n78097, n78098, 
        n77863, n77785, n78223, n76621, n78257, n78258, n17_adj_4719, 
        n19_adj_4720, n21_adj_4721, n33_adj_4722, n25973, n75982, 
        n76945, n77413, n77409, n75984, n10_adj_4723, n77591, n77592, 
        n36_adj_4724, n75974, n77866, n76629, n22_adj_4725, n77860, 
        n77861, n77857, n77775, n78231, n76627, n78269, n78270, 
        n78268, n75188, n75185, n75182, n70156, n70162, n25979, 
        n6_adj_4726, n69436, n14_adj_4727, n15_adj_4728, n70328, n70334, 
        n70104, n70344, n70350, n70264, n70270, n70312, n70318, 
        n70296, n70302, n70376, n70382, n70624, n3_adj_4729, n70360, 
        n70366, n70628, n5_adj_4730, n70632, n8_adj_4731, n70196, 
        n70202, n72154, n72220, n2, n11917, n70138, n70062;
    
    SB_LUT4 r_Clock_Count_2053_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n60285), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_5 (.CI(n60285), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n60286));
    SB_LUT4 r_Clock_Count_2053_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n60284), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_4 (.CI(n60284), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n60285));
    SB_LUT4 r_Clock_Count_2053_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n60283), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_3 (.CI(n60283), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n60284));
    SB_LUT4 r_Clock_Count_2053_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n60283));
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8683[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8683[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8683[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8683[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8683[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8683[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28240), 
            .D(n479[1]), .R(n67800));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8683[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28240), 
            .D(n479[2]), .R(n67800));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 i60358_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5217), .I3(n66790), .O(n75177));
    defparam i60358_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i60355_4_lut (.I0(n75177), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n75174));
    defparam i60355_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n75174), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n28117));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i1_4_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70280), .O(n70286));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_968 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70286), .O(n70292));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_968.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8683[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8683[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8683[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8683[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8683[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8683[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8683[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8657[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8657[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8657[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8657[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8657[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8657[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8657[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8657[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8657[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8657[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4455));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4456));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8657[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8657[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4457));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8657[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8657[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8657[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8657[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8657[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8657[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8657[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60057_4_lut (.I0(n31), .I1(n19), .I2(n17), .I3(n15), .O(n75913));
    defparam i60057_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61029_4_lut (.I0(n13), .I1(n11), .I2(n3065), .I3(baudrate[2]), 
            .O(n76885));
    defparam i61029_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i61525_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n76885), 
            .O(n77381));
    defparam i61525_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i56337_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), .I2(baudrate[12]), 
            .I3(baudrate[11]), .O(n72184));
    defparam i56337_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61521_4_lut (.I0(n25), .I1(n23_adj_4457), .I2(n21), .I3(n77381), 
            .O(n77377));
    defparam i61521_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60061_4_lut (.I0(n31), .I1(n29_adj_4456), .I2(n27_adj_4455), 
            .I3(n77377), .O(n75917));
    defparam i60061_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i56383_2_lut_3_lut (.I0(baudrate[13]), .I1(baudrate[14]), .I2(n72228), 
            .I3(GND_net), .O(n72230));
    defparam i56383_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61725_3_lut (.I0(n8), .I1(baudrate[13]), .I2(n31), .I3(GND_net), 
            .O(n77581));   // verilog/uart_rx.v(119[33:55])
    defparam i61725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61726_3_lut (.I0(n77581), .I1(baudrate[14]), .I2(n33), .I3(GND_net), 
            .O(n77582));   // verilog/uart_rx.v(119[33:55])
    defparam i61726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16), .I1(baudrate[17]), 
            .I2(n39), .I3(GND_net), .O(n34_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(n78173), .I1(baudrate[11]), .I2(n1831), 
            .I3(n70074), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 i60050_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n75913), 
            .O(n75906));
    defparam i60050_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62014_4_lut (.I0(n34_c), .I1(n14), .I2(n39), .I3(n75902), 
            .O(n77870));   // verilog/uart_rx.v(119[33:55])
    defparam i62014_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60785_3_lut (.I0(n77582), .I1(baudrate[15]), .I2(n35), .I3(GND_net), 
            .O(n76641));   // verilog/uart_rx.v(119[33:55])
    defparam i60785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61727_3_lut (.I0(n10), .I1(baudrate[10]), .I2(n25), .I3(GND_net), 
            .O(n77583));   // verilog/uart_rx.v(119[33:55])
    defparam i61727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61728_3_lut (.I0(n77583), .I1(baudrate[11]), .I2(n27_adj_4455), 
            .I3(GND_net), .O(n77584));   // verilog/uart_rx.v(119[33:55])
    defparam i61728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61009_4_lut (.I0(n27_adj_4455), .I1(n25), .I2(n23_adj_4457), 
            .I3(n75928), .O(n76865));
    defparam i61009_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12), .I1(baudrate[9]), 
            .I2(n23_adj_4457), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60783_3_lut (.I0(n77584), .I1(baudrate[12]), .I2(n29_adj_4456), 
            .I3(GND_net), .O(n76639));   // verilog/uart_rx.v(119[33:55])
    defparam i60783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61905_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n75917), 
            .O(n77761));
    defparam i61905_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62377_4_lut (.I0(n76641), .I1(n77870), .I2(n39), .I3(n75906), 
            .O(n78233));   // verilog/uart_rx.v(119[33:55])
    defparam i62377_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61814_4_lut (.I0(n76639), .I1(n20), .I2(n29_adj_4456), .I3(n76865), 
            .O(n77670));   // verilog/uart_rx.v(119[33:55])
    defparam i61814_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i63199_2_lut_4_lut (.I0(n78173), .I1(baudrate[11]), .I2(n1831), 
            .I3(n72232), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i63199_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i62403_4_lut (.I0(n77670), .I1(n78233), .I2(n39), .I3(n77761), 
            .O(n78259));   // verilog/uart_rx.v(119[33:55])
    defparam i62403_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62404_3_lut (.I0(n78259), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n78260));   // verilog/uart_rx.v(119[33:55])
    defparam i62404_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62028_3_lut (.I0(n78260), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n77884));   // verilog/uart_rx.v(119[33:55])
    defparam i62028_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62029_3_lut (.I0(n77884), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n77885));   // verilog/uart_rx.v(119[33:55])
    defparam i62029_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8631[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8631[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i63191_2_lut_4_lut (.I0(n77243), .I1(baudrate[8]), .I2(n1408), 
            .I3(n72242), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i63191_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8631[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4458));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8631[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8631[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8631[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8631[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8631[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4461));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4462));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8631[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8631[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8631[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4463));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4464));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4465));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_969 (.I0(n77243), .I1(baudrate[8]), .I2(n1408), 
            .I3(n70072), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_969.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8631[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8631[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8631[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4466));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4467));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8631[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8631[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8605[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8605[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8605[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4468));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8605[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4469));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8605[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4470));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8605[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4471));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8605[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8605[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8605[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4472));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4473));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4474));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8605[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8605[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8605[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(n71350), .I1(n72232), .I2(n8371[14]), 
            .I3(n48), .O(n1702));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4475));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8605[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8605[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8605[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29937));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29936));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29934));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29915));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8579[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8579[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8579[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29914));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29910));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29906));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8579[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8579[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n79649));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8579[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8579[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8579[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8579[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8579[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8579[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8579[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8579[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8579[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i56395_2_lut_3_lut (.I0(n71350), .I1(n72232), .I2(baudrate[9]), 
            .I3(GND_net), .O(n72242));
    defparam i56395_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i63196_2_lut_3_lut (.I0(n71350), .I1(n72232), .I2(n48), .I3(GND_net), 
            .O(n294[14]));
    defparam i63196_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i59616_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n75472));   // verilog/uart_rx.v(119[33:55])
    defparam i59616_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8579[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4491));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4492));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4493));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4494));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR r_Clock_Count_2053__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n28161), .D(n1[0]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n28161), .D(n1[1]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n28161), .D(n1[2]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n28161), .D(n1[3]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n28161), .D(n1[4]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n28161), .D(n1[5]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n28161), .D(n1[6]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n28161), .D(n1[7]), .R(n29423));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i60236_4_lut (.I0(n37_adj_4494), .I1(n25_adj_4493), .I2(n23_adj_4492), 
            .I3(n21_adj_4491), .O(n76092));
    defparam i60236_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61181_4_lut (.I0(n19_adj_4490), .I1(n17_adj_4489), .I2(n2729), 
            .I3(baudrate[2]), .O(n77037));
    defparam i61181_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i61603_4_lut (.I0(n25_adj_4493), .I1(n23_adj_4492), .I2(n21_adj_4491), 
            .I3(n77037), .O(n77459));
    defparam i61603_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61601_4_lut (.I0(n31_adj_4486), .I1(n29_adj_4485), .I2(n27_adj_4484), 
            .I3(n77459), .O(n77457));
    defparam i61601_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60238_4_lut (.I0(n37_adj_4494), .I1(n35_adj_4488), .I2(n33_adj_4487), 
            .I3(n77457), .O(n76094));
    defparam i60238_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_4497));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61745_3_lut (.I0(n14_adj_4497), .I1(baudrate[13]), .I2(n37_adj_4494), 
            .I3(GND_net), .O(n77601));   // verilog/uart_rx.v(119[33:55])
    defparam i61745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61746_3_lut (.I0(n77601), .I1(baudrate[14]), .I2(n39_adj_4482), 
            .I3(GND_net), .O(n77602));   // verilog/uart_rx.v(119[33:55])
    defparam i61746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22), .I1(baudrate[17]), 
            .I2(n45_adj_4481), .I3(GND_net), .O(n40_adj_4498));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60226_4_lut (.I0(n43_adj_4483), .I1(n41_adj_4480), .I2(n39_adj_4482), 
            .I3(n76092), .O(n76082));
    defparam i60226_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61808_4_lut (.I0(n40_adj_4498), .I1(n20_adj_4499), .I2(n45_adj_4481), 
            .I3(n76078), .O(n77664));   // verilog/uart_rx.v(119[33:55])
    defparam i61808_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i60761_3_lut (.I0(n77602), .I1(baudrate[15]), .I2(n41_adj_4480), 
            .I3(GND_net), .O(n76617));   // verilog/uart_rx.v(119[33:55])
    defparam i60761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18), .I1(baudrate[9]), 
            .I2(n29_adj_4485), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62237_4_lut (.I0(n26), .I1(n16_adj_4500), .I2(n29_adj_4485), 
            .I3(n76108), .O(n78093));   // verilog/uart_rx.v(119[33:55])
    defparam i62237_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62238_3_lut (.I0(n78093), .I1(baudrate[10]), .I2(n31_adj_4486), 
            .I3(GND_net), .O(n78094));   // verilog/uart_rx.v(119[33:55])
    defparam i62238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62017_3_lut (.I0(n78094), .I1(baudrate[11]), .I2(n33_adj_4487), 
            .I3(GND_net), .O(n77873));   // verilog/uart_rx.v(119[33:55])
    defparam i62017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61939_4_lut (.I0(n43_adj_4483), .I1(n41_adj_4480), .I2(n39_adj_4482), 
            .I3(n76094), .O(n77795));
    defparam i61939_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62249_4_lut (.I0(n76617), .I1(n77664), .I2(n45_adj_4481), 
            .I3(n76082), .O(n78105));   // verilog/uart_rx.v(119[33:55])
    defparam i62249_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2903_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n60147), 
            .O(n8709[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2903_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n60146), 
            .O(n8709[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_24 (.CI(n60146), .I0(n3152), .I1(n3082), .CO(n60147));
    SB_LUT4 add_2903_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n60145), 
            .O(n8709[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60759_3_lut (.I0(n77873), .I1(baudrate[12]), .I2(n35_adj_4488), 
            .I3(GND_net), .O(n76615));   // verilog/uart_rx.v(119[33:55])
    defparam i60759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62251_4_lut (.I0(n76615), .I1(n78105), .I2(n45_adj_4481), 
            .I3(n77795), .O(n78107));   // verilog/uart_rx.v(119[33:55])
    defparam i62251_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2903_23 (.CI(n60145), .I0(n3153), .I1(n3188), .CO(n60146));
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8579[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8605[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2903_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n60144), 
            .O(n8709[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_22 (.CI(n60144), .I0(n3154), .I1(n3084), .CO(n60145));
    SB_LUT4 add_2903_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n60143), 
            .O(n8709[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_21 (.CI(n60143), .I0(n3155), .I1(n2977), .CO(n60144));
    SB_LUT4 add_2903_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n60142), 
            .O(n8709[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_20 (.CI(n60142), .I0(n3156), .I1(n2867), .CO(n60143));
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8553[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8553[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2903_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n60141), 
            .O(n8709[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_19 (.CI(n60141), .I0(n3157), .I1(n2754), .CO(n60142));
    SB_LUT4 add_2903_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n60140), 
            .O(n8709[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n30762));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n62510));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30758));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8553[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2903_18 (.CI(n60140), .I0(n3158), .I1(n2638), .CO(n60141));
    SB_LUT4 add_2903_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n60139), 
            .O(n8709[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_17 (.CI(n60139), .I0(n3159), .I1(n2519), .CO(n60140));
    SB_LUT4 add_2903_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n60138), 
            .O(n8709[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_16 (.CI(n60138), .I0(n3160), .I1(n2397), .CO(n60139));
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4501));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2903_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n60137), 
            .O(n8709[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_15 (.CI(n60137), .I0(n3161), .I1(n2272), .CO(n60138));
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8553[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2903_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n60136), 
            .O(n8709[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_14 (.CI(n60136), .I0(n3162), .I1(n2144), .CO(n60137));
    SB_LUT4 add_2903_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n60135), 
            .O(n8709[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_13 (.CI(n60135), .I0(n3163), .I1(n2013), .CO(n60136));
    SB_LUT4 add_2903_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n60134), 
            .O(n8709[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_12 (.CI(n60134), .I0(n3164), .I1(n1879), .CO(n60135));
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4502));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8553[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2903_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n60133), 
            .O(n8709[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_11 (.CI(n60133), .I0(n3165), .I1(n1742), .CO(n60134));
    SB_LUT4 i56398_1_lut_2_lut (.I0(baudrate[8]), .I1(n72242), .I2(GND_net), 
            .I3(GND_net), .O(n67928));
    defparam i56398_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 add_2903_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n60132), 
            .O(n8709[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_10 (.CI(n60132), .I0(n3166), .I1(n1602), .CO(n60133));
    SB_LUT4 add_2903_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n60131), 
            .O(n8709[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_9 (.CI(n60131), .I0(n3167), .I1(n1459), .CO(n60132));
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4503));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8553[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2903_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n60130), 
            .O(n8709[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_8 (.CI(n60130), .I0(n3168), .I1(n1460), .CO(n60131));
    SB_LUT4 add_2903_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n60129), 
            .O(n8709[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_7 (.CI(n60129), .I0(n3169), .I1(n1011), .CO(n60130));
    SB_LUT4 add_2903_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n60128), 
            .O(n8709[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4504));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2903_6 (.CI(n60128), .I0(n3170), .I1(n856), .CO(n60129));
    SB_LUT4 add_2903_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n60127), 
            .O(n8709[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_5 (.CI(n60127), .I0(n3171), .I1(n698), .CO(n60128));
    SB_LUT4 add_2903_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n60126), 
            .O(n8709[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_4 (.CI(n60126), .I0(n3172), .I1(n858), .CO(n60127));
    SB_LUT4 add_2903_3_lut (.I0(n67874), .I1(GND_net), .I2(n538), .I3(n60125), 
            .O(n70092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8553[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2903_3 (.CI(n60125), .I0(GND_net), .I1(n538), .CO(n60126));
    SB_CARRY add_2903_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n60125));
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8553[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4505));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4506));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2902_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n60124), 
            .O(n8683[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i56399_2_lut_3_lut (.I0(baudrate[8]), .I1(n72242), .I2(baudrate[7]), 
            .I3(GND_net), .O(n72246));
    defparam i56399_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 add_2902_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n60123), 
            .O(n8683[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8553[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2902_22 (.CI(n60123), .I0(n3047), .I1(n3188), .CO(n60124));
    SB_LUT4 add_2902_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n60122), 
            .O(n8683[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_21 (.CI(n60122), .I0(n3048), .I1(n3084), .CO(n60123));
    SB_LUT4 add_2902_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n60121), 
            .O(n8683[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8553[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2902_20 (.CI(n60121), .I0(n3049), .I1(n2977), .CO(n60122));
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8553[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i63188_2_lut_3_lut (.I0(baudrate[8]), .I1(n72242), .I2(n48_adj_4507), 
            .I3(GND_net), .O(n294[16]));
    defparam i63188_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8553[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2902_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n60120), 
            .O(n8683[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4508));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4509));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2902_19 (.CI(n60120), .I0(n3050), .I1(n2867), .CO(n60121));
    SB_LUT4 add_2902_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n60119), 
            .O(n8683[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4510));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2902_18 (.CI(n60119), .I0(n3051), .I1(n2754), .CO(n60120));
    SB_LUT4 add_2902_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n60118), 
            .O(n8683[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_17 (.CI(n60118), .I0(n3052), .I1(n2638), .CO(n60119));
    SB_LUT4 add_2902_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n60117), 
            .O(n8683[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8709[20]), .I3(n294[1]), .O(n41_adj_4511));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8709[19]), .I3(n294[1]), .O(n39_adj_4512));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8553[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8709[14]), .I3(n294[1]), .O(n29_adj_4513));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4514));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8709[15]), .I3(n294[1]), .O(n31_adj_4515));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8709[18]), .I3(n294[1]), .O(n37_adj_4516));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8709[11]), .I3(n294[1]), .O(n23_adj_4517));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8709[12]), .I3(n294[1]), .O(n25_adj_4518));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8709[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8709[22]), .I3(n294[1]), .O(n45_adj_4519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8709[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4520));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8709[8]), .I3(n294[1]), .O(n17_adj_4521));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2902_16 (.CI(n60117), .I0(n3053), .I1(n2519), .CO(n60118));
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8527[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2902_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n60116), 
            .O(n8683[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8527[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8527[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2902_15 (.CI(n60116), .I0(n3054), .I1(n2397), .CO(n60117));
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8709[10]), .I3(n294[1]), .O(n21_adj_4522));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8709[9]), .I3(n294[1]), .O(n19_adj_4523));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8709[21]), .I3(n294[1]), .O(n43_adj_4524));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8709[16]), .I3(n294[1]), .O(n33_adj_4525));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4526));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8709[17]), .I3(n294[1]), .O(n35_adj_4527));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8709[5]), .I3(n294[1]), .O(n11_adj_4528));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8709[6]), .I3(n294[1]), .O(n13_adj_4529));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8709[7]), .I3(n294[1]), .O(n15_adj_4530));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8709[13]), .I3(n294[1]), .O(n27_adj_4531));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8527[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59963_4_lut (.I0(n27_adj_4531), .I1(n15_adj_4530), .I2(n13_adj_4529), 
            .I3(n11_adj_4528), .O(n75819));
    defparam i59963_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2902_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n60115), 
            .O(n8683[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4532));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2902_14 (.CI(n60115), .I0(n3055), .I1(n2272), .CO(n60116));
    SB_LUT4 add_2902_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n60114), 
            .O(n8683[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_13 (.CI(n60114), .I0(n3056), .I1(n2144), .CO(n60115));
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8527[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_4525), .I3(GND_net), .O(n12_adj_4533));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59955_2_lut (.I0(n33_adj_4525), .I1(n15_adj_4530), .I2(GND_net), 
            .I3(GND_net), .O(n75811));
    defparam i59955_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13_adj_4529), .I3(GND_net), .O(n10_adj_4534));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2902_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n60113), 
            .O(n8683[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_12 (.CI(n60113), .I0(n3057), .I1(n2013), .CO(n60114));
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4535));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_4533), .I1(baudrate[17]), 
            .I2(n35_adj_4527), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2902_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n60112), 
            .O(n8683[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_11 (.CI(n60112), .I0(n3058), .I1(n1879), .CO(n60113));
    SB_LUT4 add_2902_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n60111), 
            .O(n8683[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_10 (.CI(n60111), .I0(n3059), .I1(n1742), .CO(n60112));
    SB_LUT4 add_2902_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n60110), 
            .O(n8683[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_9 (.CI(n60110), .I0(n3060), .I1(n1602), .CO(n60111));
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8527[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2902_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n60109), 
            .O(n8683[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59971_4_lut (.I0(n21_adj_4522), .I1(n19_adj_4523), .I2(n17_adj_4521), 
            .I3(n9), .O(n75827));
    defparam i59971_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2902_8 (.CI(n60109), .I0(n3061), .I1(n1459), .CO(n60110));
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_4524), .I3(GND_net), .O(n16_adj_4536));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4537));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2902_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n60108), 
            .O(n8683[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59943_2_lut (.I0(n43_adj_4524), .I1(n19_adj_4523), .I2(GND_net), 
            .I3(GND_net), .O(n75799));
    defparam i59943_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8527[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2902_7 (.CI(n60108), .I0(n3062), .I1(n1460), .CO(n60109));
    SB_LUT4 add_2902_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n60107), 
            .O(n8683[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_6 (.CI(n60107), .I0(n3063), .I1(n1011), .CO(n60108));
    SB_LUT4 add_2902_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n60106), 
            .O(n8683[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_4521), .I3(GND_net), .O(n8_adj_4538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8527[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_4536), .I1(baudrate[22]), 
            .I2(n45_adj_4519), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2902_5 (.CI(n60106), .I0(n3064), .I1(n856), .CO(n60107));
    SB_LUT4 add_2902_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n60105), 
            .O(n8683[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8709[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59981_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n75837));
    defparam i59981_3_lut.LUT_INIT = 16'hbebe;
    SB_CARRY add_2902_4 (.CI(n60105), .I0(n3065), .I1(n698), .CO(n60106));
    SB_LUT4 add_2902_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n60104), 
            .O(n8683[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60933_4_lut (.I0(n13_adj_4529), .I1(n11_adj_4528), .I2(n9), 
            .I3(n75837), .O(n76789));
    defparam i60933_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2902_3 (.CI(n60104), .I0(n3066), .I1(n858), .CO(n60105));
    SB_LUT4 add_2902_2_lut (.I0(n67878), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2902_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n60104));
    SB_LUT4 add_2901_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n60103), 
            .O(n8657[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60927_4_lut (.I0(n19_adj_4523), .I1(n17_adj_4521), .I2(n15_adj_4530), 
            .I3(n76789), .O(n76783));
    defparam i60927_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2901_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n60102), 
            .O(n8657[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8527[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2901_21 (.CI(n60102), .I0(n2939), .I1(n3084), .CO(n60103));
    SB_LUT4 i62100_4_lut (.I0(n25_adj_4518), .I1(n23_adj_4517), .I2(n21_adj_4522), 
            .I3(n76783), .O(n77956));
    defparam i62100_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4539));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2901_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n60101), 
            .O(n8657[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4540));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4541));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2901_20 (.CI(n60101), .I0(n2940), .I1(n2977), .CO(n60102));
    SB_LUT4 i61463_4_lut (.I0(n31_adj_4515), .I1(n29_adj_4513), .I2(n27_adj_4531), 
            .I3(n77956), .O(n77319));
    defparam i61463_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i62264_4_lut (.I0(n37_adj_4516), .I1(n35_adj_4527), .I2(n33_adj_4525), 
            .I3(n77319), .O(n78120));
    defparam i62264_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2901_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n60100), 
            .O(n8657[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_19 (.CI(n60100), .I0(n2941), .I1(n2867), .CO(n60101));
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2901_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n60099), 
            .O(n8657[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_18 (.CI(n60099), .I0(n2942), .I1(n2754), .CO(n60100));
    SB_LUT4 add_2901_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n60098), 
            .O(n8657[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_17 (.CI(n60098), .I0(n2943), .I1(n2638), .CO(n60099));
    SB_LUT4 i61689_3_lut (.I0(n6), .I1(baudrate[10]), .I2(n21_adj_4522), 
            .I3(GND_net), .O(n77545));   // verilog/uart_rx.v(119[33:55])
    defparam i61689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2901_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n60097), 
            .O(n8657[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_16 (.CI(n60097), .I0(n2944), .I1(n2519), .CO(n60098));
    SB_LUT4 i61690_3_lut (.I0(n77545), .I1(baudrate[11]), .I2(n23_adj_4517), 
            .I3(GND_net), .O(n77546));   // verilog/uart_rx.v(119[33:55])
    defparam i61690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n70092), .I3(n48_adj_4542), .O(n4));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 add_2901_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n60096), 
            .O(n8657[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_15 (.CI(n60096), .I0(n2945), .I1(n2397), .CO(n60097));
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8527[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61687_3_lut (.I0(n4), .I1(baudrate[13]), .I2(n27_adj_4531), 
            .I3(GND_net), .O(n77543));   // verilog/uart_rx.v(119[33:55])
    defparam i61687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2901_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n60095), 
            .O(n8657[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_14 (.CI(n60095), .I0(n2946), .I1(n2272), .CO(n60096));
    SB_LUT4 add_2901_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n60094), 
            .O(n8657[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_13 (.CI(n60094), .I0(n2947), .I1(n2144), .CO(n60095));
    SB_LUT4 add_2901_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n60093), 
            .O(n8657[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_12 (.CI(n60093), .I0(n2948), .I1(n2013), .CO(n60094));
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8527[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61688_3_lut (.I0(n77543), .I1(baudrate[14]), .I2(n29_adj_4513), 
            .I3(GND_net), .O(n77544));   // verilog/uart_rx.v(119[33:55])
    defparam i61688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59957_4_lut (.I0(n33_adj_4525), .I1(n31_adj_4515), .I2(n29_adj_4513), 
            .I3(n75819), .O(n75813));
    defparam i59957_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62148_4_lut (.I0(n30), .I1(n10_adj_4534), .I2(n35_adj_4527), 
            .I3(n75811), .O(n78004));   // verilog/uart_rx.v(119[33:55])
    defparam i62148_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2901_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n60092), 
            .O(n8657[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_11 (.CI(n60092), .I0(n2949), .I1(n1879), .CO(n60093));
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_4543));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59639_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n75495));   // verilog/uart_rx.v(119[33:55])
    defparam i59639_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i56409_2_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(n72246), 
            .I3(GND_net), .O(n72256));
    defparam i56409_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i60810_3_lut (.I0(n77544), .I1(baudrate[15]), .I2(n31_adj_4515), 
            .I3(GND_net), .O(n76666));   // verilog/uart_rx.v(119[33:55])
    defparam i60810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62355_4_lut (.I0(n76666), .I1(n78004), .I2(n35_adj_4527), 
            .I3(n75813), .O(n78211));   // verilog/uart_rx.v(119[33:55])
    defparam i62355_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62356_3_lut (.I0(n78211), .I1(baudrate[18]), .I2(n37_adj_4516), 
            .I3(GND_net), .O(n78212));   // verilog/uart_rx.v(119[33:55])
    defparam i62356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62288_3_lut (.I0(n78212), .I1(baudrate[19]), .I2(n39_adj_4512), 
            .I3(GND_net), .O(n78144));   // verilog/uart_rx.v(119[33:55])
    defparam i62288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2901_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n60091), 
            .O(n8657[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_10 (.CI(n60091), .I0(n2950), .I1(n1742), .CO(n60092));
    SB_LUT4 add_2901_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n60090), 
            .O(n8657[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_9 (.CI(n60090), .I0(n2951), .I1(n1602), .CO(n60091));
    SB_LUT4 add_2901_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n60089), 
            .O(n8657[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_8 (.CI(n60089), .I0(n2952), .I1(n1459), .CO(n60090));
    SB_LUT4 i59945_4_lut (.I0(n43_adj_4524), .I1(n25_adj_4518), .I2(n23_adj_4517), 
            .I3(n75827), .O(n75801));
    defparam i59945_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2901_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n60088), 
            .O(n8657[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_7 (.CI(n60088), .I0(n2953), .I1(n1460), .CO(n60089));
    SB_LUT4 i61822_4_lut (.I0(n24), .I1(n8_adj_4538), .I2(n45_adj_4519), 
            .I3(n75799), .O(n77678));   // verilog/uart_rx.v(119[33:55])
    defparam i61822_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4544));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2901_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n60087), 
            .O(n8657[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60808_3_lut (.I0(n77546), .I1(baudrate[12]), .I2(n25_adj_4518), 
            .I3(GND_net), .O(n76664));   // verilog/uart_rx.v(119[33:55])
    defparam i60808_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2901_6 (.CI(n60087), .I0(n2954), .I1(n1011), .CO(n60088));
    SB_LUT4 i59947_4_lut (.I0(n43_adj_4524), .I1(n41_adj_4511), .I2(n39_adj_4512), 
            .I3(n78120), .O(n75803));
    defparam i59947_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4545));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62252_4_lut (.I0(n76664), .I1(n77678), .I2(n45_adj_4519), 
            .I3(n75801), .O(n78108));   // verilog/uart_rx.v(119[33:55])
    defparam i62252_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2901_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n60086), 
            .O(n8657[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_5 (.CI(n60086), .I0(n2955), .I1(n856), .CO(n60087));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[4]), 
            .I3(baudrate[3]), .O(n70554));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8527[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60816_3_lut (.I0(n78144), .I1(baudrate[20]), .I2(n41_adj_4511), 
            .I3(GND_net), .O(n76672));   // verilog/uart_rx.v(119[33:55])
    defparam i60816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8527[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8709[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2901_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n60085), 
            .O(n8657[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_4 (.CI(n60085), .I0(n2956), .I1(n698), .CO(n60086));
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4546));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4547));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62254_4_lut (.I0(n76672), .I1(n78108), .I2(n45_adj_4519), 
            .I3(n75803), .O(n78110));   // verilog/uart_rx.v(119[33:55])
    defparam i62254_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8501[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2901_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n60084), 
            .O(n8657[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8501[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2901_3 (.CI(n60084), .I0(n2957), .I1(n858), .CO(n60085));
    SB_LUT4 add_2901_2_lut (.I0(n67882), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2901_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n60084));
    SB_LUT4 i62838_4_lut (.I0(n70018), .I1(n78110), .I2(baudrate[23]), 
            .I3(n3253), .O(n69091));   // verilog/uart_rx.v(119[33:55])
    defparam i62838_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 add_2900_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n60083), 
            .O(n8631[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2900_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n60082), 
            .O(n8631[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_20 (.CI(n60082), .I0(n2828), .I1(n2977), .CO(n60083));
    SB_LUT4 add_2900_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n60081), 
            .O(n8631[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_4548), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4549));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2900_19 (.CI(n60081), .I0(n2829), .I1(n2867), .CO(n60082));
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4550));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2900_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n60080), 
            .O(n8631[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_18 (.CI(n60080), .I0(n2830), .I1(n2754), .CO(n60081));
    SB_LUT4 add_2900_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n60079), 
            .O(n8631[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4551));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2900_17 (.CI(n60079), .I0(n2831), .I1(n2638), .CO(n60080));
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i56413_3_lut_4_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(baudrate[2]), 
            .I3(n72256), .O(n72260));
    defparam i56413_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8501[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8501[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2900_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n60078), 
            .O(n8631[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4560));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2900_16 (.CI(n60078), .I0(n2832), .I1(n2519), .CO(n60079));
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4561));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4562));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2900_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n60077), 
            .O(n8631[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4563));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2900_15 (.CI(n60077), .I0(n2833), .I1(n2397), .CO(n60078));
    SB_LUT4 add_2900_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n60076), 
            .O(n8631[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_14 (.CI(n60076), .I0(n2834), .I1(n2272), .CO(n60077));
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4564));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60010_4_lut (.I0(n29_adj_4563), .I1(n17_adj_4562), .I2(n15_adj_4561), 
            .I3(n13_adj_4560), .O(n75866));
    defparam i60010_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60979_4_lut (.I0(n11_adj_4558), .I1(n9_adj_4557), .I2(n3171), 
            .I3(baudrate[2]), .O(n76835));
    defparam i60979_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i61499_4_lut (.I0(n17_adj_4562), .I1(n15_adj_4561), .I2(n13_adj_4560), 
            .I3(n76835), .O(n77355));
    defparam i61499_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61497_4_lut (.I0(n23_adj_4554), .I1(n21_adj_4553), .I2(n19_adj_4559), 
            .I3(n77355), .O(n77353));
    defparam i61497_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60012_4_lut (.I0(n29_adj_4563), .I1(n27_adj_4556), .I2(n25_adj_4555), 
            .I3(n77353), .O(n75868));
    defparam i60012_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_4565));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61717_3_lut (.I0(n6_adj_4565), .I1(baudrate[13]), .I2(n29_adj_4563), 
            .I3(GND_net), .O(n77573));   // verilog/uart_rx.v(119[33:55])
    defparam i61717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8501[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2900_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n60075), 
            .O(n8631[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4566));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2900_13 (.CI(n60075), .I0(n2835), .I1(n2144), .CO(n60076));
    SB_LUT4 add_2900_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n60074), 
            .O(n8631[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_4567), .I1(baudrate[17]), 
            .I2(n37_adj_4551), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_12 (.CI(n60074), .I0(n2836), .I1(n2013), .CO(n60075));
    SB_LUT4 add_2900_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n60073), 
            .O(n8631[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61718_3_lut (.I0(n77573), .I1(baudrate[14]), .I2(n31_adj_4550), 
            .I3(GND_net), .O(n77574));   // verilog/uart_rx.v(119[33:55])
    defparam i61718_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_11 (.CI(n60073), .I0(n2837), .I1(n1879), .CO(n60074));
    SB_LUT4 i59999_4_lut (.I0(n35_adj_4552), .I1(n33_adj_4549), .I2(n31_adj_4550), 
            .I3(n75866), .O(n75855));
    defparam i59999_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62126_4_lut (.I0(n32), .I1(n12_adj_4568), .I2(n37_adj_4551), 
            .I3(n75853), .O(n77982));   // verilog/uart_rx.v(119[33:55])
    defparam i62126_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60796_3_lut (.I0(n77574), .I1(baudrate[15]), .I2(n33_adj_4549), 
            .I3(GND_net), .O(n76652));   // verilog/uart_rx.v(119[33:55])
    defparam i60796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61818_3_lut (.I0(n8_adj_4569), .I1(baudrate[10]), .I2(n23_adj_4554), 
            .I3(GND_net), .O(n77674));   // verilog/uart_rx.v(119[33:55])
    defparam i61818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61819_3_lut (.I0(n77674), .I1(baudrate[11]), .I2(n25_adj_4555), 
            .I3(GND_net), .O(n77675));   // verilog/uart_rx.v(119[33:55])
    defparam i61819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60965_4_lut (.I0(n25_adj_4555), .I1(n23_adj_4554), .I2(n21_adj_4553), 
            .I3(n75876), .O(n76821));
    defparam i60965_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61820_3_lut (.I0(n10_adj_4570), .I1(baudrate[9]), .I2(n21_adj_4553), 
            .I3(GND_net), .O(n77676));   // verilog/uart_rx.v(119[33:55])
    defparam i61820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60794_3_lut (.I0(n77675), .I1(baudrate[12]), .I2(n27_adj_4556), 
            .I3(GND_net), .O(n76650));   // verilog/uart_rx.v(119[33:55])
    defparam i60794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61899_4_lut (.I0(n35_adj_4552), .I1(n33_adj_4549), .I2(n31_adj_4550), 
            .I3(n75868), .O(n77755));
    defparam i61899_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62351_4_lut (.I0(n76652), .I1(n77982), .I2(n37_adj_4551), 
            .I3(n75855), .O(n78207));   // verilog/uart_rx.v(119[33:55])
    defparam i62351_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2900_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n60072), 
            .O(n8631[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61979_4_lut (.I0(n76650), .I1(n77676), .I2(n27_adj_4556), 
            .I3(n76821), .O(n77835));   // verilog/uart_rx.v(119[33:55])
    defparam i61979_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8501[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62415_4_lut (.I0(n77835), .I1(n78207), .I2(n37_adj_4551), 
            .I3(n77755), .O(n78271));   // verilog/uart_rx.v(119[33:55])
    defparam i62415_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2900_10 (.CI(n60072), .I0(n2838), .I1(n1742), .CO(n60073));
    SB_LUT4 i62416_3_lut (.I0(n78271), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n78272));   // verilog/uart_rx.v(119[33:55])
    defparam i62416_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62408_3_lut (.I0(n78272), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n78264));   // verilog/uart_rx.v(119[33:55])
    defparam i62408_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2900_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n60071), 
            .O(n8631[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62180_3_lut (.I0(n78264), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n78036));   // verilog/uart_rx.v(119[33:55])
    defparam i62180_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62181_3_lut (.I0(n78036), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n78037));   // verilog/uart_rx.v(119[33:55])
    defparam i62181_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60806_3_lut (.I0(n78037), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_4542));   // verilog/uart_rx.v(119[33:55])
    defparam i60806_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2900_9 (.CI(n60071), .I0(n2839), .I1(n1602), .CO(n60072));
    SB_LUT4 add_2900_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n60070), 
            .O(n8631[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_8 (.CI(n60070), .I0(n2840), .I1(n1459), .CO(n60071));
    SB_LUT4 add_2900_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n60069), 
            .O(n8631[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4571));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8501[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4572));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2900_7 (.CI(n60069), .I0(n2841), .I1(n1460), .CO(n60070));
    SB_LUT4 add_2900_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n60068), 
            .O(n8631[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_6 (.CI(n60068), .I0(n2842), .I1(n1011), .CO(n60069));
    SB_LUT4 add_2900_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n60067), 
            .O(n8631[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_5 (.CI(n60067), .I0(n2843), .I1(n856), .CO(n60068));
    SB_LUT4 add_2900_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n60066), 
            .O(n8631[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8501[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_4 (.CI(n60066), .I0(n2844), .I1(n698), .CO(n60067));
    SB_LUT4 add_2900_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n60065), 
            .O(n8631[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8501[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_3 (.CI(n60065), .I0(n2845), .I1(n858), .CO(n60066));
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8501[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2900_2_lut (.I0(n67886), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4573));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4574));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4575));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8501[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n60065));
    SB_LUT4 add_2899_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n60064), 
            .O(n8605[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2899_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n60063), 
            .O(n8605[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_19 (.CI(n60063), .I0(n2714), .I1(n2867), .CO(n60064));
    SB_LUT4 add_2899_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n60062), 
            .O(n8605[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_18 (.CI(n60062), .I0(n2715), .I1(n2754), .CO(n60063));
    SB_LUT4 i1_2_lut (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n71350));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_970 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n71354));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'heeee;
    SB_LUT4 add_2899_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n60061), 
            .O(n8605[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_17 (.CI(n60061), .I0(n2716), .I1(n2638), .CO(n60062));
    SB_LUT4 add_2899_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n60060), 
            .O(n8605[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_16 (.CI(n60060), .I0(n2717), .I1(n2519), .CO(n60061));
    SB_LUT4 add_2899_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n60059), 
            .O(n8605[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_15 (.CI(n60059), .I0(n2718), .I1(n2397), .CO(n60060));
    SB_LUT4 i1_2_lut_adj_971 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n71352));
    defparam i1_2_lut_adj_971.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_972 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n70588));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_973 (.I0(n70588), .I1(n71352), .I2(n71354), .I3(n71350), 
            .O(n70662));
    defparam i1_4_lut_adj_973.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_974 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n71474));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_975 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n71468));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_976 (.I0(baudrate[31]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n71470));
    defparam i1_2_lut_adj_976.LUT_INIT = 16'heeee;
    SB_LUT4 add_2899_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n60058), 
            .O(n8605[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_14 (.CI(n60058), .I0(n2719), .I1(n2272), .CO(n60059));
    SB_LUT4 add_2899_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n60057), 
            .O(n8605[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_13 (.CI(n60057), .I0(n2720), .I1(n2144), .CO(n60058));
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8501[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2899_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n60056), 
            .O(n8605[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8501[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_977 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n71472));
    defparam i1_2_lut_adj_977.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_978 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4576));
    defparam i1_2_lut_adj_978.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_979 (.I0(baudrate[24]), .I1(baudrate[26]), .I2(baudrate[25]), 
            .I3(baudrate[29]), .O(n14_adj_4577));
    defparam i1_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_CARRY add_2899_12 (.CI(n60056), .I0(n2721), .I1(n2013), .CO(n60057));
    SB_LUT4 i1_3_lut (.I0(n71468), .I1(n71474), .I2(baudrate[17]), .I3(GND_net), 
            .O(n71480));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 add_2899_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n60055), 
            .O(n8605[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_980 (.I0(n14_adj_4577), .I1(n9_adj_4576), .I2(n71480), 
            .I3(n71478), .O(n26019));
    defparam i1_4_lut_adj_980.LUT_INIT = 16'hfffe;
    SB_LUT4 i30763_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44852));
    defparam i30763_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2899_11 (.CI(n60055), .I0(n2722), .I1(n1879), .CO(n60056));
    SB_LUT4 add_2899_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n60054), 
            .O(n8605[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_981 (.I0(baudrate[2]), .I1(n42_adj_4578), 
            .I2(baudrate[3]), .I3(n21181), .O(n68370));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_981.LUT_INIT = 16'hff4f;
    SB_CARRY add_2899_10 (.CI(n60054), .I0(n2723), .I1(n1742), .CO(n60055));
    SB_LUT4 i16_4_lut (.I0(n70654), .I1(baudrate[16]), .I2(n28), .I3(n26019), 
            .O(n34));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2899_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n60053), 
            .O(n8605[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_9 (.CI(n60053), .I0(n2724), .I1(n1602), .CO(n60054));
    SB_LUT4 add_2899_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n60052), 
            .O(n8605[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_8 (.CI(n60052), .I0(n2725), .I1(n1459), .CO(n60053));
    SB_LUT4 add_2899_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n60051), 
            .O(n8605[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_7 (.CI(n60051), .I0(n2726), .I1(n1460), .CO(n60052));
    SB_LUT4 add_2899_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n60050), 
            .O(n8605[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_6 (.CI(n60050), .I0(n2727), .I1(n1011), .CO(n60051));
    SB_LUT4 add_2899_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n60049), 
            .O(n8605[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_5 (.CI(n60049), .I0(n2728), .I1(n856), .CO(n60050));
    SB_LUT4 add_2899_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n60048), 
            .O(n8605[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_4 (.CI(n60048), .I0(n2729), .I1(n698), .CO(n60049));
    SB_LUT4 add_2899_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n60047), 
            .O(n8605[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_3 (.CI(n60047), .I0(n2730), .I1(n858), .CO(n60048));
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4580));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2899_2_lut (.I0(n67890), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i63080_2_lut_4_lut (.I0(n77656), .I1(baudrate[6]), .I2(n1111), 
            .I3(n72246), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i63080_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY add_2899_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n60047));
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4581));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2898_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n60046), 
            .O(n8579[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4582));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8475[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2898_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n60045), 
            .O(n8579[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_18 (.CI(n60045), .I0(n2597), .I1(n2754), .CO(n60046));
    SB_LUT4 add_2898_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n60044), 
            .O(n8579[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8475[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2898_17 (.CI(n60044), .I0(n2598), .I1(n2638), .CO(n60045));
    SB_LUT4 i62878_3_lut_4_lut_3_lut (.I0(n72260), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n72264));
    defparam i62878_3_lut_4_lut_3_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2898_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n60043), 
            .O(n8579[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i56400_1_lut (.I0(n72246), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67932));
    defparam i56400_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2898_16 (.CI(n60043), .I0(n2599), .I1(n2519), .CO(n60044));
    SB_LUT4 add_2898_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n60042), 
            .O(n8579[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_15 (.CI(n60042), .I0(n2600), .I1(n2397), .CO(n60043));
    SB_LUT4 add_2898_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n60041), 
            .O(n8579[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8449[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8475[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2898_14 (.CI(n60041), .I0(n2601), .I1(n2272), .CO(n60042));
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4583));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2898_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n60040), 
            .O(n8579[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_13 (.CI(n60040), .I0(n2602), .I1(n2144), .CO(n60041));
    SB_LUT4 add_2898_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n60039), 
            .O(n8579[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_12 (.CI(n60039), .I0(n2603), .I1(n2013), .CO(n60040));
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8475[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n4_adj_4584));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4585));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8475[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4586));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2898_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n60038), 
            .O(n8579[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_11 (.CI(n60038), .I0(n2604), .I1(n1879), .CO(n60039));
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8475[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4587));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2898_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n60037), 
            .O(n8579[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_10 (.CI(n60037), .I0(n2605), .I1(n1742), .CO(n60038));
    SB_LUT4 add_2898_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n60036), 
            .O(n8579[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_9 (.CI(n60036), .I0(n2606), .I1(n1602), .CO(n60037));
    SB_LUT4 add_2898_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n60035), 
            .O(n8579[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_8 (.CI(n60035), .I0(n2607), .I1(n1459), .CO(n60036));
    SB_LUT4 add_2898_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n60034), 
            .O(n8579[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_7 (.CI(n60034), .I0(n2608), .I1(n1460), .CO(n60035));
    SB_LUT4 add_2898_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n60033), 
            .O(n8579[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_6 (.CI(n60033), .I0(n2609), .I1(n1011), .CO(n60034));
    SB_LUT4 add_2898_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n60032), 
            .O(n8579[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_5 (.CI(n60032), .I0(n2610), .I1(n856), .CO(n60033));
    SB_LUT4 add_2898_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n60031), 
            .O(n8579[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_4 (.CI(n60031), .I0(n2611), .I1(n698), .CO(n60032));
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8475[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2898_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n60030), 
            .O(n8579[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8475[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2898_3 (.CI(n60030), .I0(n2612), .I1(n858), .CO(n60031));
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8475[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4588));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2898_2_lut (.I0(n67894), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i56396_1_lut (.I0(n72242), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67924));
    defparam i56396_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2898_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n60030));
    SB_LUT4 add_2897_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n60029), 
            .O(n8553[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4589));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4590));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2897_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n60028), 
            .O(n8553[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8475[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2897_17 (.CI(n60028), .I0(n2477), .I1(n2638), .CO(n60029));
    SB_LUT4 add_2897_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n60027), 
            .O(n8553[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_16 (.CI(n60027), .I0(n2478), .I1(n2519), .CO(n60028));
    SB_LUT4 add_2897_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n60026), 
            .O(n8553[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_15 (.CI(n60026), .I0(n2479), .I1(n2397), .CO(n60027));
    SB_LUT4 add_2897_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n60025), 
            .O(n8553[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_14 (.CI(n60025), .I0(n2480), .I1(n2272), .CO(n60026));
    SB_LUT4 add_2897_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n60024), 
            .O(n8553[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_13 (.CI(n60024), .I0(n2481), .I1(n2144), .CO(n60025));
    SB_LUT4 add_2897_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n60023), 
            .O(n8553[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8475[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2897_12 (.CI(n60023), .I0(n2482), .I1(n2013), .CO(n60024));
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8475[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2897_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n60022), 
            .O(n8553[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_11 (.CI(n60022), .I0(n2483), .I1(n1879), .CO(n60023));
    SB_LUT4 add_2897_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n60021), 
            .O(n8553[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_10 (.CI(n60021), .I0(n2484), .I1(n1742), .CO(n60022));
    SB_LUT4 add_2897_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n60020), 
            .O(n8553[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_9 (.CI(n60020), .I0(n2485), .I1(n1602), .CO(n60021));
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4591));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4592));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2897_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n60019), 
            .O(n8553[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_8 (.CI(n60019), .I0(n2486), .I1(n1459), .CO(n60020));
    SB_LUT4 add_2897_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n60018), 
            .O(n8553[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_982 (.I0(n77656), .I1(baudrate[6]), .I2(n1111), 
            .I3(n70068), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_982.LUT_INIT = 16'h7100;
    SB_CARRY add_2897_7 (.CI(n60018), .I0(n2487), .I1(n1460), .CO(n60019));
    SB_LUT4 add_2897_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n60017), 
            .O(n8553[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_6 (.CI(n60017), .I0(n2488), .I1(n1011), .CO(n60018));
    SB_LUT4 add_2897_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n60016), 
            .O(n8553[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_5 (.CI(n60016), .I0(n2489), .I1(n856), .CO(n60017));
    SB_LUT4 add_2897_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n60015), 
            .O(n8553[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_4 (.CI(n60015), .I0(n2490), .I1(n698), .CO(n60016));
    SB_LUT4 add_2897_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n60014), 
            .O(n8553[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_3 (.CI(n60014), .I0(n2491), .I1(n858), .CO(n60015));
    SB_LUT4 add_2897_2_lut (.I0(n67898), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_4593));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4594));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2897_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n60014));
    SB_LUT4 add_2896_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n60013), 
            .O(n8527[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2896_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n60012), 
            .O(n8527[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8449[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2896_16 (.CI(n60012), .I0(n2354), .I1(n2519), .CO(n60013));
    SB_LUT4 add_2896_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n60011), 
            .O(n8527[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_15 (.CI(n60011), .I0(n2355), .I1(n2397), .CO(n60012));
    SB_LUT4 add_2896_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n60010), 
            .O(n8527[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_14 (.CI(n60010), .I0(n2356), .I1(n2272), .CO(n60011));
    SB_LUT4 add_2896_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n60009), 
            .O(n8527[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_13 (.CI(n60009), .I0(n2357), .I1(n2144), .CO(n60010));
    SB_LUT4 add_2896_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n60008), 
            .O(n8527[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_12 (.CI(n60008), .I0(n2358), .I1(n2013), .CO(n60009));
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8449[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2896_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n60007), 
            .O(n8527[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n59030), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_11 (.CI(n60007), .I0(n2359), .I1(n1879), .CO(n60008));
    SB_LUT4 add_2896_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n60006), 
            .O(n8527[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_10 (.CI(n60006), .I0(n2360), .I1(n1742), .CO(n60007));
    SB_LUT4 add_2896_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n60005), 
            .O(n8527[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i56382_1_lut (.I0(n72228), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67906));
    defparam i56382_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n70030), .I1(n294[23]), .I2(VCC_net), 
            .I3(n59029), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8449[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8449[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2896_9 (.CI(n60005), .I0(n2361), .I1(n1602), .CO(n60006));
    SB_CARRY sub_38_add_2_25 (.CI(n59029), .I0(n294[23]), .I1(VCC_net), 
            .CO(n59030));
    SB_LUT4 sub_38_add_2_24_lut (.I0(n70132), .I1(n72264), .I2(VCC_net), 
            .I3(n59028), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2896_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n60004), 
            .O(n8527[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4595));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_24 (.CI(n59028), .I0(n72264), .I1(VCC_net), 
            .CO(n59029));
    SB_CARRY add_2896_8 (.CI(n60004), .I0(n2362), .I1(n1459), .CO(n60005));
    SB_LUT4 add_2896_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n60003), 
            .O(n8527[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_7 (.CI(n60003), .I0(n2363), .I1(n1460), .CO(n60004));
    SB_LUT4 add_2896_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n60002), 
            .O(n8527[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_6 (.CI(n60002), .I0(n2364), .I1(n1011), .CO(n60003));
    SB_LUT4 add_2896_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n60001), 
            .O(n8527[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_5 (.CI(n60001), .I0(n2365), .I1(n856), .CO(n60002));
    SB_LUT4 add_2896_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n60000), 
            .O(n8527[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_4 (.CI(n60000), .I0(n2366), .I1(n698), .CO(n60001));
    SB_LUT4 add_2896_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n59999), 
            .O(n8527[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_3 (.CI(n59999), .I0(n2367), .I1(n858), .CO(n60000));
    SB_LUT4 add_2896_2_lut (.I0(n67902), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2896_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59999));
    SB_LUT4 add_2895_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n59998), 
            .O(n8501[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2895_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n59997), 
            .O(n8501[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_15 (.CI(n59997), .I0(n2228), .I1(n2397), .CO(n59998));
    SB_LUT4 add_2895_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n59996), 
            .O(n8501[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8449[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8449[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2895_14 (.CI(n59996), .I0(n2229), .I1(n2272), .CO(n59997));
    SB_LUT4 add_2895_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n59995), 
            .O(n8501[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8449[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2895_13 (.CI(n59995), .I0(n2230), .I1(n2144), .CO(n59996));
    SB_LUT4 add_2895_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n59994), 
            .O(n8501[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_12 (.CI(n59994), .I0(n2231), .I1(n2013), .CO(n59995));
    SB_LUT4 add_2895_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n59993), 
            .O(n8501[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_11 (.CI(n59993), .I0(n2232), .I1(n1879), .CO(n59994));
    SB_LUT4 add_2895_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n59992), 
            .O(n8501[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59654_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n75510));   // verilog/uart_rx.v(119[33:55])
    defparam i59654_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2895_10 (.CI(n59992), .I0(n2233), .I1(n1742), .CO(n59993));
    SB_LUT4 add_2895_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n59991), 
            .O(n8501[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_9 (.CI(n59991), .I0(n2234), .I1(n1602), .CO(n59992));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n59027), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2895_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n59990), 
            .O(n8501[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_8 (.CI(n59990), .I0(n2235), .I1(n1459), .CO(n59991));
    SB_LUT4 add_2895_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n59989), 
            .O(n8501[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_7 (.CI(n59989), .I0(n2236), .I1(n1460), .CO(n59990));
    SB_LUT4 add_2895_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n59988), 
            .O(n8501[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_6 (.CI(n59988), .I0(n2237), .I1(n1011), .CO(n59989));
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_23 (.CI(n59027), .I0(n294[21]), .I1(VCC_net), 
            .CO(n59028));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n70130), .I1(n294[20]), .I2(VCC_net), 
            .I3(n59026), .O(n70132)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2895_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n59987), 
            .O(n8501[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_5 (.CI(n59987), .I0(n2238), .I1(n856), .CO(n59988));
    SB_LUT4 add_2895_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n59986), 
            .O(n8501[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_4 (.CI(n59986), .I0(n2239), .I1(n698), .CO(n59987));
    SB_LUT4 add_2895_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n59985), 
            .O(n8501[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_3 (.CI(n59985), .I0(n2240), .I1(n858), .CO(n59986));
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8449[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2895_2_lut (.I0(n67906), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2895_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59985));
    SB_CARRY sub_38_add_2_22 (.CI(n59026), .I0(n294[20]), .I1(VCC_net), 
            .CO(n59027));
    SB_LUT4 add_2894_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n59984), 
            .O(n8475[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n70128), .I1(n294[19]), .I2(VCC_net), 
            .I3(n59025), .O(n70130)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2894_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n59983), 
            .O(n8475[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_13 (.CI(n59983), .I0(n2099), .I1(n2272), .CO(n59984));
    SB_LUT4 add_2894_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n59982), 
            .O(n8475[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_12 (.CI(n59982), .I0(n2100), .I1(n2144), .CO(n59983));
    SB_LUT4 add_2894_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n59981), 
            .O(n8475[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_11 (.CI(n59981), .I0(n2101), .I1(n2013), .CO(n59982));
    SB_LUT4 add_2894_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n59980), 
            .O(n8475[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_10 (.CI(n59980), .I0(n2102), .I1(n1879), .CO(n59981));
    SB_LUT4 add_2894_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n59979), 
            .O(n8475[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_983 (.I0(baudrate[3]), .I1(n42_adj_4599), 
            .I2(baudrate[4]), .I3(n21191), .O(n68354));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_983.LUT_INIT = 16'hff4f;
    SB_CARRY add_2894_9 (.CI(n59979), .I0(n2103), .I1(n1742), .CO(n59980));
    SB_LUT4 add_2894_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n59978), 
            .O(n8475[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_8 (.CI(n59978), .I0(n2104), .I1(n1602), .CO(n59979));
    SB_CARRY sub_38_add_2_21 (.CI(n59025), .I0(n294[19]), .I1(VCC_net), 
            .CO(n59026));
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n59024), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n59024), .I0(n294[18]), .I1(VCC_net), 
            .CO(n59025));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n70126), .I1(n294[17]), .I2(VCC_net), 
            .I3(n59023), .O(n70128)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2894_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n59977), 
            .O(n8475[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8449[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2894_7 (.CI(n59977), .I0(n2105), .I1(n1459), .CO(n59978));
    SB_LUT4 add_2894_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n59976), 
            .O(n8475[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_6 (.CI(n59976), .I0(n2106), .I1(n1460), .CO(n59977));
    SB_LUT4 add_2894_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n59975), 
            .O(n8475[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_5 (.CI(n59975), .I0(n2107), .I1(n1011), .CO(n59976));
    SB_LUT4 add_2894_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n59974), 
            .O(n8475[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_4 (.CI(n59974), .I0(n2108), .I1(n856), .CO(n59975));
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8449[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2894_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n59973), 
            .O(n8475[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_19 (.CI(n59023), .I0(n294[17]), .I1(VCC_net), 
            .CO(n59024));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n70124), .I1(n294[16]), .I2(VCC_net), 
            .I3(n59022), .O(n70126)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2894_3 (.CI(n59973), .I0(n2109), .I1(n698), .CO(n59974));
    SB_LUT4 add_2894_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8475[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2894_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n59973));
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_18 (.CI(n59022), .I0(n294[16]), .I1(VCC_net), 
            .CO(n59023));
    SB_LUT4 add_2893_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n59972), 
            .O(n8449[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2893_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n59971), 
            .O(n8449[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n70028), .I1(n294[15]), .I2(VCC_net), 
            .I3(n59021), .O(n70030)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8423[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2893_13 (.CI(n59971), .I0(n1967), .I1(n2144), .CO(n59972));
    SB_LUT4 add_2893_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n59970), 
            .O(n8449[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_12 (.CI(n59970), .I0(n1968), .I1(n2013), .CO(n59971));
    SB_LUT4 add_2893_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n59969), 
            .O(n8449[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_11 (.CI(n59969), .I0(n1969), .I1(n1879), .CO(n59970));
    SB_LUT4 add_2893_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n59968), 
            .O(n8449[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_17 (.CI(n59021), .I0(n294[15]), .I1(VCC_net), 
            .CO(n59022));
    SB_CARRY add_2893_10 (.CI(n59968), .I0(n1970), .I1(n1742), .CO(n59969));
    SB_LUT4 add_2893_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n59967), 
            .O(n8449[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_9 (.CI(n59967), .I0(n1971), .I1(n1602), .CO(n59968));
    SB_LUT4 add_2893_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n59966), 
            .O(n8449[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_16_lut (.I0(n70122), .I1(n294[14]), .I2(VCC_net), 
            .I3(n59020), .O(n70124)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_16 (.CI(n59020), .I0(n294[14]), .I1(VCC_net), 
            .CO(n59021));
    SB_CARRY add_2893_8 (.CI(n59966), .I0(n1972), .I1(n1459), .CO(n59967));
    SB_LUT4 add_2893_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n59965), 
            .O(n8449[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_7 (.CI(n59965), .I0(n1973), .I1(n1460), .CO(n59966));
    SB_LUT4 add_2893_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n59964), 
            .O(n8449[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_6 (.CI(n59964), .I0(n1974), .I1(n1011), .CO(n59965));
    SB_LUT4 add_2893_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n59963), 
            .O(n8449[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_5 (.CI(n59963), .I0(n1975), .I1(n856), .CO(n59964));
    SB_LUT4 add_2893_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n59962), 
            .O(n8449[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8423[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8423[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2893_4 (.CI(n59962), .I0(n1976), .I1(n698), .CO(n59963));
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n59019), .O(n70122)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2893_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n59961), 
            .O(n8449[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n59019), .I0(n294[13]), .I1(VCC_net), 
            .CO(n59020));
    SB_CARRY add_2893_3 (.CI(n59961), .I0(n1977), .I1(n858), .CO(n59962));
    SB_LUT4 add_2893_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8449[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59961));
    SB_LUT4 add_2892_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n59960), 
            .O(n8423[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2892_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n59959), 
            .O(n8423[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_12 (.CI(n59959), .I0(n1832), .I1(n2013), .CO(n59960));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n59018), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2892_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n59958), 
            .O(n8423[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_11 (.CI(n59958), .I0(n1833), .I1(n1879), .CO(n59959));
    SB_LUT4 add_2892_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n59957), 
            .O(n8423[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_14 (.CI(n59018), .I0(n294[12]), .I1(VCC_net), 
            .CO(n59019));
    SB_CARRY add_2892_10 (.CI(n59957), .I0(n1834), .I1(n1742), .CO(n59958));
    SB_LUT4 add_2892_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n59956), 
            .O(n8423[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_9 (.CI(n59956), .I0(n1835), .I1(n1602), .CO(n59957));
    SB_LUT4 add_2892_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n59955), 
            .O(n8423[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_8 (.CI(n59955), .I0(n1836), .I1(n1459), .CO(n59956));
    SB_LUT4 i52089_1_lut (.I0(n26019), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67898));
    defparam i52089_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2892_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n59954), 
            .O(n8423[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_7 (.CI(n59954), .I0(n1837), .I1(n1460), .CO(n59955));
    SB_LUT4 add_2892_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n59953), 
            .O(n8423[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59607_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n75463));   // verilog/uart_rx.v(119[33:55])
    defparam i59607_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2892_6 (.CI(n59953), .I0(n1838), .I1(n1011), .CO(n59954));
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8423[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2892_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n59952), 
            .O(n8423[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_5 (.CI(n59952), .I0(n1839), .I1(n856), .CO(n59953));
    SB_LUT4 add_2892_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n59951), 
            .O(n8423[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8423[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2892_4 (.CI(n59951), .I0(n1840), .I1(n698), .CO(n59952));
    SB_LUT4 add_2892_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n59950), 
            .O(n8423[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_3 (.CI(n59950), .I0(n1841), .I1(n858), .CO(n59951));
    SB_LUT4 add_2892_2_lut (.I0(n67915), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2892_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59950));
    SB_LUT4 add_2891_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n59949), 
            .O(n8397[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2891_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n59948), 
            .O(n8397[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_10 (.CI(n59948), .I0(n1694), .I1(n1879), .CO(n59949));
    SB_LUT4 add_2891_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n59947), 
            .O(n8397[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_9 (.CI(n59947), .I0(n1695), .I1(n1742), .CO(n59948));
    SB_LUT4 add_2891_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n59946), 
            .O(n8397[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n59017), .O(n70028)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2891_8 (.CI(n59946), .I0(n1696), .I1(n1602), .CO(n59947));
    SB_LUT4 add_2891_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n59945), 
            .O(n8397[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_7 (.CI(n59945), .I0(n1697), .I1(n1459), .CO(n59946));
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8423[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2891_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n59944), 
            .O(n8397[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_6 (.CI(n59944), .I0(n1698), .I1(n1460), .CO(n59945));
    SB_LUT4 add_2891_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n59943), 
            .O(n8397[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_5 (.CI(n59943), .I0(n1699), .I1(n1011), .CO(n59944));
    SB_LUT4 add_2891_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n59942), 
            .O(n8397[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_4 (.CI(n59942), .I0(n1700), .I1(n856), .CO(n59943));
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_13 (.CI(n59017), .I0(n294[11]), .I1(VCC_net), 
            .CO(n59018));
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n59016), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2891_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n59941), 
            .O(n8397[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8423[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2891_3 (.CI(n59941), .I0(n1701), .I1(n698), .CO(n59942));
    SB_LUT4 add_2891_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8397[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n59941));
    SB_LUT4 add_2890_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n59940), 
            .O(n8371[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2890_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n59939), 
            .O(n8371[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2890_10 (.CI(n59939), .I0(n1553), .I1(n1742), .CO(n59940));
    SB_LUT4 add_2890_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n59938), 
            .O(n8371[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_9 (.CI(n59938), .I0(n1554), .I1(n1602), .CO(n59939));
    SB_CARRY sub_38_add_2_12 (.CI(n59016), .I0(n294[10]), .I1(VCC_net), 
            .CO(n59017));
    SB_LUT4 add_2890_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n59937), 
            .O(n8371[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_4607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_2890_8 (.CI(n59937), .I0(n1555), .I1(n1459), .CO(n59938));
    SB_LUT4 add_2890_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n59936), 
            .O(n8371[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_7 (.CI(n59936), .I0(n1556), .I1(n1460), .CO(n59937));
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8423[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2890_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n59935), 
            .O(n8371[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_6 (.CI(n59935), .I0(n1557), .I1(n1011), .CO(n59936));
    SB_LUT4 add_2890_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n59934), 
            .O(n8371[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_5 (.CI(n59934), .I0(n1558), .I1(n856), .CO(n59935));
    SB_LUT4 add_2890_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n59933), 
            .O(n8371[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_4 (.CI(n59933), .I0(n1559), .I1(n698), .CO(n59934));
    SB_LUT4 add_2890_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n59932), 
            .O(n8371[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_3 (.CI(n59932), .I0(n1560), .I1(n858), .CO(n59933));
    SB_LUT4 add_2890_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8371[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59932));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n59015), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2889_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n59931), 
            .O(n8345[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2889_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n59930), 
            .O(n8345[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_9 (.CI(n59930), .I0(n1409), .I1(n1602), .CO(n59931));
    SB_LUT4 add_2889_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n59929), 
            .O(n8345[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8397[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2889_8 (.CI(n59929), .I0(n1410), .I1(n1459), .CO(n59930));
    SB_LUT4 add_2889_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n59928), 
            .O(n8345[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_7 (.CI(n59928), .I0(n1411), .I1(n1460), .CO(n59929));
    SB_LUT4 add_2889_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n59927), 
            .O(n8345[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_6 (.CI(n59927), .I0(n1412), .I1(n1011), .CO(n59928));
    SB_LUT4 add_2889_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n59926), 
            .O(n8345[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_5 (.CI(n59926), .I0(n1413), .I1(n856), .CO(n59927));
    SB_LUT4 add_2889_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n59925), 
            .O(n8345[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n59015), .I0(n294[9]), .I1(VCC_net), 
            .CO(n59016));
    SB_CARRY add_2889_4 (.CI(n59925), .I0(n1414), .I1(n698), .CO(n59926));
    SB_LUT4 add_2889_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n59924), 
            .O(n8345[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_3 (.CI(n59924), .I0(n1415), .I1(n858), .CO(n59925));
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8397[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8397[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2889_2_lut (.I0(n67924), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8397[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2889_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59924));
    SB_LUT4 add_2888_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n59923), 
            .O(n8319[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2888_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n59922), 
            .O(n8319[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_8 (.CI(n59922), .I0(n1262), .I1(n1459), .CO(n59923));
    SB_LUT4 add_2888_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n59921), 
            .O(n8319[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_7 (.CI(n59921), .I0(n1263), .I1(n1460), .CO(n59922));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n59014), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2888_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n59920), 
            .O(n8319[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_6 (.CI(n59920), .I0(n1264), .I1(n1011), .CO(n59921));
    SB_LUT4 add_2888_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n59919), 
            .O(n8319[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_10 (.CI(n59014), .I0(n294[8]), .I1(VCC_net), 
            .CO(n59015));
    SB_CARRY add_2888_5 (.CI(n59919), .I0(n1265), .I1(n856), .CO(n59920));
    SB_LUT4 add_2888_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n59918), 
            .O(n8319[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_4 (.CI(n59918), .I0(n1266), .I1(n698), .CO(n59919));
    SB_LUT4 add_2888_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n59917), 
            .O(n8319[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n59013), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_3 (.CI(n59917), .I0(n1267), .I1(n858), .CO(n59918));
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2888_2_lut (.I0(n67928), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2888_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59917));
    SB_LUT4 add_2887_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n59916), 
            .O(n8293[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2887_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n59915), 
            .O(n8293[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_7 (.CI(n59915), .I0(n1112), .I1(n1460), .CO(n59916));
    SB_LUT4 add_2887_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n59914), 
            .O(n8293[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_6 (.CI(n59914), .I0(n1113), .I1(n1011), .CO(n59915));
    SB_LUT4 add_2887_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n59913), 
            .O(n8293[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n59013), .I0(n294[7]), .I1(VCC_net), 
            .CO(n59014));
    SB_CARRY add_2887_5 (.CI(n59913), .I0(n1114), .I1(n856), .CO(n59914));
    SB_LUT4 add_2887_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n59912), 
            .O(n8293[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_4 (.CI(n59912), .I0(n1115), .I1(n698), .CO(n59913));
    SB_LUT4 add_2887_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n59911), 
            .O(n8293[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_3 (.CI(n59911), .I0(n1116), .I1(n858), .CO(n59912));
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n59012), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8397[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2887_2_lut (.I0(n67932), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n70068)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2887_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59911));
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8397[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_8 (.CI(n59012), .I0(n294[6]), .I1(VCC_net), 
            .CO(n59013));
    SB_LUT4 i1_3_lut_adj_984 (.I0(n26029), .I1(n48_adj_4611), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_984.LUT_INIT = 16'hefef;
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n59011), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n59011), .I0(n294[5]), .I1(VCC_net), 
            .CO(n59012));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n59010), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8397[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_6 (.CI(n59010), .I0(n294[4]), .I1(VCC_net), 
            .CO(n59011));
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4612));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n59009), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n59009), .I0(n294[3]), .I1(VCC_net), 
            .CO(n59010));
    SB_LUT4 i59590_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n75446));   // verilog/uart_rx.v(119[33:55])
    defparam i59590_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8397[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n8371[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_4613));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n8371[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n8371[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4614));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n8371[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n59008), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n59008), .I0(n294[2]), .I1(VCC_net), 
            .CO(n59009));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n59007), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n59007), .I0(n294[1]), .I1(VCC_net), 
            .CO(n59008));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n69091), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4615));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n69091), .I1(GND_net), 
            .CO(n59007));
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n8371[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4616));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n8371[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52065_1_lut_4_lut (.I0(n9_adj_4576), .I1(n14_adj_4577), .I2(n71486), 
            .I3(baudrate[30]), .O(n67874));
    defparam i52065_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4617));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n8371[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n8371[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_985 (.I0(n71472), .I1(n71488), .I2(n71486), .I3(baudrate[11]), 
            .O(n71416));
    defparam i1_4_lut_adj_985.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_986 (.I0(n71418), .I1(n70620), .I2(n71416), .I3(GND_net), 
            .O(n26029));
    defparam i1_3_lut_adj_986.LUT_INIT = 16'hfefe;
    SB_LUT4 i30793_rep_5_2_lut (.I0(n8371[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n67918));   // verilog/uart_rx.v(119[33:55])
    defparam i30793_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n67918), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_4618));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i62050_3_lut (.I0(n32_adj_4618), .I1(baudrate[6]), .I2(n39_adj_4617), 
            .I3(GND_net), .O(n77906));   // verilog/uart_rx.v(119[33:55])
    defparam i62050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62051_3_lut (.I0(n77906), .I1(baudrate[7]), .I2(n41_adj_4616), 
            .I3(GND_net), .O(n77907));   // verilog/uart_rx.v(119[33:55])
    defparam i62051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60536_4_lut (.I0(n41_adj_4616), .I1(n39_adj_4617), .I2(n37_adj_4615), 
            .I3(n75446), .O(n76392));
    defparam i60536_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i62455_2_lut_3_lut_4_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n28240));
    defparam i62455_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i61391_3_lut (.I0(n34_adj_4613), .I1(baudrate[5]), .I2(n37_adj_4615), 
            .I3(GND_net), .O(n77247));   // verilog/uart_rx.v(119[33:55])
    defparam i61391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61776_3_lut (.I0(n77907), .I1(baudrate[8]), .I2(n43_adj_4614), 
            .I3(GND_net), .O(n77632));   // verilog/uart_rx.v(119[33:55])
    defparam i61776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62048_4_lut (.I0(n77632), .I1(n77247), .I2(n43_adj_4614), 
            .I3(n76392), .O(n77904));   // verilog/uart_rx.v(119[33:55])
    defparam i62048_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62049_3_lut (.I0(n77904), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n77905));   // verilog/uart_rx.v(119[33:55])
    defparam i62049_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61778_3_lut (.I0(n77905), .I1(baudrate[10]), .I2(n1693), 
            .I3(GND_net), .O(n48_adj_4611));   // verilog/uart_rx.v(119[33:55])
    defparam i61778_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n8345[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n8345[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n8345[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_987 (.I0(n71358), .I1(baudrate[18]), 
            .I2(baudrate[19]), .I3(n71472), .O(n71364));
    defparam i1_2_lut_3_lut_4_lut_adj_987.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4619));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n8345[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4620));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n8345[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4621));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n8345[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4622));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n8345[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52081_1_lut (.I0(n25967), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67890));
    defparam i52081_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_4623));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_988 (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n70588), .I3(n71362), .O(n70602));
    defparam i1_3_lut_4_lut_adj_988.LUT_INIT = 16'hfffe;
    SB_LUT4 i61789_3_lut (.I0(n32_adj_4623), .I1(baudrate[5]), .I2(n39_adj_4622), 
            .I3(GND_net), .O(n77645));   // verilog/uart_rx.v(119[33:55])
    defparam i61789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61790_3_lut (.I0(n77645), .I1(baudrate[6]), .I2(n41_adj_4621), 
            .I3(GND_net), .O(n77646));   // verilog/uart_rx.v(119[33:55])
    defparam i61790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60552_4_lut (.I0(n41_adj_4621), .I1(n39_adj_4622), .I2(n37_adj_4620), 
            .I3(n75463), .O(n76408));
    defparam i60552_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61389_3_lut (.I0(n34_adj_4607), .I1(baudrate[4]), .I2(n37_adj_4620), 
            .I3(GND_net), .O(n77245));   // verilog/uart_rx.v(119[33:55])
    defparam i61389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61772_3_lut (.I0(n77646), .I1(baudrate[7]), .I2(n43_adj_4619), 
            .I3(GND_net), .O(n77628));   // verilog/uart_rx.v(119[33:55])
    defparam i61772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61783_4_lut (.I0(n77628), .I1(n77245), .I2(n43_adj_4619), 
            .I3(n76408), .O(n77639));   // verilog/uart_rx.v(119[33:55])
    defparam i61783_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61784_3_lut (.I0(n77639), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n77640));   // verilog/uart_rx.v(119[33:55])
    defparam i61784_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61774_3_lut (.I0(n77640), .I1(baudrate[9]), .I2(n1552), .I3(GND_net), 
            .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i61774_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n8319[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n8319[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4624));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n8319[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4625));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n8319[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_989 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[15]), .I3(baudrate[14]), .O(n70654));
    defparam i1_2_lut_3_lut_4_lut_adj_989.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4626));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n8319[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4627));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_990 (.I0(n70070), .I1(n48_adj_4507), .I2(GND_net), 
            .I3(GND_net), .O(n1415));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n8293[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n8293[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n8293[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n8293[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4628));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5844_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n68354), .I3(n44_adj_4629), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i5844_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i742_4_lut (.I0(n67645), .I1(n294[18]), .I2(n46), .I3(baudrate[5]), 
            .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 i7317_4_lut (.I0(n960), .I1(n11692), .I2(n21189), .I3(baudrate[3]), 
            .O(n21191));   // verilog/uart_rx.v(119[33:55])
    defparam i7317_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_4629), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_4630), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i5822_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_4630));   // verilog/uart_rx.v(119[33:55])
    defparam i5822_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i7316_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n21189));   // verilog/uart_rx.v(119[33:55])
    defparam i7316_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i5830_2_lut (.I0(n21189), .I1(n11692), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_4599));   // verilog/uart_rx.v(119[33:55])
    defparam i5830_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_4599), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4631));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_991 (.I0(n26035), .I1(n48_adj_4632), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_991.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_4633));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_4593), .I1(baudrate[4]), 
            .I2(n43_adj_4631), .I3(GND_net), .O(n42_adj_4634));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61799_4_lut (.I0(n42_adj_4634), .I1(n38_adj_4633), .I2(n43_adj_4631), 
            .I3(n75510), .O(n77655));   // verilog/uart_rx.v(119[33:55])
    defparam i61799_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61800_3_lut (.I0(n77655), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n77656));   // verilog/uart_rx.v(119[33:55])
    defparam i61800_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5673_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n68370), .I3(n44_adj_4635), 
            .O(n46_adj_4636));   // verilog/uart_rx.v(119[33:55])
    defparam i5673_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i639_4_lut (.I0(n67643), .I1(n294[19]), .I2(n46_adj_4636), 
            .I3(baudrate[4]), .O(n67645));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 r_Clock_Count_2053_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n60289), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n60288), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_8 (.CI(n60288), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n60289));
    SB_LUT4 r_Clock_Count_2053_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n60287), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7310_4_lut (.I0(n804), .I1(n44852), .I2(n21179), .I3(baudrate[2]), 
            .O(n21181));   // verilog/uart_rx.v(119[33:55])
    defparam i7310_4_lut.LUT_INIT = 16'ha2aa;
    SB_CARRY r_Clock_Count_2053_add_4_7 (.CI(n60287), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n60288));
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_4635), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 r_Clock_Count_2053_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n60286), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52077_1_lut (.I0(n25970), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67886));
    defparam i52077_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_4578), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i1_4_lut_adj_992 (.I0(n25991), .I1(n48_adj_4637), .I2(n44854), 
            .I3(baudrate[2]), .O(n68378));
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hefff;
    SB_LUT4 i5504_4_lut (.I0(n644), .I1(baudrate[2]), .I2(n68378), .I3(n44_adj_4638), 
            .O(n46_adj_4639));   // verilog/uart_rx.v(119[33:55])
    defparam i5504_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i534_4_lut (.I0(n67641), .I1(n294[20]), .I2(n46_adj_4639), 
            .I3(baudrate[3]), .O(n67643));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 i60377_4_lut (.I0(n25991), .I1(n75551), .I2(n48_adj_4637), 
            .I3(baudrate[0]), .O(n804));
    defparam i60377_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i1_2_lut_4_lut_adj_993 (.I0(n78107), .I1(baudrate[18]), .I2(n2713), 
            .I3(n70084), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_993.LUT_INIT = 16'h7100;
    SB_LUT4 i62613_2_lut (.I0(n48_adj_4640), .I1(n26022), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i62613_2_lut.LUT_INIT = 16'h1111;
    SB_CARRY r_Clock_Count_2053_add_4_6 (.CI(n60286), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n60287));
    SB_LUT4 i63220_2_lut_4_lut (.I0(n78107), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25967), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i63220_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i535_4_lut (.I0(n644), .I1(n44_adj_4638), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_3_lut_adj_994 (.I0(n25988), .I1(n48_adj_4641), .I2(n44854), 
            .I3(GND_net), .O(n68402));
    defparam i1_3_lut_adj_994.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i427_4_lut (.I0(n5), .I1(n68402), .I2(n294[21]), .I3(baudrate[2]), 
            .O(n67641));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_4_lut_adj_995 (.I0(n70620), .I1(n71478), .I2(n71468), .I3(baudrate[19]), 
            .O(n25967));
    defparam i1_4_lut_adj_995.LUT_INIT = 16'hfffe;
    SB_LUT4 i63237_2_lut (.I0(n48_adj_4637), .I1(n25991), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i63237_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i62841_2_lut (.I0(baudrate[1]), .I1(n72260), .I2(GND_net), 
            .I3(GND_net), .O(n294[23]));
    defparam i62841_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i56355_4_lut (.I0(baudrate[1]), .I1(n71362), .I2(n70588), 
            .I3(baudrate[3]), .O(n72202));
    defparam i56355_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_996 (.I0(n72202), .I1(n72228), .I2(n71360), .I3(n70512), 
            .O(n48_adj_4641));
    defparam i1_4_lut_adj_996.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_997 (.I0(n70602), .I1(n25937), .I2(n71360), .I3(n71358), 
            .O(n25988));
    defparam i1_4_lut_adj_997.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_998 (.I0(baudrate[23]), .I1(baudrate[1]), .I2(GND_net), 
            .I3(GND_net), .O(n70444));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'h4444;
    SB_LUT4 i56359_4_lut (.I0(baudrate[19]), .I1(n70588), .I2(baudrate[3]), 
            .I3(baudrate[20]), .O(n72206));
    defparam i56359_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i56343_3_lut (.I0(baudrate[21]), .I1(baudrate[10]), .I2(baudrate[22]), 
            .I3(GND_net), .O(n72190));
    defparam i56343_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_999 (.I0(n72184), .I1(n72116), .I2(n71470), .I3(n70444), 
            .O(n70486));
    defparam i1_4_lut_adj_999.LUT_INIT = 16'h0100;
    SB_LUT4 i56369_4_lut (.I0(n14_adj_4577), .I1(n72206), .I2(n72118), 
            .I3(baudrate[2]), .O(n72216));
    defparam i56369_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i56371_4_lut (.I0(n9_adj_4576), .I1(n71352), .I2(n71354), 
            .I3(n72190), .O(n72218));
    defparam i56371_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1000 (.I0(n45376), .I1(n72218), .I2(n72216), 
            .I3(n70486), .O(n5));   // verilog/uart_rx.v(119[33:55])
    defparam i1_4_lut_adj_1000.LUT_INIT = 16'habaa;
    SB_LUT4 div_37_LessThan_341_i48_4_lut (.I0(n72260), .I1(baudrate[2]), 
            .I2(n5), .I3(n44854), .O(n48_adj_4637));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_4_lut.LUT_INIT = 16'hd4c0;
    SB_LUT4 i60380_4_lut (.I0(n25988), .I1(n75548), .I2(n48_adj_4641), 
            .I3(baudrate[0]), .O(n644));
    defparam i60380_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i56271_2_lut (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n72118));
    defparam i56271_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i30765_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44854));
    defparam i30765_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(baudrate[7]), .I1(baudrate[9]), .I2(baudrate[8]), 
            .I3(baudrate[10]), .O(n70552));
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1002 (.I0(n72184), .I1(n72116), .I2(n72118), 
            .I3(GND_net), .O(n70556));
    defparam i1_3_lut_adj_1002.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1003 (.I0(n70554), .I1(n25967), .I2(n70556), 
            .I3(n70552), .O(n25991));
    defparam i1_4_lut_adj_1003.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n75234), .I1(baudrate[2]), 
            .I2(n644), .I3(n48_adj_4637), .O(n46_adj_4642));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_4642), .I1(baudrate[3]), 
            .I2(n67641), .I3(GND_net), .O(n48_adj_4640));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_3_lut_adj_1004 (.I0(n70662), .I1(n25970), .I2(n71418), 
            .I3(GND_net), .O(n26022));
    defparam i1_3_lut_adj_1004.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1005 (.I0(n26022), .I1(n48_adj_4640), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1005.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_4643));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61810_3_lut (.I0(n42_adj_4643), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n77666));   // verilog/uart_rx.v(119[33:55])
    defparam i61810_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61811_3_lut (.I0(n77666), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n77667));   // verilog/uart_rx.v(119[33:55])
    defparam i61811_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61760_3_lut (.I0(n77667), .I1(baudrate[4]), .I2(n67643), 
            .I3(GND_net), .O(n48_adj_4644));   // verilog/uart_rx.v(119[33:55])
    defparam i61760_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(n71362), .I1(n25976), .I2(n71364), 
            .I3(n71360), .O(n26035));
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'hfffe;
    SB_LUT4 i30770_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n67935));   // verilog/uart_rx.v(119[33:55])
    defparam i30770_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n67935), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_4645));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61806_3_lut (.I0(n42_adj_4645), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n77662));   // verilog/uart_rx.v(119[33:55])
    defparam i61806_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61807_3_lut (.I0(n77662), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n77663));   // verilog/uart_rx.v(119[33:55])
    defparam i61807_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1007 (.I0(n77885), .I1(baudrate[21]), .I2(n3046), 
            .I3(n70090), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1007.LUT_INIT = 16'h7100;
    SB_LUT4 i61762_3_lut (.I0(n77663), .I1(baudrate[5]), .I2(n67645), 
            .I3(GND_net), .O(n48_adj_4632));   // verilog/uart_rx.v(119[33:55])
    defparam i61762_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i63240_2_lut_4_lut (.I0(n77885), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25976), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i63240_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_adj_1008 (.I0(n72256), .I1(n48_adj_4644), .I2(baudrate[0]), 
            .I3(GND_net), .O(n962));
    defparam i1_3_lut_adj_1008.LUT_INIT = 16'h1010;
    SB_LUT4 i60368_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i60368_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n8293[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_4646));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_4543), .I1(baudrate[4]), 
            .I2(n41_adj_4628), .I3(GND_net), .O(n40_adj_4647));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62297_4_lut (.I0(n40_adj_4647), .I1(n36_adj_4646), .I2(n41_adj_4628), 
            .I3(n75495), .O(n78153));   // verilog/uart_rx.v(119[33:55])
    defparam i62297_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62298_3_lut (.I0(n78153), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n78154));   // verilog/uart_rx.v(119[33:55])
    defparam i62298_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_4648));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62234_3_lut (.I0(n78154), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n78090));   // verilog/uart_rx.v(119[33:55])
    defparam i62234_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62039_3_lut (.I0(n78090), .I1(baudrate[7]), .I2(n1261), .I3(GND_net), 
            .O(n48_adj_4507));   // verilog/uart_rx.v(119[33:55])
    defparam i62039_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60138_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n75994));
    defparam i60138_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_4649));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n8293[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n8319[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62040_3_lut (.I0(n34_adj_4650), .I1(baudrate[5]), .I2(n41_adj_4627), 
            .I3(GND_net), .O(n77896));   // verilog/uart_rx.v(119[33:55])
    defparam i62040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62041_3_lut (.I0(n77896), .I1(baudrate[6]), .I2(n43_adj_4626), 
            .I3(GND_net), .O(n77897));   // verilog/uart_rx.v(119[33:55])
    defparam i62041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60558_4_lut (.I0(n43_adj_4626), .I1(n41_adj_4627), .I2(n39_adj_4625), 
            .I3(n75472), .O(n76414));
    defparam i60558_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36), .I1(baudrate[4]), .I2(n39_adj_4625), 
            .I3(GND_net), .O(n38_adj_4651));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61768_3_lut (.I0(n77897), .I1(baudrate[7]), .I2(n45_adj_4624), 
            .I3(GND_net), .O(n44_adj_4652));   // verilog/uart_rx.v(119[33:55])
    defparam i61768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61387_4_lut (.I0(n44_adj_4652), .I1(n38_adj_4651), .I2(n45_adj_4624), 
            .I3(n76414), .O(n77243));   // verilog/uart_rx.v(119[33:55])
    defparam i61387_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_4653));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60112_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n75968));
    defparam i60112_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n8319[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_4654));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n8345[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n8371[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8397[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4655));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60213_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5217), .I3(\o_Rx_DV_N_3488[8] ), .O(n75205));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i60213_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4656));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4657));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60345_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n66553), 
            .I3(r_SM_Main[0]), .O(n75211));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i60345_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i60208_4_lut (.I0(n75205), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n75202));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i60208_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i56385_2_lut (.I0(baudrate[12]), .I1(n72230), .I2(GND_net), 
            .I3(GND_net), .O(n72232));
    defparam i56385_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4658));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60218_4_lut (.I0(n75211), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n75208));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i60218_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i59572_4_lut (.I0(n35_adj_4657), .I1(n33_adj_4656), .I2(n31_adj_4655), 
            .I3(n29_adj_4658), .O(n75428));
    defparam i59572_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n75208), .I1(n75202), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_4548));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_4659), .I1(baudrate[9]), 
            .I2(n43_adj_4610), .I3(GND_net), .O(n40_adj_4660));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_4661));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62044_3_lut (.I0(n28_adj_4661), .I1(baudrate[5]), .I2(n35_adj_4657), 
            .I3(GND_net), .O(n77900));   // verilog/uart_rx.v(119[33:55])
    defparam i62044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62045_3_lut (.I0(n77900), .I1(baudrate[6]), .I2(n37_adj_4609), 
            .I3(GND_net), .O(n77901));   // verilog/uart_rx.v(119[33:55])
    defparam i62045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59566_4_lut (.I0(n41_adj_4612), .I1(n39_adj_4608), .I2(n37_adj_4609), 
            .I3(n75428), .O(n75422));
    defparam i59566_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62042_4_lut (.I0(n40_adj_4660), .I1(n30_adj_4662), .I2(n43_adj_4610), 
            .I3(n75416), .O(n77898));   // verilog/uart_rx.v(119[33:55])
    defparam i62042_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61780_3_lut (.I0(n77901), .I1(baudrate[7]), .I2(n39_adj_4608), 
            .I3(GND_net), .O(n77636));   // verilog/uart_rx.v(119[33:55])
    defparam i61780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62316_4_lut (.I0(n77636), .I1(n77898), .I2(n43_adj_4610), 
            .I3(n75422), .O(n78172));   // verilog/uart_rx.v(119[33:55])
    defparam i62316_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62317_3_lut (.I0(n78172), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n78173));   // verilog/uart_rx.v(119[33:55])
    defparam i62317_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_1009 (.I0(baudrate[31]), .I1(baudrate[23]), 
            .I2(baudrate[21]), .I3(GND_net), .O(n71490));
    defparam i1_2_lut_3_lut_adj_1009.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1010 (.I0(n71438), .I1(baudrate[22]), 
            .I2(baudrate[23]), .I3(n71470), .O(n71442));
    defparam i1_2_lut_3_lut_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8397[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8423[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8423[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4663));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4664));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4665));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4666));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59530_4_lut (.I0(n33_adj_4665), .I1(n31_adj_4664), .I2(n29_adj_4663), 
            .I3(n27_adj_4666), .O(n75386));
    defparam i59530_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_4667), .I1(baudrate[9]), 
            .I2(n41_adj_4603), .I3(GND_net), .O(n38_adj_4668));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_4669));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62036_3_lut (.I0(n26_adj_4669), .I1(baudrate[5]), .I2(n33_adj_4665), 
            .I3(GND_net), .O(n77892));   // verilog/uart_rx.v(119[33:55])
    defparam i62036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62037_3_lut (.I0(n77892), .I1(baudrate[6]), .I2(n35_adj_4605), 
            .I3(GND_net), .O(n77893));   // verilog/uart_rx.v(119[33:55])
    defparam i62037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59526_4_lut (.I0(n39_adj_4606), .I1(n37_adj_4604), .I2(n35_adj_4605), 
            .I3(n75386), .O(n75382));
    defparam i59526_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62299_4_lut (.I0(n38_adj_4668), .I1(n28_adj_4670), .I2(n41_adj_4603), 
            .I3(n75379), .O(n78155));   // verilog/uart_rx.v(119[33:55])
    defparam i62299_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61786_3_lut (.I0(n77893), .I1(baudrate[7]), .I2(n37_adj_4604), 
            .I3(GND_net), .O(n77642));   // verilog/uart_rx.v(119[33:55])
    defparam i61786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62397_4_lut (.I0(n77642), .I1(n78155), .I2(n41_adj_4603), 
            .I3(n75382), .O(n78253));   // verilog/uart_rx.v(119[33:55])
    defparam i62397_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62398_3_lut (.I0(n78253), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n78254));   // verilog/uart_rx.v(119[33:55])
    defparam i62398_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62372_3_lut (.I0(n78254), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n78228));   // verilog/uart_rx.v(119[33:55])
    defparam i62372_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62321_3_lut (.I0(n78228), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_4671));   // verilog/uart_rx.v(119[33:55])
    defparam i62321_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8423[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8449[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(n71442), .I1(n9_adj_4576), .I2(n14_adj_4577), 
            .I3(n71358), .O(n26010));
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4672));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59512_4_lut (.I0(n33_adj_4602), .I1(n31_adj_4601), .I2(n29_adj_4600), 
            .I3(n27_adj_4672), .O(n75368));
    defparam i59512_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_4673), .I1(baudrate[10]), 
            .I2(n41_adj_4597), .I3(GND_net), .O(n38_adj_4674));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30802_rep_4_2_lut (.I0(n8449[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n67909));   // verilog/uart_rx.v(119[33:55])
    defparam i30802_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n67909), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_4675));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i62032_3_lut (.I0(n26_adj_4675), .I1(baudrate[6]), .I2(n33_adj_4602), 
            .I3(GND_net), .O(n77888));   // verilog/uart_rx.v(119[33:55])
    defparam i62032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62033_3_lut (.I0(n77888), .I1(baudrate[7]), .I2(n35_adj_4595), 
            .I3(GND_net), .O(n77889));   // verilog/uart_rx.v(119[33:55])
    defparam i62033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59506_4_lut (.I0(n39_adj_4598), .I1(n37_adj_4596), .I2(n35_adj_4595), 
            .I3(n75368), .O(n75362));
    defparam i59506_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62303_4_lut (.I0(n38_adj_4674), .I1(n28_adj_4676), .I2(n41_adj_4597), 
            .I3(n75359), .O(n78159));   // verilog/uart_rx.v(119[33:55])
    defparam i62303_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61792_3_lut (.I0(n77889), .I1(baudrate[8]), .I2(n37_adj_4596), 
            .I3(GND_net), .O(n77648));   // verilog/uart_rx.v(119[33:55])
    defparam i61792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62399_4_lut (.I0(n77648), .I1(n78159), .I2(n41_adj_4597), 
            .I3(n75362), .O(n78255));   // verilog/uart_rx.v(119[33:55])
    defparam i62399_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62400_3_lut (.I0(n78255), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n78256));   // verilog/uart_rx.v(119[33:55])
    defparam i62400_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62370_3_lut (.I0(n78256), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n78226));   // verilog/uart_rx.v(119[33:55])
    defparam i62370_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62323_3_lut (.I0(n78226), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_4677));   // verilog/uart_rx.v(119[33:55])
    defparam i62323_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1012 (.I0(n72230), .I1(n48_adj_4671), .I2(n8449[11]), 
            .I3(GND_net), .O(n2110));
    defparam i1_3_lut_adj_1012.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8475[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56269_2_lut (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n72116));
    defparam i56269_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i56377_4_lut (.I0(n71486), .I1(n9_adj_4576), .I2(n71474), 
            .I3(baudrate[17]), .O(n72224));
    defparam i56377_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i56381_4_lut (.I0(n72196), .I1(n72224), .I2(n14_adj_4577), 
            .I3(n72116), .O(n72228));
    defparam i56381_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4678));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59492_4_lut (.I0(n29_adj_4594), .I1(n27_adj_4592), .I2(n25_adj_4591), 
            .I3(n23_adj_4678), .O(n75348));
    defparam i59492_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59488_4_lut (.I0(n35_adj_4590), .I1(n33_adj_4589), .I2(n31_adj_4588), 
            .I3(n75348), .O(n75344));
    defparam i59488_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_4679));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_4680), .I1(baudrate[7]), 
            .I2(n33_adj_4589), .I3(GND_net), .O(n30_adj_4681));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_4682), .I1(baudrate[9]), 
            .I2(n37_adj_4587), .I3(GND_net), .O(n34_adj_4683));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62217_4_lut (.I0(n34_adj_4683), .I1(n24_adj_4684), .I2(n37_adj_4587), 
            .I3(n75338), .O(n78073));   // verilog/uart_rx.v(119[33:55])
    defparam i62217_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62218_3_lut (.I0(n78073), .I1(baudrate[10]), .I2(n39_adj_4586), 
            .I3(GND_net), .O(n78074));   // verilog/uart_rx.v(119[33:55])
    defparam i62218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62069_3_lut (.I0(n78074), .I1(baudrate[11]), .I2(n41_adj_4585), 
            .I3(GND_net), .O(n77925));   // verilog/uart_rx.v(119[33:55])
    defparam i62069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61665_4_lut (.I0(n41_adj_4585), .I1(n39_adj_4586), .I2(n37_adj_4587), 
            .I3(n75344), .O(n77521));
    defparam i61665_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62225_4_lut (.I0(n30_adj_4681), .I1(n22_adj_4679), .I2(n33_adj_4589), 
            .I3(n75346), .O(n78081));   // verilog/uart_rx.v(119[33:55])
    defparam i62225_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60727_3_lut (.I0(n77925), .I1(baudrate[12]), .I2(n43_adj_4583), 
            .I3(GND_net), .O(n76583));   // verilog/uart_rx.v(119[33:55])
    defparam i60727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62309_4_lut (.I0(n76583), .I1(n78081), .I2(n43_adj_4583), 
            .I3(n77521), .O(n78165));   // verilog/uart_rx.v(119[33:55])
    defparam i62309_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62310_3_lut (.I0(n78165), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n78166));   // verilog/uart_rx.v(119[33:55])
    defparam i62310_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1013 (.I0(n26010), .I1(n48_adj_4677), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1013.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8501[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_4685));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(n14_adj_4577), .I1(n9_adj_4576), .I2(n71462), 
            .I3(n71438), .O(n26016));
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4686));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60437_4_lut (.I0(n27_adj_4582), .I1(n25_adj_4581), .I2(n23_adj_4580), 
            .I3(n21_adj_4686), .O(n76293));
    defparam i60437_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60429_4_lut (.I0(n33_adj_4575), .I1(n31_adj_4574), .I2(n29_adj_4573), 
            .I3(n76293), .O(n76285));
    defparam i60429_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_4687));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_4688), .I1(baudrate[7]), 
            .I2(n31_adj_4574), .I3(GND_net), .O(n28_adj_4689));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_4690), .I1(baudrate[9]), 
            .I2(n35_adj_4572), .I3(GND_net), .O(n32_adj_4691));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62219_4_lut (.I0(n32_adj_4691), .I1(n22_adj_4692), .I2(n35_adj_4572), 
            .I3(n76283), .O(n78075));   // verilog/uart_rx.v(119[33:55])
    defparam i62219_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62220_3_lut (.I0(n78075), .I1(baudrate[10]), .I2(n37_adj_4566), 
            .I3(GND_net), .O(n78076));   // verilog/uart_rx.v(119[33:55])
    defparam i62220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62067_3_lut (.I0(n78076), .I1(baudrate[11]), .I2(n39_adj_4571), 
            .I3(GND_net), .O(n77923));   // verilog/uart_rx.v(119[33:55])
    defparam i62067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61957_4_lut (.I0(n39_adj_4571), .I1(n37_adj_4566), .I2(n35_adj_4572), 
            .I3(n76285), .O(n77813));
    defparam i61957_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62221_4_lut (.I0(n28_adj_4689), .I1(n20_adj_4687), .I2(n31_adj_4574), 
            .I3(n76289), .O(n78077));   // verilog/uart_rx.v(119[33:55])
    defparam i62221_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60731_3_lut (.I0(n77923), .I1(baudrate[12]), .I2(n41_adj_4564), 
            .I3(GND_net), .O(n76587));   // verilog/uart_rx.v(119[33:55])
    defparam i60731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62293_4_lut (.I0(n76587), .I1(n78077), .I2(n41_adj_4564), 
            .I3(n77813), .O(n78149));   // verilog/uart_rx.v(119[33:55])
    defparam i62293_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62294_3_lut (.I0(n78149), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n78150));   // verilog/uart_rx.v(119[33:55])
    defparam i62294_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62257_3_lut (.I0(n78150), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n78113));   // verilog/uart_rx.v(119[33:55])
    defparam i62257_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60198_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n76054));
    defparam i60198_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_4693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_4694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8527[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60383_4_lut (.I0(n25_adj_4695), .I1(n23_adj_4547), .I2(n21_adj_4546), 
            .I3(n19_adj_4697), .O(n76239));
    defparam i60383_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60371_4_lut (.I0(n31_adj_4545), .I1(n29_adj_4544), .I2(n27_adj_4696), 
            .I3(n76239), .O(n76227));
    defparam i60371_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60166_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n76022));
    defparam i60166_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i61951_4_lut (.I0(n37_adj_4541), .I1(n35_adj_4540), .I2(n33_adj_4539), 
            .I3(n76227), .O(n77807));
    defparam i61951_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2491), .I3(GND_net), .O(n18_adj_4698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61757_3_lut (.I0(n18_adj_4698), .I1(baudrate[13]), .I2(n41_adj_4537), 
            .I3(GND_net), .O(n77613));   // verilog/uart_rx.v(119[33:55])
    defparam i61757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61758_3_lut (.I0(n77613), .I1(baudrate[14]), .I2(n43_adj_4535), 
            .I3(GND_net), .O(n77614));   // verilog/uart_rx.v(119[33:55])
    defparam i61758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61229_4_lut (.I0(n43_adj_4535), .I1(n41_adj_4537), .I2(n29_adj_4544), 
            .I3(n76234), .O(n77085));
    defparam i61229_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_4699), .I1(baudrate[7]), 
            .I2(n29_adj_4544), .I3(GND_net), .O(n26_adj_4700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60743_3_lut (.I0(n77614), .I1(baudrate[15]), .I2(n45_adj_4532), 
            .I3(GND_net), .O(n76599));   // verilog/uart_rx.v(119[33:55])
    defparam i60743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_4701), .I1(baudrate[9]), 
            .I2(n33_adj_4539), .I3(GND_net), .O(n30_adj_4702));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62231_4_lut (.I0(n30_adj_4702), .I1(n20_adj_4703), .I2(n33_adj_4539), 
            .I3(n76215), .O(n78087));   // verilog/uart_rx.v(119[33:55])
    defparam i62231_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62232_3_lut (.I0(n78087), .I1(baudrate[10]), .I2(n35_adj_4540), 
            .I3(GND_net), .O(n78088));   // verilog/uart_rx.v(119[33:55])
    defparam i62232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62047_3_lut (.I0(n78088), .I1(baudrate[11]), .I2(n37_adj_4541), 
            .I3(GND_net), .O(n77903));   // verilog/uart_rx.v(119[33:55])
    defparam i62047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61231_4_lut (.I0(n43_adj_4535), .I1(n41_adj_4537), .I2(n39_adj_4526), 
            .I3(n77807), .O(n77087));
    defparam i61231_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61801_4_lut (.I0(n76599), .I1(n26_adj_4700), .I2(n45_adj_4532), 
            .I3(n77085), .O(n77657));   // verilog/uart_rx.v(119[33:55])
    defparam i61801_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60741_3_lut (.I0(n77903), .I1(baudrate[12]), .I2(n39_adj_4526), 
            .I3(GND_net), .O(n76597));   // verilog/uart_rx.v(119[33:55])
    defparam i60741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61803_4_lut (.I0(n76597), .I1(n77657), .I2(n45_adj_4532), 
            .I3(n77087), .O(n77659));   // verilog/uart_rx.v(119[33:55])
    defparam i61803_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_4704));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8527[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8553[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8553[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4705));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4706));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(n70620), .I1(n71442), .I2(GND_net), 
            .I3(GND_net), .O(n25937));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4707));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60319_4_lut (.I0(n23_adj_4705), .I1(n21_adj_4520), .I2(n19_adj_4514), 
            .I3(n17_adj_4707), .O(n76175));
    defparam i60319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60311_4_lut (.I0(n29_adj_4506), .I1(n27_adj_4505), .I2(n25_adj_4706), 
            .I3(n76175), .O(n76167));
    defparam i60311_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61947_4_lut (.I0(n35_adj_4510), .I1(n33_adj_4509), .I2(n31_adj_4508), 
            .I3(n76167), .O(n77803));
    defparam i61947_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_4708));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61751_3_lut (.I0(n16_adj_4708), .I1(baudrate[13]), .I2(n39_adj_4504), 
            .I3(GND_net), .O(n77607));   // verilog/uart_rx.v(119[33:55])
    defparam i61751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61752_3_lut (.I0(n77607), .I1(baudrate[14]), .I2(n41_adj_4503), 
            .I3(GND_net), .O(n77608));   // verilog/uart_rx.v(119[33:55])
    defparam i61752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61187_4_lut (.I0(n41_adj_4503), .I1(n39_adj_4504), .I2(n27_adj_4505), 
            .I3(n76171), .O(n77043));
    defparam i61187_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61804_3_lut (.I0(n22_adj_4709), .I1(baudrate[7]), .I2(n27_adj_4505), 
            .I3(GND_net), .O(n77660));   // verilog/uart_rx.v(119[33:55])
    defparam i61804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60751_3_lut (.I0(n77608), .I1(baudrate[15]), .I2(n43_adj_4502), 
            .I3(GND_net), .O(n76607));   // verilog/uart_rx.v(119[33:55])
    defparam i60751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1016 (.I0(baudrate[22]), .I1(baudrate[23]), 
            .I2(baudrate[31]), .I3(baudrate[30]), .O(n71436));
    defparam i1_2_lut_4_lut_adj_1016.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_4710), .I1(baudrate[9]), 
            .I2(n31_adj_4508), .I3(GND_net), .O(n28_adj_4711));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62235_4_lut (.I0(n28_adj_4711), .I1(n18_adj_4712), .I2(n31_adj_4508), 
            .I3(n76160), .O(n78091));   // verilog/uart_rx.v(119[33:55])
    defparam i62235_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62236_3_lut (.I0(n78091), .I1(baudrate[10]), .I2(n33_adj_4509), 
            .I3(GND_net), .O(n78092));   // verilog/uart_rx.v(119[33:55])
    defparam i62236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62025_3_lut (.I0(n78092), .I1(baudrate[11]), .I2(n35_adj_4510), 
            .I3(GND_net), .O(n77881));   // verilog/uart_rx.v(119[33:55])
    defparam i62025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61189_4_lut (.I0(n41_adj_4503), .I1(n39_adj_4504), .I2(n37_adj_4501), 
            .I3(n77803), .O(n77045));
    defparam i61189_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i62020_4_lut (.I0(n76607), .I1(n77660), .I2(n43_adj_4502), 
            .I3(n77043), .O(n77876));   // verilog/uart_rx.v(119[33:55])
    defparam i62020_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60749_3_lut (.I0(n77881), .I1(baudrate[12]), .I2(n37_adj_4501), 
            .I3(GND_net), .O(n76605));   // verilog/uart_rx.v(119[33:55])
    defparam i60749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62314_4_lut (.I0(n76605), .I1(n77876), .I2(n43_adj_4502), 
            .I3(n77045), .O(n78170));   // verilog/uart_rx.v(119[33:55])
    defparam i62314_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62315_3_lut (.I0(n78170), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n78171));   // verilog/uart_rx.v(119[33:55])
    defparam i62315_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8553[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8579[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8605[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_4712));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(n71436), .I1(n14_adj_4577), .I2(n9_adj_4576), 
            .I3(n71472), .O(n25970));
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'hfffe;
    SB_LUT4 i60180_4_lut (.I0(n35_adj_4479), .I1(n23_adj_4715), .I2(n21_adj_4714), 
            .I3(n19_adj_4713), .O(n76036));
    defparam i60180_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61143_4_lut (.I0(n17_adj_4476), .I1(n15_adj_4475), .I2(n2844), 
            .I3(baudrate[2]), .O(n76999));
    defparam i61143_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i61585_4_lut (.I0(n23_adj_4715), .I1(n21_adj_4714), .I2(n19_adj_4713), 
            .I3(n76999), .O(n77441));
    defparam i61585_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60304_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n76160));
    defparam i60304_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i61581_4_lut (.I0(n29_adj_4474), .I1(n27_adj_4473), .I2(n25_adj_4472), 
            .I3(n77441), .O(n77437));
    defparam i61581_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60184_4_lut (.I0(n35_adj_4479), .I1(n33_adj_4478), .I2(n31_adj_4477), 
            .I3(n77437), .O(n76040));
    defparam i60184_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_4716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_4710));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61741_3_lut (.I0(n12_adj_4716), .I1(baudrate[13]), .I2(n35_adj_4479), 
            .I3(GND_net), .O(n77597));   // verilog/uart_rx.v(119[33:55])
    defparam i61741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_4704), .I1(baudrate[17]), 
            .I2(n43_adj_4470), .I3(GND_net), .O(n38_adj_4717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61742_3_lut (.I0(n77597), .I1(baudrate[14]), .I2(n37_adj_4469), 
            .I3(GND_net), .O(n77598));   // verilog/uart_rx.v(119[33:55])
    defparam i61742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60172_4_lut (.I0(n41_adj_4471), .I1(n39_adj_4468), .I2(n37_adj_4469), 
            .I3(n76036), .O(n76028));
    defparam i60172_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62223_4_lut (.I0(n38_adj_4717), .I1(n18_adj_4694), .I2(n43_adj_4470), 
            .I3(n76022), .O(n78079));   // verilog/uart_rx.v(119[33:55])
    defparam i62223_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60767_3_lut (.I0(n77598), .I1(baudrate[15]), .I2(n39_adj_4468), 
            .I3(GND_net), .O(n76623));   // verilog/uart_rx.v(119[33:55])
    defparam i60767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_4693), .I1(baudrate[9]), 
            .I2(n27_adj_4473), .I3(GND_net), .O(n24_adj_4718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62241_4_lut (.I0(n24_adj_4718), .I1(n14_adj_4685), .I2(n27_adj_4473), 
            .I3(n76054), .O(n78097));   // verilog/uart_rx.v(119[33:55])
    defparam i62241_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62242_3_lut (.I0(n78097), .I1(baudrate[10]), .I2(n29_adj_4474), 
            .I3(GND_net), .O(n78098));   // verilog/uart_rx.v(119[33:55])
    defparam i62242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_4709));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62007_3_lut (.I0(n78098), .I1(baudrate[11]), .I2(n31_adj_4477), 
            .I3(GND_net), .O(n77863));   // verilog/uart_rx.v(119[33:55])
    defparam i62007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61929_4_lut (.I0(n41_adj_4471), .I1(n39_adj_4468), .I2(n37_adj_4469), 
            .I3(n76040), .O(n77785));
    defparam i61929_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62367_4_lut (.I0(n76623), .I1(n78079), .I2(n43_adj_4470), 
            .I3(n76028), .O(n78223));   // verilog/uart_rx.v(119[33:55])
    defparam i62367_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60765_3_lut (.I0(n77863), .I1(baudrate[12]), .I2(n33_adj_4478), 
            .I3(GND_net), .O(n76621));   // verilog/uart_rx.v(119[33:55])
    defparam i60765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62401_4_lut (.I0(n76621), .I1(n78223), .I2(n43_adj_4470), 
            .I3(n77785), .O(n78257));   // verilog/uart_rx.v(119[33:55])
    defparam i62401_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62402_3_lut (.I0(n78257), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n78258));   // verilog/uart_rx.v(119[33:55])
    defparam i62402_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60315_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n76171));
    defparam i60315_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8605[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8631[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8631[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1018 (.I0(n14_adj_4577), .I1(baudrate[28]), 
            .I2(baudrate[27]), .I3(GND_net), .O(n70620));
    defparam i1_2_lut_3_lut_adj_1018.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(baudrate[30]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n71488));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(baudrate[31]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n71486));
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1021 (.I0(n71490), .I1(n14_adj_4577), .I2(n9_adj_4576), 
            .I3(n71488), .O(n25973));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i60126_4_lut (.I0(n33_adj_4722), .I1(n21_adj_4721), .I2(n19_adj_4720), 
            .I3(n17_adj_4719), .O(n75982));
    defparam i60126_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61089_4_lut (.I0(n15_adj_4467), .I1(n13_adj_4466), .I2(n2956), 
            .I3(baudrate[2]), .O(n76945));
    defparam i61089_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i61557_4_lut (.I0(n21_adj_4721), .I1(n19_adj_4720), .I2(n17_adj_4719), 
            .I3(n76945), .O(n77413));
    defparam i61557_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61553_4_lut (.I0(n27_adj_4465), .I1(n25_adj_4464), .I2(n23_adj_4463), 
            .I3(n77413), .O(n77409));
    defparam i61553_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60128_4_lut (.I0(n33_adj_4722), .I1(n31_adj_4462), .I2(n29_adj_4461), 
            .I3(n77409), .O(n75984));
    defparam i60128_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_adj_1022 (.I0(baudrate[18]), .I1(baudrate[19]), 
            .I2(baudrate[20]), .I3(baudrate[21]), .O(n71438));
    defparam i1_2_lut_4_lut_adj_1022.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_4723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61735_3_lut (.I0(n10_adj_4723), .I1(baudrate[13]), .I2(n33_adj_4722), 
            .I3(GND_net), .O(n77591));   // verilog/uart_rx.v(119[33:55])
    defparam i61735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61736_3_lut (.I0(n77591), .I1(baudrate[14]), .I2(n35_adj_4459), 
            .I3(GND_net), .O(n77592));   // verilog/uart_rx.v(119[33:55])
    defparam i61736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_4654), .I1(baudrate[17]), 
            .I2(n41), .I3(GND_net), .O(n36_adj_4724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60118_4_lut (.I0(n39_adj_4460), .I1(n37_adj_4458), .I2(n35_adj_4459), 
            .I3(n75982), .O(n75974));
    defparam i60118_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i62010_4_lut (.I0(n36_adj_4724), .I1(n16_adj_4653), .I2(n41), 
            .I3(n75968), .O(n77866));   // verilog/uart_rx.v(119[33:55])
    defparam i62010_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60773_3_lut (.I0(n77592), .I1(baudrate[15]), .I2(n37_adj_4458), 
            .I3(GND_net), .O(n76629));   // verilog/uart_rx.v(119[33:55])
    defparam i60773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_4649), .I1(baudrate[9]), 
            .I2(n25_adj_4464), .I3(GND_net), .O(n22_adj_4725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62004_4_lut (.I0(n22_adj_4725), .I1(n12_adj_4648), .I2(n25_adj_4464), 
            .I3(n75994), .O(n77860));   // verilog/uart_rx.v(119[33:55])
    defparam i62004_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62005_3_lut (.I0(n77860), .I1(baudrate[10]), .I2(n27_adj_4465), 
            .I3(GND_net), .O(n77861));   // verilog/uart_rx.v(119[33:55])
    defparam i62005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62001_3_lut (.I0(n77861), .I1(baudrate[11]), .I2(n29_adj_4461), 
            .I3(GND_net), .O(n77857));   // verilog/uart_rx.v(119[33:55])
    defparam i62001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61919_4_lut (.I0(n39_adj_4460), .I1(n37_adj_4458), .I2(n35_adj_4459), 
            .I3(n75984), .O(n77775));
    defparam i61919_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62375_4_lut (.I0(n76629), .I1(n77866), .I2(n41), .I3(n75974), 
            .O(n78231));   // verilog/uart_rx.v(119[33:55])
    defparam i62375_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_4703));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60771_3_lut (.I0(n77857), .I1(baudrate[12]), .I2(n31_adj_4462), 
            .I3(GND_net), .O(n76627));   // verilog/uart_rx.v(119[33:55])
    defparam i60771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60359_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n76215));
    defparam i60359_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i62413_4_lut (.I0(n76627), .I1(n78231), .I2(n41), .I3(n77775), 
            .O(n78269));   // verilog/uart_rx.v(119[33:55])
    defparam i62413_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62414_3_lut (.I0(n78269), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n78270));   // verilog/uart_rx.v(119[33:55])
    defparam i62414_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62412_3_lut (.I0(n78270), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n78268));   // verilog/uart_rx.v(119[33:55])
    defparam i62412_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_4701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52069_1_lut (.I0(n25976), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67878));
    defparam i52069_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8631[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8657[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8683[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_4699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60378_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n76234));
    defparam i60378_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_4692));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60427_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n76283));
    defparam i60427_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_4690));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60433_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n76289));
    defparam i60433_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_4688));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_4684));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59482_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n75338));
    defparam i59482_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_4682));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59490_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n75346));
    defparam i59490_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_4680));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i56349_2_lut_4_lut (.I0(baudrate[20]), .I1(baudrate[21]), .I2(baudrate[30]), 
            .I3(baudrate[22]), .O(n72196));
    defparam i56349_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i60410_2_lut (.I0(n66553), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n75188));
    defparam i60410_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i62790_2_lut_4_lut (.I0(n78226), .I1(baudrate[13]), .I2(n2098), 
            .I3(n26010), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i62790_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i60400_4_lut (.I0(n75188), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n75185));
    defparam i60400_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i59728_4_lut (.I0(n75185), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n75182));
    defparam i59728_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i62850_4_lut (.I0(\r_SM_Main[2] ), .I1(n75182), .I2(r_SM_Main_2__N_3446[1]), 
            .I3(\r_SM_Main[1] ), .O(n29423));
    defparam i62850_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1023 (.I0(n66553), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n70156));
    defparam i1_4_lut_adj_1023.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1024 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n70156), .O(n70162));
    defparam i1_4_lut_adj_1024.LUT_INIT = 16'h0100;
    SB_LUT4 i62458_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n70162), .O(n28161));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i62458_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(n9_adj_4576), .I1(n14_adj_4577), .I2(n71486), 
            .I3(baudrate[30]), .O(n25979));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8683[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_4676));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8683[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59503_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n75359));
    defparam i59503_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_4673));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i63202_2_lut_4_lut (.I0(n78228), .I1(baudrate[12]), .I2(n1966), 
            .I3(n72230), .O(n294[11]));
    defparam i63202_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_4670));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i59523_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n75379));
    defparam i59523_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_4667));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8683[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52073_1_lut_4_lut (.I0(n71490), .I1(n14_adj_4577), .I2(n9_adj_4576), 
            .I3(n71488), .O(n67882));
    defparam i52073_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_4662));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59560_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n75416));
    defparam i59560_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_4659));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62696_2_lut_4_lut (.I0(n77905), .I1(baudrate[10]), .I2(n1693), 
            .I3(n26029), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i62696_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_965_i34_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n70070), .I3(n48_adj_4507), .O(n34_adj_4650));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i62616_2_lut_4_lut (.I0(n77663), .I1(baudrate[5]), .I2(n67645), 
            .I3(n26035), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i62616_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i1_2_lut_4_lut_adj_1026 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n71362));
    defparam i1_2_lut_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1027 (.I0(baudrate[28]), .I1(baudrate[27]), 
            .I2(n14_adj_4577), .I3(n71436), .O(n25976));
    defparam i1_3_lut_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8683[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62969_2_lut_4_lut (.I0(n77667), .I1(baudrate[4]), .I2(n67643), 
            .I3(n72256), .O(n294[19]));
    defparam i62969_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i60351_2_lut_3_lut (.I0(n25991), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n75234));   // verilog/uart_rx.v(119[33:55])
    defparam i60351_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i62999_4_lut_4_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(n6_adj_4726), .I3(n69436), .O(n67800));
    defparam i62999_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i59692_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4637), .I2(n25991), 
            .I3(GND_net), .O(n75548));   // verilog/uart_rx.v(119[33:55])
    defparam i59692_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_4727));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5217), 
            .O(n15_adj_4728));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4728), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_4727), 
            .I3(n66790), .O(n79649));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_3_lut_4_lut_adj_1028 (.I0(baudrate[14]), .I1(baudrate[2]), 
            .I2(baudrate[1]), .I3(baudrate[0]), .O(n70512));
    defparam i1_3_lut_4_lut_adj_1028.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_adj_1029 (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n72260), .I3(GND_net), .O(n45376));
    defparam i1_2_lut_3_lut_adj_1029.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_1030 (.I0(n25991), .I1(n48_adj_4637), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_4638));
    defparam i1_3_lut_4_lut_adj_1030.LUT_INIT = 16'hefff;
    SB_LUT4 i59695_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4640), .I2(n26022), 
            .I3(GND_net), .O(n75551));   // verilog/uart_rx.v(119[33:55])
    defparam i59695_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i5659_2_lut_3_lut (.I0(n21179), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_4578));   // verilog/uart_rx.v(119[33:55])
    defparam i5659_2_lut_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 i7309_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n21179));   // verilog/uart_rx.v(119[33:55])
    defparam i7309_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70328), .O(n70334));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70334), .O(n70340));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1033 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n5220), 
            .I3(GND_net), .O(n70104));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n70104), .O(\r_SM_Main_2__N_3536[1] ));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i5828_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n11692));   // verilog/uart_rx.v(119[33:55])
    defparam i5828_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70344), .O(n70350));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70350), .O(n70356));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70264), .O(n70270));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70270), .O(n70276));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1039 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[10]), .I3(baudrate[11]), .O(n71360));
    defparam i1_2_lut_3_lut_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1040 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70312), .O(n70318));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1041 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70318), .O(n70324));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n28));
    defparam i10_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1042 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70296), .O(n70302));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1042.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70302), .O(n70308));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70376), .O(n70382));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n70624));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_271_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4729));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70382), .O(n70388));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1047 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70376));
    defparam i1_3_lut_4_lut_adj_1047.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_4_lut_adj_1048 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n70360), .O(n70366));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1048.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1049 (.I0(r_Clock_Count[3]), .I1(n3_adj_4729), 
            .I2(\o_Rx_DV_N_3488[4] ), .I3(n70624), .O(n70628));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1049.LUT_INIT = 16'hffde;
    SB_LUT4 equal_271_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4730));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1050 (.I0(r_Clock_Count[5]), .I1(n5_adj_4730), 
            .I2(\o_Rx_DV_N_3488[6] ), .I3(n70628), .O(n70632));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1050.LUT_INIT = 16'hffde;
    SB_LUT4 equal_271_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4731));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1051 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70360));
    defparam i1_3_lut_4_lut_adj_1051.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_4_lut_adj_1052 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70366), .O(n70372));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1052.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1053 (.I0(r_Clock_Count[6]), .I1(n8_adj_4731), 
            .I2(n70632), .I3(\o_Rx_DV_N_3488[7] ), .O(n66553));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1053.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_3_lut_4_lut_adj_1054 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70296));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1054.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1055 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70312));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1055.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut_4_lut_adj_1056 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70344));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1056.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_3_lut_4_lut_adj_1057 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70264));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1057.LUT_INIT = 16'hffdf;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5217), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n69436), .O(n70196));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1059 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n70196), .O(n70202));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1059.LUT_INIT = 16'hfffe;
    SB_LUT4 i56307_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n66553), .I2(GND_net), 
            .I3(GND_net), .O(n72154));
    defparam i56307_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8683[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56373_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n72154), .O(n72220));
    defparam i56373_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n70202), .I1(r_SM_Main_2__N_3446[1]), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n72220), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n11917));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n11917), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_3_lut_4_lut_adj_1060 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70328));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1060.LUT_INIT = 16'hffef;
    SB_LUT4 i1_3_lut_4_lut_adj_1061 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4584), .O(n70280));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1061.LUT_INIT = 16'hfffe;
    SB_LUT4 i52085_1_lut_2_lut (.I0(n70620), .I1(n71442), .I2(GND_net), 
            .I3(GND_net), .O(n67894));
    defparam i52085_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i5837_2_lut_3_lut_4_lut (.I0(baudrate[3]), .I1(n21189), .I2(n11692), 
            .I3(n960), .O(n44_adj_4629));   // verilog/uart_rx.v(119[33:55])
    defparam i5837_2_lut_3_lut_4_lut.LUT_INIT = 16'hfd54;
    SB_LUT4 i52093_1_lut_4_lut (.I0(n14_adj_4577), .I1(n9_adj_4576), .I2(n71462), 
            .I3(n71438), .O(n67902));
    defparam i52093_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i56386_1_lut_2_lut (.I0(baudrate[12]), .I1(n72230), .I2(GND_net), 
            .I3(GND_net), .O(n67915));
    defparam i56386_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i5666_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(n21179), .I2(n44852), 
            .I3(n804), .O(n44_adj_4635));   // verilog/uart_rx.v(119[33:55])
    defparam i5666_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf45;
    SB_LUT4 i1_4_lut_adj_1062 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n5220), 
            .I3(\r_SM_Main[0] ), .O(n70138));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1062.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1063 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n70138), .O(n68353));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1063.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1064 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[31]), .I3(baudrate[30]), .O(n71478));
    defparam i1_2_lut_4_lut_adj_1064.LUT_INIT = 16'hfffe;
    SB_LUT4 i63245_2_lut_4_lut (.I0(n78037), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25979), .O(n294[1]));
    defparam i63245_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_4569));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_4568));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59997_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n75853));
    defparam i59997_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_4567));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_4570));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60020_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n75876));
    defparam i60020_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1065 (.I0(baudrate[28]), .I1(baudrate[27]), 
            .I2(n14_adj_4577), .I3(n71470), .O(n70018));
    defparam i1_3_lut_4_lut_adj_1065.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8683[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_4500));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60252_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n76108));
    defparam i60252_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_4499));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60222_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n76078));
    defparam i60222_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1066 (.I0(n78268), .I1(baudrate[20]), .I2(n2938), 
            .I3(n70088), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1066.LUT_INIT = 16'h7100;
    SB_LUT4 i63226_2_lut_4_lut (.I0(n78268), .I1(baudrate[20]), .I2(n2938), 
            .I3(n25973), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i63226_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1067 (.I0(n78258), .I1(baudrate[19]), .I2(n2827), 
            .I3(n70086), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1067.LUT_INIT = 16'h7100;
    SB_LUT4 i63223_2_lut_4_lut (.I0(n78258), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25970), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i63223_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1068 (.I0(n78171), .I1(baudrate[17]), .I2(n2596), 
            .I3(n70082), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1068.LUT_INIT = 16'h7100;
    SB_LUT4 i63217_2_lut_4_lut (.I0(n78171), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25937), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i63217_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1069 (.I0(n77659), .I1(baudrate[16]), .I2(n2476), 
            .I3(n70080), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1069.LUT_INIT = 16'h7100;
    SB_LUT4 i63214_2_lut_4_lut (.I0(n77659), .I1(baudrate[16]), .I2(n2476), 
            .I3(n26019), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i63214_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i2314_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2314_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_2_lut_4_lut_adj_1070 (.I0(n78113), .I1(baudrate[15]), .I2(n2353), 
            .I3(n70078), .O(n2491));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1070.LUT_INIT = 16'h7100;
    SB_LUT4 i63211_2_lut_4_lut (.I0(n78113), .I1(baudrate[15]), .I2(n2353), 
            .I3(n26016), .O(n294[8]));   // verilog/uart_rx.v(119[33:55])
    defparam i63211_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60046_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n75902));
    defparam i60046_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n5217), 
            .I3(\o_Rx_DV_N_3488[8] ), .O(n70062));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n70062), .O(r_SM_Main_2__N_3446[1]));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1073 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n71474), .I3(n70654), .O(n71418));
    defparam i1_3_lut_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4726));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n69436));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i60072_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n75928));
    defparam i60072_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1074 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[15]), .I3(baudrate[14]), .O(n71358));
    defparam i1_2_lut_3_lut_4_lut_adj_1074.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1075 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n71436), .I3(GND_net), .O(n71462));
    defparam i1_2_lut_3_lut_adj_1075.LUT_INIT = 16'hfefe;
    SB_LUT4 i2307_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2307_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i63208_2_lut_4_lut (.I0(n78166), .I1(baudrate[14]), .I2(n2227), 
            .I3(n72228), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i63208_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1076 (.I0(n78166), .I1(baudrate[14]), .I2(n2227), 
            .I3(n70076), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1076.LUT_INIT = 16'h7100;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (GND_net, VCC_net, n5, n5_adj_3, n5_adj_4, state_7__N_4319, 
            n44711, clk16MHz, CS_c, CS_CLK_c, n30119, \data[15] , 
            n30118, \data[12] , n30117, \data[11] , n30116, \data[10] , 
            n30115, \data[9] , n30114, \data[8] , n30113, \data[7] , 
            n30112, \data[6] , n30111, \data[5] , n30110, \data[4] , 
            n30109, \data[3] , n30108, \data[2] , n30107, \data[1] , 
            n29947, \current[0] , n30767, \data[0] , n30677, \current[1] , 
            n30676, \current[2] , n30675, \current[3] , n30674, \current[4] , 
            n30673, \current[5] , n30672, \current[6] , n30671, \current[7] , 
            n30670, \current[8] , n30669, \current[9] , n30668, \current[10] , 
            n30667, \current[11] , n28099, \current[15] , n25895, 
            n11, n25912, n25869, n25885) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    output n5;
    output n5_adj_3;
    output n5_adj_4;
    output state_7__N_4319;
    output n44711;
    input clk16MHz;
    output CS_c;
    output CS_CLK_c;
    input n30119;
    output \data[15] ;
    input n30118;
    output \data[12] ;
    input n30117;
    output \data[11] ;
    input n30116;
    output \data[10] ;
    input n30115;
    output \data[9] ;
    input n30114;
    output \data[8] ;
    input n30113;
    output \data[7] ;
    input n30112;
    output \data[6] ;
    input n30111;
    output \data[5] ;
    input n30110;
    output \data[4] ;
    input n30109;
    output \data[3] ;
    input n30108;
    output \data[2] ;
    input n30107;
    output \data[1] ;
    input n29947;
    output \current[0] ;
    input n30767;
    output \data[0] ;
    input n30677;
    output \current[1] ;
    input n30676;
    output \current[2] ;
    input n30675;
    output \current[3] ;
    input n30674;
    output \current[4] ;
    input n30673;
    output \current[5] ;
    input n30672;
    output \current[6] ;
    input n30671;
    output \current[7] ;
    input n30670;
    output \current[8] ;
    input n30669;
    output \current[9] ;
    input n30668;
    output \current[10] ;
    input n30667;
    output \current[11] ;
    output n28099;
    output \current[15] ;
    output n25895;
    output n11;
    output n25912;
    output n25869;
    output n25885;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n60282, n60281;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n60280, n60279, n60278, n60277, n60276, n60275;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n60274, n60273;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n60272, n60271, n60270, clk_slow_N_4232;
    wire [7:0]n37;
    
    wire n60256, n60255, n60254, n60253, n75191, n60252, n2, n75180, 
        n60251, n75172, n60250, n75192, clk_out, n29949, n15, 
        n9, n12495, n28263, n29167, n22862, n28156, delay_counter_15__N_4314, 
        clk_slow_N_4233, n22864, n22866, n22868, n29435;
    wire [13:0]n241;
    
    wire n45285, n4, n8, n12, n10;
    
    SB_LUT4 counter_2050_2051_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n60282), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2050_2051_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n60281), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_3 (.CI(n60281), .I0(GND_net), .I1(counter[1]), 
            .CO(n60282));
    SB_LUT4 counter_2050_2051_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n60281));
    SB_LUT4 delay_counter_2048_2049_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n60280), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2048_2049_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n60279), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_12 (.CI(n60279), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n60280));
    SB_LUT4 delay_counter_2048_2049_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n60278), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_11 (.CI(n60278), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n60279));
    SB_LUT4 delay_counter_2048_2049_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n60277), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_10 (.CI(n60277), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n60278));
    SB_LUT4 delay_counter_2048_2049_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n60276), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_9 (.CI(n60276), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n60277));
    SB_LUT4 delay_counter_2048_2049_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n60275), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 equal_337_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_337_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_328_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_CARRY delay_counter_2048_2049_add_4_8 (.CI(n60275), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n60276));
    SB_LUT4 delay_counter_2048_2049_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n60274), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_7 (.CI(n60274), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n60275));
    SB_LUT4 equal_330_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4));   // verilog/tli4970.v(54[9:26])
    defparam equal_330_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 delay_counter_2048_2049_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n60273), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4319));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_CARRY delay_counter_2048_2049_add_4_6 (.CI(n60273), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n60274));
    SB_LUT4 delay_counter_2048_2049_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n60272), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_5 (.CI(n60272), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n60273));
    SB_LUT4 delay_counter_2048_2049_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n60271), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_4 (.CI(n60271), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n60272));
    SB_LUT4 delay_counter_2048_2049_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n60270), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_3 (.CI(n60270), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n60271));
    SB_LUT4 i30622_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n44711));
    defparam i30622_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 delay_counter_2048_2049_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n60270));
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4232));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 bit_counter_2044_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n60256), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2044_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n60255), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_8 (.CI(n60255), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n60256));
    SB_LUT4 bit_counter_2044_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n60254), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_7 (.CI(n60254), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n60255));
    SB_LUT4 bit_counter_2044_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n60253), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_6 (.CI(n60253), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n60254));
    SB_LUT4 bit_counter_2044_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n60252), .O(n75191)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_5 (.CI(n60252), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n60253));
    SB_LUT4 bit_counter_2044_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n60251), .O(n75180)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_4 (.CI(n60251), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n60252));
    SB_LUT4 bit_counter_2044_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n60250), .O(n75172)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_3 (.CI(n60250), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n60251));
    SB_LUT4 bit_counter_2044_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n75192)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n60250));
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n30119));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n30118));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n30117));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n30116));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n30115));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n30114));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n30113));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n30112));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n30111));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n30110));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n30109));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n30108));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n30107));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i15735_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n29949));
    defparam i15735_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i63229_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9));
    defparam i63229_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n28263), .D(n12495), 
            .R(n29167));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29949));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29947));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n28156), 
            .D(n22862));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2050_2051__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2050_2051__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_2048_2049__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNE bit_counter_2044__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n28156), 
            .D(n22864));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2044__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n28156), 
            .D(n22866));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2044__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n28156), 
            .D(n22868));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n28156), 
            .D(n37[4]), .R(n29435));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n28156), 
            .D(n37[5]), .R(n29435));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n28156), 
            .D(n37[6]), .R(n29435));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n28156), 
            .D(n37[7]), .R(n29435));   // verilog/tli4970.v(55[24:39])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30767));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n30677));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n30676));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n30675));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n30674));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n30673));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n30672));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n30671));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n30670));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n30669));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n30668));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n30667));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(delay_counter_15__N_4314), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n28263));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 i14953_2_lut_4_lut (.I0(delay_counter_15__N_4314), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n29167));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14953_2_lut_4_lut.LUT_INIT = 16'h2202;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n28099), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(state[0]), .I3(state[1]), .O(n25895));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_268_i11_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n11));   // verilog/tli4970.v(54[9:26])
    defparam equal_268_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n28263), .D(n45285), 
            .S(n29167));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_966 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n25912));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_966.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_967 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n25869));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_967.LUT_INIT = 16'hffbf;
    SB_LUT4 i62479_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n45285));
    defparam i62479_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i15222_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29435));   // verilog/tli4970.v(55[24:39])
    defparam i15222_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2243_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2243_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2521_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));
    defparam i2521_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8936_3_lut (.I0(state[0]), .I1(n75172), .I2(state[1]), .I3(GND_net), 
            .O(n22868));   // verilog/tli4970.v(55[24:39])
    defparam i8936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8934_3_lut (.I0(state[0]), .I1(n75180), .I2(state[1]), .I3(GND_net), 
            .O(n22866));   // verilog/tli4970.v(55[24:39])
    defparam i8934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8932_3_lut (.I0(state[0]), .I1(n75191), .I2(state[1]), .I3(GND_net), 
            .O(n22864));   // verilog/tli4970.v(55[24:39])
    defparam i8932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14096_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n28156));
    defparam i14096_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8930_3_lut (.I0(state[0]), .I1(n75192), .I2(state[1]), .I3(GND_net), 
            .O(n22862));   // verilog/tli4970.v(55[24:39])
    defparam i8930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2179_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4233));
    defparam i2179_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4233), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4232));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62471_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n28099));
    defparam i62471_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut (.I0(bit_counter[4]), .I1(bit_counter[6]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(n11), .I1(bit_counter[5]), .I2(bit_counter[7]), 
            .I3(n4), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i2_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2180_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2180_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(delay_counter[11]), .I1(delay_counter[7]), .I2(delay_counter[8]), 
            .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4314));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 mux_2153_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n12495));
    defparam mux_2153_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(state[0]), 
            .I3(state[1]), .O(n25885));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2874, pwm_out, clk32MHz, \pwm_counter[7] , GND_net, \pwm_counter[16] , 
            \pwm_counter[20] , \pwm_counter[19] , \pwm_counter[12] , \pwm_setpoint[18] , 
            \pwm_setpoint[17] , \pwm_counter[4] , VCC_net, reset, \pwm_setpoint[22] , 
            \pwm_setpoint[21] , \pwm_setpoint[11] , \pwm_setpoint[10] , 
            \pwm_setpoint[9] , \pwm_setpoint[6] , \pwm_setpoint[8] , \pwm_setpoint[3] , 
            \pwm_setpoint[5] , \pwm_setpoint[2] , n9, n15, \pwm_setpoint[1] , 
            \pwm_setpoint[0] , \pwm_setpoint[7] , \pwm_setpoint[12] , 
            n25, \pwm_setpoint[13] , \pwm_setpoint[14] , \pwm_setpoint[15] , 
            n32, n34, \pwm_setpoint[20] , n41, n39, \pwm_setpoint[19] , 
            \pwm_setpoint[23] , \pwm_setpoint[4] ) /* synthesis syn_module_defined=1 */ ;
    input n2874;
    output pwm_out;
    input clk32MHz;
    output \pwm_counter[7] ;
    input GND_net;
    output \pwm_counter[16] ;
    output \pwm_counter[20] ;
    output \pwm_counter[19] ;
    output \pwm_counter[12] ;
    input \pwm_setpoint[18] ;
    input \pwm_setpoint[17] ;
    output \pwm_counter[4] ;
    input VCC_net;
    input reset;
    input \pwm_setpoint[22] ;
    input \pwm_setpoint[21] ;
    input \pwm_setpoint[11] ;
    input \pwm_setpoint[10] ;
    input \pwm_setpoint[9] ;
    input \pwm_setpoint[6] ;
    input \pwm_setpoint[8] ;
    input \pwm_setpoint[3] ;
    input \pwm_setpoint[5] ;
    input \pwm_setpoint[2] ;
    input n9;
    input n15;
    input \pwm_setpoint[1] ;
    input \pwm_setpoint[0] ;
    input \pwm_setpoint[7] ;
    input \pwm_setpoint[12] ;
    input n25;
    input \pwm_setpoint[13] ;
    input \pwm_setpoint[14] ;
    input \pwm_setpoint[15] ;
    output n32;
    input n34;
    input \pwm_setpoint[20] ;
    input n41;
    input n39;
    input \pwm_setpoint[19] ;
    input \pwm_setpoint[23] ;
    input \pwm_setpoint[4] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_577;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n69874, n22, n15_c, n20, n24, n19, n45, n76231, n65178, 
        n60187, n65218, n60186, n65250, n60185, n65290, n60184, 
        n65330, n60183, n36, n65370, n60182, n65408, n60181, n65446, 
        n60180, n65480, n60179, n65524, n60178, n65560, n60177, 
        n65598, n60176, n65632, n60175, n65664, n60174, n65704, 
        n60173, n65756, n60172, n65798, n60171, n65860, n60170, 
        n65968, n60169, n66136, n60168, n66278, n60167, n66280, 
        n60166, n66282, n60165, n66268, n45_adj_4450, n43, n23, 
        n21, n19_adj_4451, n13, n17, n7, n11, n5, n76275, n76264, 
        n4, n10, n12, n8, n16, n6, n76262, n78055, n78056, 
        n77959, n77809, n76270, n77954, n76431, n78057, n78058, 
        n77953, n77739, n77740, n77095, n38, n76439, n77547;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2874), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(\pwm_counter[7] ), 
            .I3(GND_net), .O(n69874));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[11]), .I1(pwm_counter[18]), .I2(pwm_counter[15]), 
            .I3(pwm_counter[13]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n69874), .I1(\pwm_counter[16] ), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_c));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(\pwm_counter[20] ), .I1(pwm_counter[22]), .I2(pwm_counter[14]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_c), .I1(n22), .I2(\pwm_counter[19] ), .I3(\pwm_counter[12] ), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[17]), .I1(pwm_counter[21]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(n45));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60375_3_lut_4_lut (.I0(pwm_counter[18]), .I1(\pwm_setpoint[18] ), 
            .I2(\pwm_setpoint[17] ), .I3(pwm_counter[17]), .O(n76231));   // verilog/pwm.v(21[8:24])
    defparam i60375_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 pwm_counter_2040_add_4_25_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n60187), .O(n65178)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_2040_add_4_24_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n60186), .O(n65218)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_24 (.CI(n60186), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n60187));
    SB_LUT4 pwm_counter_2040_add_4_23_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n60185), .O(n65250)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_23 (.CI(n60185), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n60186));
    SB_LUT4 pwm_counter_2040_add_4_22_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[20] ), 
            .I3(n60184), .O(n65290)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_22 (.CI(n60184), .I0(GND_net), .I1(\pwm_counter[20] ), 
            .CO(n60185));
    SB_LUT4 pwm_counter_2040_add_4_21_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[19] ), 
            .I3(n60183), .O(n65330)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_21 (.CI(n60183), .I0(GND_net), .I1(\pwm_counter[19] ), 
            .CO(n60184));
    SB_LUT4 duty_23__I_0_i36_3_lut_3_lut (.I0(pwm_counter[18]), .I1(\pwm_setpoint[18] ), 
            .I2(\pwm_setpoint[17] ), .I3(GND_net), .O(n36));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 pwm_counter_2040_add_4_20_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n60182), .O(n65370)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_20 (.CI(n60182), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n60183));
    SB_LUT4 pwm_counter_2040_add_4_19_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n60181), .O(n65408)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_19 (.CI(n60181), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n60182));
    SB_LUT4 pwm_counter_2040_add_4_18_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[16] ), 
            .I3(n60180), .O(n65446)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_18 (.CI(n60180), .I0(GND_net), .I1(\pwm_counter[16] ), 
            .CO(n60181));
    SB_LUT4 pwm_counter_2040_add_4_17_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n60179), .O(n65480)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_17 (.CI(n60179), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n60180));
    SB_LUT4 pwm_counter_2040_add_4_16_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n60178), .O(n65524)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_16 (.CI(n60178), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n60179));
    SB_LUT4 pwm_counter_2040_add_4_15_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n60177), .O(n65560)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_15 (.CI(n60177), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n60178));
    SB_LUT4 pwm_counter_2040_add_4_14_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[12] ), 
            .I3(n60176), .O(n65598)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_14 (.CI(n60176), .I0(GND_net), .I1(\pwm_counter[12] ), 
            .CO(n60177));
    SB_LUT4 pwm_counter_2040_add_4_13_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n60175), .O(n65632)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_13 (.CI(n60175), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n60176));
    SB_LUT4 pwm_counter_2040_add_4_12_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n60174), .O(n65664)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_12 (.CI(n60174), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n60175));
    SB_LUT4 pwm_counter_2040_add_4_11_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n60173), .O(n65704)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_11 (.CI(n60173), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n60174));
    SB_LUT4 pwm_counter_2040_add_4_10_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n60172), .O(n65756)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_10 (.CI(n60172), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n60173));
    SB_LUT4 pwm_counter_2040_add_4_9_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[7] ), 
            .I3(n60171), .O(n65798)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_9 (.CI(n60171), .I0(GND_net), .I1(\pwm_counter[7] ), 
            .CO(n60172));
    SB_LUT4 pwm_counter_2040_add_4_8_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n60170), .O(n65860)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_8 (.CI(n60170), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n60171));
    SB_LUT4 pwm_counter_2040_add_4_7_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n60169), .O(n65968)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_7 (.CI(n60169), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n60170));
    SB_LUT4 pwm_counter_2040_add_4_6_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[4] ), 
            .I3(n60168), .O(n66136)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_6 (.CI(n60168), .I0(GND_net), .I1(\pwm_counter[4] ), 
            .CO(n60169));
    SB_LUT4 pwm_counter_2040_add_4_5_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n60167), .O(n66278)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_5 (.CI(n60167), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n60168));
    SB_LUT4 pwm_counter_2040_add_4_4_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n60166), .O(n66280)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_4 (.CI(n60166), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n60167));
    SB_LUT4 pwm_counter_2040_add_4_3_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n60165), .O(n66282)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_3 (.CI(n60165), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n60166));
    SB_LUT4 pwm_counter_2040_add_4_2_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n66268)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n60165));
    SB_DFFR pwm_counter_2040__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n66268), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n65178), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n65218), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n65250), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i20 (.Q(\pwm_counter[20] ), .C(clk32MHz), 
            .D(n65290), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i19 (.Q(\pwm_counter[19] ), .C(clk32MHz), 
            .D(n65330), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n65370), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n65408), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i16 (.Q(\pwm_counter[16] ), .C(clk32MHz), 
            .D(n65446), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n65480), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n65524), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n65560), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i12 (.Q(\pwm_counter[12] ), .C(clk32MHz), 
            .D(n65598), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n65632), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n65664), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n65704), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n65756), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i7 (.Q(\pwm_counter[7] ), .C(clk32MHz), .D(n65798), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n65860), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n65968), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i4 (.Q(\pwm_counter[4] ), .C(clk32MHz), .D(n66136), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n66278), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n66280), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n66282), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(\pwm_setpoint[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4450));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(\pwm_setpoint[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(\pwm_setpoint[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(\pwm_setpoint[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(\pwm_setpoint[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4451));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(\pwm_setpoint[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(\pwm_setpoint[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i7_2_lut (.I0(pwm_counter[3]), .I1(\pwm_setpoint[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(\pwm_setpoint[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i5_2_lut (.I0(pwm_counter[2]), .I1(\pwm_setpoint[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i60419_4_lut (.I0(n11), .I1(n9), .I2(n7), .I3(n5), .O(n76275));
    defparam i60419_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60408_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n76275), 
            .O(n76264));
    defparam i60408_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(\pwm_setpoint[1] ), 
            .I2(pwm_counter[1]), .I3(\pwm_setpoint[0] ), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(n10), .I1(\pwm_setpoint[7] ), .I2(n15), 
            .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(n8), .I1(\pwm_setpoint[9] ), .I2(n19_adj_4451), 
            .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62199_4_lut (.I0(n16), .I1(n6), .I2(n19_adj_4451), .I3(n76262), 
            .O(n78055));   // verilog/pwm.v(21[8:24])
    defparam i62199_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62200_3_lut (.I0(n78055), .I1(\pwm_setpoint[10] ), .I2(n21), 
            .I3(GND_net), .O(n78056));   // verilog/pwm.v(21[8:24])
    defparam i62200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62103_3_lut (.I0(n78056), .I1(\pwm_setpoint[11] ), .I2(n23), 
            .I3(GND_net), .O(n77959));   // verilog/pwm.v(21[8:24])
    defparam i62103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61953_4_lut (.I0(n23), .I1(n21), .I2(n19_adj_4451), .I3(n76264), 
            .O(n77809));
    defparam i61953_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62098_4_lut (.I0(n12), .I1(n4), .I2(n15), .I3(n76270), 
            .O(n77954));   // verilog/pwm.v(21[8:24])
    defparam i62098_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60575_3_lut (.I0(n77959), .I1(\pwm_setpoint[12] ), .I2(n25), 
            .I3(GND_net), .O(n76431));   // verilog/pwm.v(21[8:24])
    defparam i60575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62201_4_lut (.I0(n76431), .I1(n77954), .I2(n25), .I3(n77809), 
            .O(n78057));   // verilog/pwm.v(21[8:24])
    defparam i62201_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i62202_3_lut (.I0(n78057), .I1(\pwm_setpoint[13] ), .I2(pwm_counter[13]), 
            .I3(GND_net), .O(n78058));   // verilog/pwm.v(21[8:24])
    defparam i62202_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i62097_3_lut (.I0(n78058), .I1(\pwm_setpoint[14] ), .I2(pwm_counter[14]), 
            .I3(GND_net), .O(n77953));   // verilog/pwm.v(21[8:24])
    defparam i62097_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60581_3_lut (.I0(n77953), .I1(\pwm_setpoint[15] ), .I2(pwm_counter[15]), 
            .I3(GND_net), .O(n32));   // verilog/pwm.v(21[8:24])
    defparam i60581_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61883_3_lut (.I0(n34), .I1(\pwm_setpoint[20] ), .I2(n41), 
            .I3(GND_net), .O(n77739));   // verilog/pwm.v(21[8:24])
    defparam i61883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61884_3_lut (.I0(n77739), .I1(\pwm_setpoint[21] ), .I2(n43), 
            .I3(GND_net), .O(n77740));   // verilog/pwm.v(21[8:24])
    defparam i61884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61239_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n76231), 
            .O(n77095));
    defparam i61239_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 duty_23__I_0_i38_3_lut (.I0(n36), .I1(\pwm_setpoint[19] ), .I2(n39), 
            .I3(GND_net), .O(n38));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60583_3_lut (.I0(n77740), .I1(\pwm_setpoint[22] ), .I2(n45_adj_4450), 
            .I3(GND_net), .O(n76439));   // verilog/pwm.v(21[8:24])
    defparam i60583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61691_4_lut (.I0(n76439), .I1(n38), .I2(n45_adj_4450), .I3(n77095), 
            .O(n77547));   // verilog/pwm.v(21[8:24])
    defparam i61691_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61692_3_lut (.I0(n77547), .I1(pwm_counter[23]), .I2(\pwm_setpoint[23] ), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i61692_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(\pwm_setpoint[2] ), .I1(\pwm_setpoint[3] ), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60406_2_lut_4_lut (.I0(pwm_counter[8]), .I1(\pwm_setpoint[8] ), 
            .I2(\pwm_counter[4] ), .I3(\pwm_setpoint[4] ), .O(n76262));
    defparam i60406_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(\pwm_setpoint[4] ), .I1(\pwm_setpoint[8] ), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60414_2_lut_4_lut (.I0(pwm_counter[6]), .I1(\pwm_setpoint[6] ), 
            .I2(pwm_counter[5]), .I3(\pwm_setpoint[5] ), .O(n76270));
    defparam i60414_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(\pwm_setpoint[5] ), .I1(\pwm_setpoint[6] ), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, enable_slow_N_4213, clk16MHz, data, baudrate, 
            n28272, \state_7__N_3918[0] , data_ready, ID, n30714, 
            n30713, n30712, n30711, n30710, n30709, n30708, n30707, 
            n30697, n30696, n30695, n30694, n30693, n30692, n30691, 
            n30690, \state[0] , n28274, \state_7__N_4110[0] , scl_enable, 
            sda_enable, sda_out, n29970, n29969, n29967, n29966, 
            n29965, n29961, n29960, n6707, n30751, n8, VCC_net, 
            n11, \state_7__N_4126[3] , n44639, n10, n4, n4_adj_2, 
            n25890, n25932, n44782, scl) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    output enable_slow_N_4213;
    input clk16MHz;
    output [7:0]data;
    output [31:0]baudrate;
    output n28272;
    input \state_7__N_3918[0] ;
    output data_ready;
    output [7:0]ID;
    input n30714;
    input n30713;
    input n30712;
    input n30711;
    input n30710;
    input n30709;
    input n30708;
    input n30707;
    input n30697;
    input n30696;
    input n30695;
    input n30694;
    input n30693;
    input n30692;
    input n30691;
    input n30690;
    output \state[0] ;
    output n28274;
    output \state_7__N_4110[0] ;
    output scl_enable;
    output sda_enable;
    output sda_out;
    input n29970;
    input n29969;
    input n29967;
    input n29966;
    input n29965;
    input n29961;
    input n29960;
    output n6707;
    input n30751;
    input n8;
    input VCC_net;
    output n11;
    input \state_7__N_4126[3] ;
    output n44639;
    output n10;
    output n4;
    output n4_adj_2;
    output n25890;
    output n25932;
    output n44782;
    output scl;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]state;   // verilog/eeprom.v(27[11:16])
    
    wire n38017, ready_prev, n44651, n117, n125, n52995, n30682;
    wire [0:0]n5927;
    
    wire enable, n52984, n30683;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n66792, n28, n4_c, n47, n4_adj_4440, n28758, n75297, 
        n10_c, n67746, n65784, n30106;
    wire [15:0]delay_counter_15__N_3956;
    
    wire n28091;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n52961, n65940, rw, n29946, n29945;
    wire [2:0]n1;
    
    wire n28163, n29432, n61529, n30721, n30720, n30719, n30718, 
        n30717, n30716, n30715, n30706, n30705, n30704, n30703, 
        n30702, n30701, n30700, n30698, n30689, n30688, n30687, 
        n30686, n30685, n30684;
    wire [7:0]state_7__N_3885;
    
    wire n69251, n25752;
    wire [15:0]n5393;
    
    wire n59150, n59149, n59148, n15, n6938, n6937, n6936, n6935, 
        n6934, n6932, n59147, n59146, n59145, n52946, n59144, 
        n59143, n59142, n59141, n59140, n59139, n59138, n59137, 
        n59136;
    wire [7:0]state_adj_4449;   // verilog/i2c_controller.v(33[12:17])
    
    wire n72174, n75328, n17, n52949, n7, n45262, n28_adj_4444, 
        n26, n27, n25, n60942, n10_adj_4445;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n66328;
    
    SB_LUT4 i1_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n38017));   // verilog/eeprom.v(27[11:16])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i30562_2_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n44651));
    defparam i30562_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4213));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i38921_4_lut (.I0(n117), .I1(n125), .I2(data[7]), .I3(baudrate[31]), 
            .O(n52995));   // verilog/eeprom.v(23[12:16])
    defparam i38921_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i38922_3_lut (.I0(n52995), .I1(baudrate[31]), .I2(state[2]), 
            .I3(GND_net), .O(n30682));   // verilog/eeprom.v(27[11:16])
    defparam i38922_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5927[0]), .R(state[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i38910_4_lut (.I0(n117), .I1(n125), .I2(data[6]), .I3(baudrate[30]), 
            .O(n52984));   // verilog/eeprom.v(23[12:16])
    defparam i38910_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i38911_3_lut (.I0(n52984), .I1(baudrate[30]), .I2(state[2]), 
            .I3(GND_net), .O(n30683));   // verilog/eeprom.v(27[11:16])
    defparam i38911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(byte_counter[1]), .I1(n66792), .I2(n28), .I3(GND_net), 
            .O(n28272));   // verilog/eeprom.v(35[8] 81[4])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_adj_954 (.I0(state[2]), .I1(byte_counter[2]), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n66792));   // verilog/eeprom.v(35[8] 81[4])
    defparam i2_3_lut_adj_954.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\state_7__N_3918[0] ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'heeee;
    SB_LUT4 i62420_3_lut (.I0(n47), .I1(n44651), .I2(state[0]), .I3(GND_net), 
            .O(n4_adj_4440));
    defparam i62420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(state[1]), .I1(state[2]), .I2(n4_adj_4440), 
            .I3(n4_c), .O(n28758));
    defparam i2_4_lut.LUT_INIT = 16'hecfd;
    SB_LUT4 i59755_3_lut (.I0(n28758), .I1(state[2]), .I2(\state_7__N_3918[0] ), 
            .I3(GND_net), .O(n75297));   // verilog/eeprom.v(27[11:16])
    defparam i59755_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i28_4_lut (.I0(n75297), .I1(n47), .I2(state[1]), .I3(n28758), 
            .O(n10_c));   // verilog/eeprom.v(27[11:16])
    defparam i28_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i27_4_lut (.I0(n10_c), .I1(n67746), .I2(state[0]), .I3(state[2]), 
            .O(n65784));   // verilog/eeprom.v(27[11:16])
    defparam i27_4_lut.LUT_INIT = 16'hfaca;
    SB_DFF state_i2 (.Q(state[2]), .C(clk16MHz), .D(n30106));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n28091), .D(delay_counter_15__N_3956[13]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n65940));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n29946));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29945));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_2047__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n28163), .D(n1[1]), .R(n29432));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2047__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n28163), .D(n1[2]), .R(n29432));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2047__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n28163), .D(n61529), .R(n29432));   // verilog/eeprom.v(68[25:39])
    SB_DFF state_i0 (.Q(state[0]), .C(clk16MHz), .D(n65784));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n30721));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n30720));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n30719));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n30718));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n30717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n30716));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n30715));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n30714));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n30713));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n30712));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n30711));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n30710));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n30709));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n30708));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n30707));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n30706));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n30705));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n30704));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n30703));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n30702));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n30701));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n30700));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n30698));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n30697));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n30696));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n30695));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n30694));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n30693));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n30692));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n30691));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n30690));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n30689));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n30688));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n30687));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n30686));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n30685));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n30684));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n30683));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n30682));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i44684_2_lut_3_lut_4_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n1[1]));   // verilog/eeprom.v(68[25:39])
    defparam i44684_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(n44651), .O(n30106));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'ha8e8;
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(n69251), .D(state_7__N_3885[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 mux_1515_Mux_0_i3_3_lut_4_lut (.I0(state[0]), .I1(enable_slow_N_4213), 
            .I2(n25752), .I3(state[1]), .O(n5927[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1515_Mux_0_i3_3_lut_4_lut.LUT_INIT = 16'h04aa;
    SB_LUT4 add_1198_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5393[9]), 
            .I3(n59150), .O(delay_counter_15__N_3956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1198_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5393[9]), 
            .I3(n59149), .O(delay_counter_15__N_3956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_16 (.CI(n59149), .I0(delay_counter[14]), .I1(n5393[9]), 
            .CO(n59150));
    SB_LUT4 add_1198_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5393[9]), 
            .I3(n59148), .O(delay_counter_15__N_3956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_4_lut (.I0(state[2]), .I1(n15), .I2(n38017), .I3(data_ready), 
            .O(n29946));   // verilog/eeprom.v(27[11:16])
    defparam i12_4_lut_4_lut.LUT_INIT = 16'hfa08;
    SB_CARRY add_1198_15 (.CI(n59148), .I0(delay_counter[13]), .I1(n5393[9]), 
            .CO(n59149));
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n28091), .D(delay_counter_15__N_3956[15]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n28091), .D(delay_counter_15__N_3956[14]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n28091), .D(delay_counter_15__N_3956[12]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n28091), .D(delay_counter_15__N_3956[11]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n28091), .D(n6938), .S(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28091), 
            .D(n6937), .S(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28091), 
            .D(n6936), .S(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28091), 
            .D(n6935), .S(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28091), 
            .D(n6934), .S(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28091), 
            .D(delay_counter_15__N_3956[5]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28091), 
            .D(n6932), .S(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28091), 
            .D(delay_counter_15__N_3956[3]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28091), 
            .D(delay_counter_15__N_3956[2]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28091), 
            .D(delay_counter_15__N_3956[1]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1198_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5393[9]), 
            .I3(n59147), .O(delay_counter_15__N_3956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_14 (.CI(n59147), .I0(delay_counter[12]), .I1(n5393[9]), 
            .CO(n59148));
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28091), 
            .D(delay_counter_15__N_3956[0]), .R(n52961));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1198_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5393[9]), 
            .I3(n59146), .O(delay_counter_15__N_3956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_13 (.CI(n59146), .I0(delay_counter[11]), .I1(n5393[9]), 
            .CO(n59147));
    SB_LUT4 add_1198_12_lut (.I0(n52946), .I1(delay_counter[10]), .I2(n5393[9]), 
            .I3(n59145), .O(n6938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_12 (.CI(n59145), .I0(delay_counter[10]), .I1(n5393[9]), 
            .CO(n59146));
    SB_LUT4 add_1198_11_lut (.I0(n52946), .I1(delay_counter[9]), .I2(n5393[9]), 
            .I3(n59144), .O(n6937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_11 (.CI(n59144), .I0(delay_counter[9]), .I1(n5393[9]), 
            .CO(n59145));
    SB_LUT4 add_1198_10_lut (.I0(n52946), .I1(delay_counter[8]), .I2(n5393[9]), 
            .I3(n59143), .O(n6936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_10 (.CI(n59143), .I0(delay_counter[8]), .I1(n5393[9]), 
            .CO(n59144));
    SB_LUT4 add_1198_9_lut (.I0(n52946), .I1(delay_counter[7]), .I2(n5393[9]), 
            .I3(n59142), .O(n6935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_9 (.CI(n59142), .I0(delay_counter[7]), .I1(n5393[9]), 
            .CO(n59143));
    SB_LUT4 add_1198_8_lut (.I0(n52946), .I1(delay_counter[6]), .I2(n5393[9]), 
            .I3(n59141), .O(n6934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_8 (.CI(n59141), .I0(delay_counter[6]), .I1(n5393[9]), 
            .CO(n59142));
    SB_LUT4 add_1198_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5393[9]), 
            .I3(n59140), .O(delay_counter_15__N_3956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_7 (.CI(n59140), .I0(delay_counter[5]), .I1(n5393[9]), 
            .CO(n59141));
    SB_LUT4 add_1198_6_lut (.I0(n52946), .I1(delay_counter[4]), .I2(n5393[9]), 
            .I3(n59139), .O(n6932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_6 (.CI(n59139), .I0(delay_counter[4]), .I1(n5393[9]), 
            .CO(n59140));
    SB_LUT4 add_1198_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5393[9]), 
            .I3(n59138), .O(delay_counter_15__N_3956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_5 (.CI(n59138), .I0(delay_counter[3]), .I1(n5393[9]), 
            .CO(n59139));
    SB_LUT4 add_1198_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5393[9]), 
            .I3(n59137), .O(delay_counter_15__N_3956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_4 (.CI(n59137), .I0(delay_counter[2]), .I1(n5393[9]), 
            .CO(n59138));
    SB_LUT4 add_1198_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5393[9]), 
            .I3(n59136), .O(delay_counter_15__N_3956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_3 (.CI(n59136), .I0(delay_counter[1]), .I1(n5393[9]), 
            .CO(n59137));
    SB_LUT4 add_1198_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5393[9]), 
            .I3(GND_net), .O(delay_counter_15__N_3956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5393[9]), 
            .CO(n59136));
    SB_LUT4 i18_2_lut (.I0(state[2]), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n52946));
    defparam i18_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i62481_2_lut (.I0(n25752), .I1(enable_slow_N_4213), .I2(GND_net), 
            .I3(GND_net), .O(n5393[9]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i62481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(\state_7__N_3918[0] ), .O(n28163));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0908;
    SB_LUT4 i15218_3_lut_4_lut (.I0(n28163), .I1(state[2]), .I2(state[0]), 
            .I3(state[1]), .O(n29432));   // verilog/eeprom.v(68[25:39])
    defparam i15218_3_lut_4_lut.LUT_INIT = 16'h8aaa;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n61529));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i56327_3_lut (.I0(\state[0] ), .I1(n25752), .I2(state_adj_4449[3]), 
            .I3(GND_net), .O(n72174));
    defparam i56327_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n75328), .I1(n67746), .I2(state[0]), .I3(n72174), 
            .O(n17));
    defparam i24_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i2_4_lut_adj_956 (.I0(n17), .I1(state[2]), .I2(\state_7__N_3918[0] ), 
            .I3(state[1]), .O(n69251));
    defparam i2_4_lut_adj_956.LUT_INIT = 16'heefe;
    SB_LUT4 i38927_4_lut (.I0(state[1]), .I1(n15), .I2(state[2]), .I3(state[0]), 
            .O(state_7__N_3885[1]));   // verilog/eeprom.v(27[11:16])
    defparam i38927_4_lut.LUT_INIT = 16'ha5ba;
    SB_LUT4 i2_3_lut_4_lut (.I0(byte_counter[1]), .I1(n28), .I2(byte_counter[2]), 
            .I3(byte_counter[0]), .O(n125));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_3_lut_adj_957 (.I0(byte_counter[1]), .I1(n28), .I2(n66792), 
            .I3(GND_net), .O(n28274));
    defparam i1_2_lut_3_lut_adj_957.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_4_lut_adj_958 (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(n28), .I3(byte_counter[2]), .O(n117));   // verilog/eeprom.v(30[11:23])
    defparam i2_3_lut_4_lut_adj_958.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_959 (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(byte_counter[2]), .I3(GND_net), .O(n15));   // verilog/eeprom.v(30[11:23])
    defparam i1_2_lut_3_lut_adj_959.LUT_INIT = 16'he0e0;
    SB_LUT4 i16484_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[7]), 
            .I3(baudrate[15]), .O(n30698));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16484_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16486_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[6]), 
            .I3(baudrate[14]), .O(n30700));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16486_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16487_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[5]), 
            .I3(baudrate[13]), .O(n30701));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16487_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16488_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[4]), 
            .I3(baudrate[12]), .O(n30702));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16488_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16489_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[3]), 
            .I3(baudrate[11]), .O(n30703));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16489_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16490_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[2]), 
            .I3(baudrate[10]), .O(n30704));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16490_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16491_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[1]), 
            .I3(baudrate[9]), .O(n30705));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16491_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i59668_2_lut_3_lut (.I0(state_adj_4449[1]), .I1(state_adj_4449[2]), 
            .I2(state[1]), .I3(GND_net), .O(n75328));
    defparam i59668_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i16492_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[0]), 
            .I3(baudrate[8]), .O(n30706));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16492_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_960 (.I0(\state[0] ), .I1(state_adj_4449[3]), 
            .I2(n7), .I3(n25752), .O(n47));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut_adj_960.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_961 (.I0(\state[0] ), .I1(state_adj_4449[3]), 
            .I2(state_adj_4449[2]), .I3(state_adj_4449[1]), .O(n45262));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut_adj_961.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(state_adj_4449[1]), .I1(state_adj_4449[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/eeprom.v(55[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16473_3_lut_4_lut (.I0(state[2]), .I1(n125), .I2(data[2]), 
            .I3(baudrate[26]), .O(n30687));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16473_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16475_3_lut_4_lut (.I0(state[2]), .I1(n125), .I2(data[0]), 
            .I3(baudrate[24]), .O(n30689));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16475_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16470_3_lut_4_lut (.I0(state[2]), .I1(n125), .I2(data[5]), 
            .I3(baudrate[29]), .O(n30684));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16470_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16471_3_lut_4_lut (.I0(state[2]), .I1(n125), .I2(data[4]), 
            .I3(baudrate[28]), .O(n30685));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16471_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16472_3_lut_4_lut (.I0(state[2]), .I1(n125), .I2(data[3]), 
            .I3(baudrate[27]), .O(n30686));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16472_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i21372_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[7]), 
            .I3(ID[7]), .O(n30715));   // verilog/eeprom.v(35[8] 81[4])
    defparam i21372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16502_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[6]), 
            .I3(ID[6]), .O(n30716));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16503_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[5]), 
            .I3(ID[5]), .O(n30717));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16474_3_lut_4_lut (.I0(state[2]), .I1(n125), .I2(data[1]), 
            .I3(baudrate[25]), .O(n30688));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16474_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16504_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[4]), 
            .I3(ID[4]), .O(n30718));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16505_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[3]), 
            .I3(ID[3]), .O(n30719));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16506_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[2]), 
            .I3(ID[2]), .O(n30720));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16507_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[1]), 
            .I3(ID[1]), .O(n30721));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15731_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52949), .I2(data[0]), 
            .I3(ID[0]), .O(n29945));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15731_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut (.I0(ready_prev), .I1(n45262), .I2(state[0]), .I3(state[1]), 
            .O(n28));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i3_4_lut_adj_962 (.I0(state[2]), .I1(byte_counter[2]), .I2(byte_counter[0]), 
            .I3(n28), .O(n52949));   // verilog/eeprom.v(35[8] 81[4])
    defparam i3_4_lut_adj_962.LUT_INIT = 16'hfeff;
    SB_LUT4 i12_4_lut (.I0(delay_counter[10]), .I1(delay_counter[15]), .I2(delay_counter[8]), 
            .I3(delay_counter[14]), .O(n28_adj_4444));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[3]), .I2(delay_counter[7]), 
            .I3(delay_counter[1]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[2]), .I1(delay_counter[12]), .I2(delay_counter[6]), 
            .I3(delay_counter[5]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28_adj_4444), 
            .O(n25752));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_963 (.I0(state[0]), .I1(enable_slow_N_4213), .I2(n25752), 
            .I3(GND_net), .O(n60942));
    defparam i2_3_lut_adj_963.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(rw), .I2(n60942), .I3(state[2]), 
            .O(n10_adj_4445));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut.LUT_INIT = 16'h888a;
    SB_LUT4 i1_4_lut_adj_964 (.I0(n10_adj_4445), .I1(rw), .I2(state[0]), 
            .I3(state[2]), .O(n65940));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_adj_964.LUT_INIT = 16'heeae;
    SB_LUT4 i1_4_lut_adj_965 (.I0(n45262), .I1(saved_addr[0]), .I2(rw), 
            .I3(\state_7__N_4110[0] ), .O(n66328));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut_adj_965.LUT_INIT = 16'hd8cc;
    SB_LUT4 i44691_3_lut_4_lut (.I0(n44651), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n1[2]));   // verilog/eeprom.v(68[25:39])
    defparam i44691_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i1_3_lut_4_lut_4_lut_4_lut (.I0(state[2]), .I1(n15), .I2(state[0]), 
            .I3(state[1]), .O(n52961));
    defparam i1_3_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'h0052;
    SB_LUT4 i51939_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(state[1]), .I3(GND_net), .O(n67746));
    defparam i51939_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(state[2]), .I1(n15), .I2(state[0]), 
            .I3(state[1]), .O(n28091));
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h0552;
    i2c_controller i2c (.clk16MHz(clk16MHz), .scl_enable(scl_enable), .\state_7__N_4110[0] (\state_7__N_4110[0] ), 
            .sda_enable(sda_enable), .sda_out(sda_out), .GND_net(GND_net), 
            .n29970(n29970), .data({data}), .n29969(n29969), .n29967(n29967), 
            .n29966(n29966), .n29965(n29965), .n29961(n29961), .n29960(n29960), 
            .n66328(n66328), .\saved_addr[0] (saved_addr[0]), .n6707(n6707), 
            .\state[1] (state_adj_4449[1]), .\state[2] (state_adj_4449[2]), 
            .\state[3] (state_adj_4449[3]), .n30751(n30751), .n8(n8), 
            .VCC_net(VCC_net), .\state[0] (\state[0] ), .n11(n11), .enable_slow_N_4213(enable_slow_N_4213), 
            .n7(n7), .\state_7__N_4126[3] (\state_7__N_4126[3] ), .enable(enable), 
            .n44639(n44639), .n10(n10), .n4(n4), .n4_adj_1(n4_adj_2), 
            .n25890(n25890), .n25932(n25932), .n44782(n44782), .scl(scl)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (clk16MHz, scl_enable, \state_7__N_4110[0] , sda_enable, 
            sda_out, GND_net, n29970, data, n29969, n29967, n29966, 
            n29965, n29961, n29960, n66328, \saved_addr[0] , n6707, 
            \state[1] , \state[2] , \state[3] , n30751, n8, VCC_net, 
            \state[0] , n11, enable_slow_N_4213, n7, \state_7__N_4126[3] , 
            enable, n44639, n10, n4, n4_adj_1, n25890, n25932, 
            n44782, scl) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output scl_enable;
    output \state_7__N_4110[0] ;
    output sda_enable;
    output sda_out;
    input GND_net;
    input n29970;
    output [7:0]data;
    input n29969;
    input n29967;
    input n29966;
    input n29965;
    input n29961;
    input n29960;
    input n66328;
    output \saved_addr[0] ;
    output n6707;
    output \state[1] ;
    output \state[2] ;
    output \state[3] ;
    input n30751;
    input n8;
    input VCC_net;
    output \state[0] ;
    output n11;
    output enable_slow_N_4213;
    input n7;
    input \state_7__N_4126[3] ;
    input enable;
    output n44639;
    output n10;
    output n4;
    output n4_adj_1;
    output n25890;
    output n25932;
    output n44782;
    output scl;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire i2c_clk_N_4199, scl_enable_N_4200, enable_slow_N_4212, n28151, 
        sda_out_adj_4430;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n29410;
    wire [7:0]n119;
    
    wire n28226;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n29179, n5, n45195, n44936, n45193, n69903, n69684, n59157, 
        n59156, n59155, n59154, n59153, n59152, n59151, n68919, 
        n28145, n66042, n69020, n28143, n11_adj_4431, n15, n11_adj_4432, 
        n60333, n60332, n60331, n60330, n60329, n28, n78295, n11_adj_4433, 
        n67720;
    wire [1:0]n6776;
    
    wire n11_adj_4434, n4_c, n6700, n44732, n9, n12, n4_adj_4435, 
        n75329, n7044, n10_adj_4436, n9_adj_4438;
    
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4199));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4200));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4110[0] ), .C(clk16MHz), .E(n28151), 
            .D(enable_slow_N_4212));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i2555_2_lut (.I0(sda_out_adj_4430), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2555_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29970));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29969));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29966));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29965));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29961));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29960));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n66328));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2057_2058__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29410));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29410));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29410));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29410));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29410));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n28226), .D(n119[1]), 
            .S(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n28226), .D(n119[2]), 
            .S(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n28226), .D(n119[3]), 
            .R(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n28226), .D(n119[4]), 
            .R(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n28226), .D(n119[5]), 
            .R(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n28226), .D(n119[6]), 
            .R(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n28226), .D(n119[7]), 
            .R(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6707), .D(n5), 
            .S(n45195));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6707), .D(n44936), 
            .S(n45193));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6707), .D(n69903), 
            .S(n69684));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2057_2058__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29410));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30751));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i62494_2_lut (.I0(enable_slow_N_4213), .I1(\state_7__N_4110[0] ), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4212));   // verilog/i2c_controller.v(44[32:47])
    defparam i62494_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n59157), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n59156), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n59156), .I0(counter[6]), .I1(VCC_net), 
            .CO(n59157));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n59155), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n59155), .I0(counter[5]), .I1(VCC_net), 
            .CO(n59156));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n59154), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n59154), .I0(counter[4]), .I1(VCC_net), 
            .CO(n59155));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n59153), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n59153), .I0(counter[3]), .I1(VCC_net), 
            .CO(n59154));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n59152), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n59152), .I0(counter[2]), .I1(VCC_net), 
            .CO(n59153));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n59151), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n59151), .I0(counter[1]), .I1(VCC_net), 
            .CO(n59152));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n59151));
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n28145), 
            .D(n68919), .S(n66042));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4430), .C(i2c_clk), .E(n28143), 
            .D(n69020), .S(n66042));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n28226), .D(n119[0]), 
            .S(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i52016_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(scl_enable_N_4200));
    defparam i52016_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4431));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n15));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4432));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 counter2_2057_2058_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n60333), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2057_2058_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n60332), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_6 (.CI(n60332), .I0(GND_net), .I1(counter2[4]), 
            .CO(n60333));
    SB_LUT4 counter2_2057_2058_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n60331), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_5 (.CI(n60331), .I0(GND_net), .I1(counter2[3]), 
            .CO(n60332));
    SB_LUT4 counter2_2057_2058_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n60330), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_4 (.CI(n60330), .I0(GND_net), .I1(counter2[2]), 
            .CO(n60331));
    SB_LUT4 counter2_2057_2058_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n60329), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_3 (.CI(n60329), .I0(GND_net), .I1(counter2[1]), 
            .CO(n60330));
    SB_LUT4 counter2_2057_2058_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n60329));
    SB_LUT4 i14965_2_lut_4_lut (.I0(n28226), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n29179));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14965_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5110;
    SB_LUT4 i62439_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n78295));
    defparam i62439_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_944 (.I0(n11_adj_4433), .I1(n78295), .I2(n28), 
            .I3(n67720), .O(n28143));
    defparam i1_4_lut_adj_944.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1830_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6776[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1830_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i31282_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n67720));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i31282_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(\state[0] ), .I1(n7), .I2(\state[3] ), .I3(n11_adj_4433), 
            .O(n66042));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_945 (.I0(n11_adj_4433), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n67720), .O(n28145));
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h0a22;
    SB_LUT4 i1_4_lut_adj_946 (.I0(\state_7__N_4126[3] ), .I1(n11_adj_4434), 
            .I2(n11_adj_4433), .I3(enable), .O(n4_c));
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h2a2f;
    SB_LUT4 i62976_3_lut (.I0(n6707), .I1(n15), .I2(n11), .I3(GND_net), 
            .O(n45193));
    defparam i62976_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i62928_2_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_4434), 
            .I2(GND_net), .I3(GND_net), .O(n44936));
    defparam i62928_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i62977_4_lut (.I0(n6707), .I1(\state[0] ), .I2(n11_adj_4431), 
            .I3(n7), .O(n45195));
    defparam i62977_4_lut.LUT_INIT = 16'h0a8a;
    SB_LUT4 i62464_4_lut (.I0(\state[3] ), .I1(n6700), .I2(n44732), .I3(n44639), 
            .O(n6707));
    defparam i62464_4_lut.LUT_INIT = 16'h5f13;
    SB_LUT4 i1_4_lut_adj_947 (.I0(n11_adj_4432), .I1(n11_adj_4434), .I2(\saved_addr[0] ), 
            .I3(\state_7__N_4126[3] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h5575;
    SB_LUT4 equal_276_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_276_i9_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6700));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(\state[3] ), .I1(n6700), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4435));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i59669_4_lut (.I0(n7), .I1(n4_adj_4435), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n75329));
    defparam i59669_4_lut.LUT_INIT = 16'hfcdd;
    SB_LUT4 i14_4_lut (.I0(n75329), .I1(n9), .I2(n7044), .I3(\state_7__N_4126[3] ), 
            .O(n28226));
    defparam i14_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i30551_3_lut_4_lut_4_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n44639));   // verilog/i2c_controller.v(151[5:14])
    defparam i30551_3_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'hfcfd;
    SB_LUT4 i62972_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6707), 
            .I3(\state[1] ), .O(n69684));   // verilog/i2c_controller.v(151[5:14])
    defparam i62972_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 equal_1562_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4433));   // verilog/i2c_controller.v(151[5:14])
    defparam equal_1562_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4434));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i62491_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(44[32:47])
    defparam i62491_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n7044));   // verilog/i2c_controller.v(44[32:47])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6776[1]), 
            .I3(\state[1] ), .O(n69020));   // verilog/i2c_controller.v(44[32:47])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4436));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4436), .I2(counter2[0]), 
            .I3(GND_net), .O(n29410));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_948 (.I0(i2c_clk), .I1(n29410), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_4199));
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_949 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n68919));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_949.LUT_INIT = 16'h1110;
    SB_LUT4 i1_2_lut_3_lut_adj_950 (.I0(enable), .I1(enable_slow_N_4213), 
            .I2(\state_7__N_4110[0] ), .I3(GND_net), .O(n28151));
    defparam i1_2_lut_3_lut_adj_950.LUT_INIT = 16'hbaba;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_355_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_355_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i30643_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(GND_net), .O(n44732));
    defparam i30643_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2_3_lut_4_lut_adj_951 (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_c), 
            .I3(n9_adj_4438), .O(n69903));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut_adj_951.LUT_INIT = 16'hf0f4;
    SB_LUT4 equal_353_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_353_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_952 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n25890));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_952.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4438));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_953 (.I0(n15), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_953.LUT_INIT = 16'hbbbb;
    SB_LUT4 i30693_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n44782));
    defparam i30693_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30585_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i30585_2_lut.LUT_INIT = 16'hbbbb;
    
endmodule
