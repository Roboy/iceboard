// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Jan 29 13:09:37 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    output SCL;   // verilog/TinyFPGA_B.v(21[10:13])
    input SDA /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, CLK_c, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, n4, 
        INHC_c, INLB_c, INHB_c, INLA_c, INHA_c;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(42[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(88[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(89[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(123[22:39])
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(124[21:45])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(125[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(126[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(127[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(128[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(129[22:24])
    
    wire n25358;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(131[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(132[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(133[22:35])
    
    wire n25228, n15590, n25357, n25227;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(163[22:33])
    wire [22:0]pwm_setpoint_22__N_3;
    
    wire RX_N_2;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [31:0]motor_state_23__N_74;
    wire [25:0]encoder0_position_scaled_23__N_26;
    wire [23:0]displacement_23__N_50;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n25356, n21945;
    wire [3:0]state_3__N_272;
    
    wire n25355, n25354, n2329, n25353, n4218, n25226, n25352, 
        n4216, n35368, n25351, n25225, n25350, n25349, n25348, 
        n445, n444, n443, n442, n441, n440, n439, n438, n437, 
        n436, n435, n434, n433, n432, n431, n430, n429, n428, 
        n427, n426, n425, n16911, n16910;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n25347, n3, n4_adj_4488, n5, n6, n7, n8, n9, n10, 
        n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
        n21, n22, n23, n24, n25, n25346, n25345, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n25224, n25344, n25343, n25223, n25222;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    
    wire n25342, n25341, tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n122, n25221, n8_adj_4489, n35073, n8868, n34025, n34029, 
        n33957, n24_adj_4490, n21_adj_4491, n20_adj_4492, n17_adj_4493, 
        n33976, n16909, n16908, n16907, n16906, n16905, n16904, 
        n16903, n16902, n16901, n16900, n16899, n16898, n16897, 
        n16896, n16894, n16893, n16892, n16891, n16890, n16889, 
        n16888, n16887, n16886, n25340, n4_adj_4494, n32219, n33956, 
        n771, n33876, n33874, n33856, n33850, n33848, n25339, 
        n25338, n25220, n25337, n25219, n25336, n25335, n25218, 
        n25217, n25334, n25216, n25333, n25332, n25215, n25331, 
        n25214, n25213, n25212, n25211, n25330, n25329, n25210, 
        n25328, n22115, n25327, n25326, n25209, n25325, n25208, 
        n25324, n25207, n25323, n25322, n25206, n25321, n25320, 
        n25205, n25319, n21885, n25204, n25203, n25202, n25201, 
        n25318, n25200, n25199, n25198, n25317, n25316, n25197, 
        n25315, n25314, n25313, n25196, n25312, n25195, n21796, 
        n25311, n25310, n25194, n25193, n25309, n33540, n25192, 
        n25191, n25308, n25307, n25190, n25189, n25306, n25305, 
        n25304, n25188, n25187, n21215, n25303, n25186, n25185, 
        n25302, n33530, n25301, n25300, n21989, n25299, n25184, 
        n25298, n25183, n25297, n25182, n25296, n25181, n25180, 
        n25295, n5_adj_4495, n30808, n25179, n25294, n25178, n22097, 
        n25293, n25292, n16885, n16884, n25291, n4452, n25177, 
        n25176, n22035, n25290, n25289, n78, n25288, n31590, n14_adj_4496, 
        n9_adj_4497, n25175, n25287, n25174, n25173, n25172, n25286, 
        n25171, n24951, n24950, n25285, n24949, n25170, n24948, 
        n25284, n25283, n18701, n28583, n33807, n25169, n33723, 
        n33247, n33241, n25168, n33725, \FRAME_MATCHER.i_31__N_2364 , 
        n25167, \FRAME_MATCHER.i_31__N_2370 , n33239, n33235, n33233, 
        n17382, n17381, n17380, n17376, n17373, n17372, n17371, 
        n17370, n17369, n17368, n17367, n17366, n17365, n17364, 
        n17363, n17362, n17361, n17360, n17359, n17358, n17357, 
        n17356, n17355, n17354, n17353, n17352, n17351, n17350, 
        n17349, n17348, n17347, n17346, n17345, n17344, n17343, 
        n17342, n17341, n17340, n17339, n17338, n17337, n17336, 
        n17335, n17334, n17333, n17332, n17331, n17330, n17329, 
        n17328, n17327, n17326, n17325, n17324, n17323, n17322, 
        n17321, n17320, n17316, n17314, n17313, n17312, n17311, 
        n17310, n17309, n17308, n17307, n17306, n17305, n17304, 
        n17303, n17302, n17301, n17300, n17299, n17298, n17297, 
        n17296, n17295, n17294, n17293, n17292, n17291, n17290, 
        n17289, n17288, n17287, n17286, n17285, n17284, n17283, 
        n17282, n17281, n17280, n17279, n17278, n17277, n17276, 
        n17275, n17274, n17273, n17272, n17271, n17270, n17269, 
        n17268, n17267, n17266, n17265, n17264, n17263, n17262, 
        n17261, n17260, n17259, n17258, n17257, n17256, n17255, 
        n17254, n17253, n17252, n17251, n17250, n17249, n17248, 
        n17247, n17246, n17245, n17244, n17243, n17242, n17241, 
        n17240, n17239, n5_adj_4498, n17238, n17237, n17236, n17235, 
        n17234, n17233, n17232, n17231, n17230, n17229, n17228, 
        n17227, n17226, n17225, n17224, n17223, n17222, n17221, 
        n17220, n17219, n17218, n17217, n17216, n17215, n17214, 
        n17213, n17212, n17211, n17210, n17209, n17208, n17207, 
        n17206, n17205, n17204, n17203, n17202, n30284, n17201, 
        n17200, n17199, n17198, n17197, n17196, n17195, n17194, 
        n17193, n17192, n17191, n17190, n17189, n17188, n17187, 
        n17186, n17185, n17184, n17183, n17182, n17181, n17180, 
        n17179, n17178, n17177, n17176, n17175, n17174, n17173, 
        n17172, n17171, n17170, n17169, n17168, n17167, n17166, 
        n17165, n17164, n17163, n17162, n17161, n17160, n17159, 
        n17158, n17157, n17156, n17155, n17154, n17153, n17152, 
        n17151, n17150, n17149, n17148, n17147, n17146, n17145, 
        n17144, n17143, n17142, n17141, n17140, n17139, n17138, 
        n17137, n17136, n17135, n17134, n17133, n17132, n26, n24_adj_4499, 
        n22_adj_4500, n31097, n18_adj_4501, n7_adj_4502, n17131, n33199, 
        n63, n17130, n17129, n17128, n17127, n17126, n17125, n17124, 
        n17123, n17122, n17121, n25282, n24947, n25166, n24946, 
        n25165, n31395, n25281, n25164, n24945, n25163, n24944, 
        n25162, n25421, n25280, n25420, n25279, n25161, n25419, 
        n25160, n24943;
    wire [23:0]duty_23__N_3516;
    
    wire quadA_debounced, quadB_debounced, n25278, n24942, n17120, 
        n25_adj_4503, n17119, quadA_debounced_adj_4504, quadB_debounced_adj_4505, 
        n17118, n17117, n25159, n17116, n25158, n24_adj_4506, n23_adj_4507, 
        n22_adj_4508, n21_adj_4509, n20_adj_4510, n19_adj_4511, n18_adj_4512, 
        n17_adj_4513, n16_adj_4514, n15_adj_4515, n14_adj_4516, n13_adj_4517, 
        n12_adj_4518, n11_adj_4519, n10_adj_4520, n9_adj_4521, n8_adj_4522, 
        n7_adj_4523, n6_adj_4524, n5_adj_4525, n4_adj_4526, n3_adj_4527, 
        n2, n17115, n24941, n25418, n25417, n22083, n17114, n25277, 
        n17113, n25276, n17112, n17111, n17110, n17109, n17108, 
        n17107, n17106, n17105, n17104, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n25416, n25275, n17103, n17102, n5_adj_4528, n17101, n17100, 
        n25076, n25075, n17099, n17098, n17097, n17096, n24940, 
        n25157, n17095, n17094, n17093, n17092, n17091, n17090, 
        n17089, n25074, n25073, n25274, n25156, n25273, n15_adj_4529, 
        n25155, n25415, n24939, n25272, n22075, n25154, n4_adj_4530, 
        n17088, n17087, n17086, n17085, n17084, n25414, n17083, 
        n17082, n17081, n17080, n17079;
    wire [2:0]r_SM_Main_adj_4704;   // verilog/uart_tx.v(31[16:25])
    
    wire n25271, n25270, n25413, n22053, n25412, n25153, n25269, 
        n25411, n25268, n25267, n15_adj_4531;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n25072, n3_adj_4532;
    wire [1:0]reg_B_adj_4715;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n25410, n17031, n17030, n17029, n17028, n17027, n17026, 
        n17025, n17024, n17023, n17022, n17021, n17020, n17019, 
        n17018, n17017, n17016, n25409, n4_adj_4535, n6_adj_4536, 
        n7_adj_4537, n8_adj_4538, n9_adj_4539, n10_adj_4540, n11_adj_4541, 
        n12_adj_4542, n13_adj_4543, n14_adj_4544, n15_adj_4545, n16_adj_4546, 
        n17_adj_4547, n18_adj_4548, n19_adj_4549, n20_adj_4550, n21_adj_4551, 
        n22_adj_4552, n23_adj_4553, n24_adj_4554, n25_adj_4555, n509, 
        n510, n511, n20_adj_4556, n18_adj_4557, n16_adj_4558, n619, 
        n29535, n34030, n25152, n674, n675, n676, n677, n678, 
        n679, n700, n4431, n4432, n4433, n4434, n728, n729, 
        n730, n731, n732, n733, n752, n753, n754, n755, n756, 
        n757, n758, n778, n33173, n806, n807, n808, n809, n810, 
        n811, n812, n830, n831, n832, n833, n834, n835, n836, 
        n837, n8_adj_4559, n856, n7_adj_4560, n34, n883, n884, 
        n885, n886, n887, n888, n889, n890, n891, n908, n909, 
        n910, n911, n912, n913, n914, n915, n916, n934, n31, 
        n961, n962, n963, n964, n965, n966, n967, n968, n969, 
        n970, n30, n28, n986, n987, n988, n989, n990, n991, 
        n992, n993, n994, n995, n1012, n1039, n1040, n1041, 
        n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
        n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
        n1072, n1073, n1074, n1090, n22_adj_4561, n21_adj_4562, 
        n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
        n1125, n1126, n1127, n1128, n1142, n1143, n1144, n1145, 
        n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
        n25408, n1168, n1195, n1196, n1197, n1198, n1199, n1200, 
        n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1220, 
        n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
        n1229, n1230, n1231, n1232, n1246, n1273, n1274, n1275, 
        n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
        n1284, n1285, n1286, n1298, n1299, n1300, n1301, n1302, 
        n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
        n1311, n25071, n1324, n1351, n1352, n1353, n1354, n1355, 
        n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
        n1364, n1365, n1376, n1377, n1378, n1379, n1380, n1381, 
        n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
        n1390, n34194, n1402, n1429, n1430, n1431, n1432, n1433, 
        n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
        n1442, n1443, n1444, n1454, n1455, n1456, n1457, n1458, 
        n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
        n1467, n1468, n1469, n1480, n1507, n1508, n1509, n1510, 
        n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
        n1519, n1520, n1521, n1522, n1523, n1532, n1533, n1534, 
        n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
        n1543, n1544, n1545, n1546, n1547, n1548, n1558, n1585, 
        n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
        n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, 
        n1602, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
        n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, 
        n1625, n1626, n1627, n1636, n1663, n1664, n1665, n1666, 
        n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, 
        n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1688, 
        n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
        n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
        n1705, n1706, n1714, n1741, n1742, n1743, n1744, n1745, 
        n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, 
        n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1766, 
        n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
        n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
        n1783, n1784, n1785, n1792, n1819, n1820, n1821, n1822, 
        n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
        n1839, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
        n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
        n1859, n1860, n1861, n1862, n1863, n1864, n1870, n1897, 
        n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
        n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, 
        n1914, n1915, n1916, n1917, n1918, n1922, n1923, n1924, 
        n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
        n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
        n1941, n1942, n1943, n1948, n1975, n1976, n1977, n1978, 
        n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
        n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
        n1995, n1996, n1997, n2000, n2001, n2002, n2003, n2004, 
        n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
        n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
        n2021, n2022, n2026, n2053, n2054, n2055, n2056, n2057, 
        n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
        n2066, n2067, n2068, n2069, n2070, n2071, n2073, n2076, 
        n22095, n4680, n4679, n4678, n4677, n4676, n4675, n4674, 
        n4673, n4672, n4671, n4670, n4669, n4668, n4667, n4666, 
        n4665, n4664, n4663, n4662, n4660, n4659, n15455, n34_adj_4563, 
        n25907, n25906, n33, n25905, n33869, n25904, n25903, n32, 
        n25266, n16802, n16710, n31_adj_4564, n16698, n25902, n30_adj_4565, 
        n63_adj_4566, n28077, n16882, n16881, n28495, n15545, n16880, 
        n16879, n16878, n16877, n16876, n16875, n33155, n33154, 
        n29, n4_adj_4567, n6_adj_4568, n7_adj_4569, n8_adj_4570, n9_adj_4571, 
        n10_adj_4572, n11_adj_4573, n12_adj_4574, n13_adj_4575, n15_adj_4576, 
        n17_adj_4577, n19_adj_4578, n21_adj_4579, n33875, n23_adj_4580, 
        n25_adj_4581, n27, n33873, n29_adj_4582, n30_adj_4583, n31_adj_4584, 
        n33_adj_4585, n35, n29542, n25407, n25406, n34028, n4429, 
        n25070, n26_adj_4586, n25_adj_4587, n24_adj_4588, n23_adj_4589, 
        n25405, n24938, n25265, n25264, n5_adj_4590, n33773, n25069, 
        n16967, n16966, n16965, n16964, n16963, n16962, n16961, 
        n16960, n16959, n16958, n16957, n16956, n16955, n16954, 
        n16953, n16874, n16872, n16871, n16870, n16867, n16952, 
        n16865, n16864, n16863, n16862, n16861, n16860, n16859, 
        n16858, n16935, n16934, n16933, n16932, n16931, n16930, 
        n16929, n16928, n30717, n31908, n30785, n29538, n25263, 
        n24937, n25404, n24936, n34057, n2_adj_4591, n3_adj_4592, 
        n4_adj_4593, n5_adj_4594, n6_adj_4595, n7_adj_4596, n8_adj_4597, 
        n9_adj_4598, n10_adj_4599, n11_adj_4600, n12_adj_4601, n13_adj_4602, 
        n14_adj_4603, n15_adj_4604, n16_adj_4605, n17_adj_4606, n18_adj_4607, 
        n19_adj_4608, n20_adj_4609, n21_adj_4610, n22_adj_4611, n23_adj_4612, 
        n24_adj_4613, n25_adj_4614, n25262, n34501, n29539, n25068, 
        n25261, n25403, n25402, n33120, n33118, n7_adj_4615, n13_adj_4616, 
        n23_adj_4617, n27_adj_4618, n29_adj_4619, n37, n39, n43, 
        n45, n49, n25067, n8_adj_4620, n7_adj_4621, n17_adj_4622, 
        n16_adj_4623, n25260, n25401, n8947, n24935, n24934, n22021, 
        n25400, n25399, n25259, n25258, n25151, n25066, n25150, 
        n25149, n16857, n25729, n30832, n30290, n30288, n30286, 
        n16856, n30267, n6_adj_4624, n25728, n25727, n4_adj_4625, 
        n25257, n12869, n29497, n25726, n25725, n25724, n31108, 
        n28_adj_4626, n27_adj_4627, n29541, n26_adj_4628, n25_adj_4629, 
        n25723, n25722, n25398, n30_adj_4630, n25721, n25720, n29_adj_4631, 
        n28_adj_4632, n27_adj_4633, n18_adj_4634, n25719, n25718, 
        n25717, n25716, n25715, n25714, n25713, n25712, n25711, 
        n25710, n25397, n25148, n25065, n25396, n25064, n25395, 
        n25709, n25708, n24933, n25256, n25255, n25707, n25706, 
        n16_adj_4635, n12_adj_4636, n10_adj_4637, n25394, n31065, 
        n2_adj_4638, n16855, n25393, n25392, n16853, n25254, n16852, 
        n5_adj_4639, n28937, n4_adj_4640, n25253, n32056, n37_adj_4641, 
        n36, n30_adj_4642, n25391, n25390, n25147, n29_adj_4643, 
        n28_adj_4644, n27_adj_4645, n26_adj_4646, n25_adj_4647, n25389, 
        n25388, n25387, n24_adj_4648, n25252, n23_adj_4649, n22_adj_4650, 
        n21_adj_4651, n25063, n24932, n25386, n25146, n25385, n31461, 
        n15450, n15595, n25384, n25145, n25251, n25383, n25382, 
        n25381, n10_adj_4652, n25380, n25062, n25379, n25378, n25377, 
        n22009, n25250, n29532, n25249, n25376, n25248, n25375, 
        n24931, n24930, n22007, n25374, n24929, n25373, n25247, 
        n25372, n25371, n25370, n25246, n12944, n25245, n25244, 
        n25061, n25243, n24928, n22003, n25369, n24927, n25060, 
        n25059, n25242, n25241, n25368, n24926, n22001, n25240, 
        n25239, n25058, n25367, n25238, n25237, n25236, n25366, 
        n25235, n25057, n25365, n25234, n25364, n25233, n25232, 
        n21971, n25231, n25363, n25230, n25056, n14_adj_4653, n10_adj_4654, 
        n22023, n25362, n24925, n25055, n22055, n25361, n25360, 
        n25054, n22041, n12_adj_4655, n15453, n25359, n6_adj_4656, 
        n22057, n6_adj_4657, n25229, n31883;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .data_o({quadA_debounced, quadB_debounced}), 
            .clk32MHz(clk32MHz), .n31883(n31883), .reg_B({reg_B}), .VCC_net(VCC_net), 
            .n16870(n16870), .ENCODER0_B_c_0(ENCODER0_B_c_0), .n17381(n17381), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(186[15] 191[4])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_28 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_50[0]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h2_27 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .GND_net(GND_net), .VCC_net(VCC_net), 
            .timer({timer}), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .\state_3__N_272[1] (state_3__N_272[1]), .start(start), .LED_c(LED_c), 
            .\state[0] (state[0]), .n21971(n21971), .\state[1] (state[1]), 
            .n22115(n22115), .neopxl_color({neopxl_color}), .n16698(n16698), 
            .n30267(n30267), .n28583(n28583), .n28495(n28495), .n17366(n17366), 
            .n17365(n17365), .n17364(n17364), .n17363(n17363), .n17362(n17362), 
            .n17361(n17361), .n17360(n17360), .n17359(n17359), .n17358(n17358), 
            .n17357(n17357), .n17356(n17356), .n17355(n17355), .n17354(n17354), 
            .n17353(n17353), .n17352(n17352), .n17351(n17351), .n17350(n17350), 
            .n17349(n17349), .n17348(n17348), .n17347(n17347), .n17346(n17346), 
            .n17345(n17345), .n17344(n17344), .n17343(n17343), .n17342(n17342), 
            .n17341(n17341), .n17340(n17340), .n17339(n17339), .n17338(n17338), 
            .n17337(n17337), .n17336(n17336), .n17316(n17316), .NEOPXL_c(NEOPXL_c), 
            .n16852(n16852)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(44[10] 50[2])
    SB_CARRY encoder0_position_23__I_0_add_566_6 (.CI(n25155), .I0(n834), 
            .I1(GND_net), .CO(n25156));
    SB_DFF dir_32 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 encoder0_position_23__I_0_add_566_5_lut (.I0(GND_net), .I1(n835), 
            .I2(VCC_net), .I3(n25154), .O(n888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_41_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[7]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_i1373_3_lut (.I0(n2010), .I1(n2063), 
            .I2(n2026), .I3(GND_net), .O(n29_adj_4619));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1374_3_lut (.I0(n2011), .I1(n2064), 
            .I2(n2026), .I3(GND_net), .O(n27_adj_4618));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1365_3_lut (.I0(n2002), .I1(n2055), 
            .I2(n2026), .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1381_3_lut (.I0(n2018), .I1(n2071), 
            .I2(n2026), .I3(GND_net), .O(n13_adj_4616));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1368_3_lut (.I0(n2005), .I1(n2058), 
            .I2(n2026), .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut (.I0(n2020), .I1(n33199), .I2(n2026), .I3(n2019), 
            .O(n5_adj_4495));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i27811_3_lut (.I0(n445), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n33154));
    defparam i27811_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 encoder0_position_23__I_0_i1363_3_lut (.I0(n2000), .I1(n2053), 
            .I2(n2026), .I3(GND_net), .O(n49));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1366_3_lut (.I0(n2003), .I1(n2056), 
            .I2(n2026), .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_41_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[22]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut (.I0(n33154), .I1(n5_adj_4495), .I2(n33155), .I3(n2026), 
            .O(n28077));
    defparam i1_4_lut.LUT_INIT = 16'h88c0;
    SB_CARRY encoder0_position_23__I_0_add_566_5 (.CI(n25154), .I0(n835), 
            .I1(VCC_net), .CO(n25155));
    SB_LUT4 i4_4_lut (.I0(n2016), .I1(n29_adj_4619), .I2(n2069), .I3(n2026), 
            .O(n24_adj_4648));
    defparam i4_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i4_4_lut_adj_1616 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4652));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i4_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4652), .I2(control_mode[2]), 
            .I3(GND_net), .O(n15545));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut (.I0(n28077), .I1(n2001), .I2(n2054), .I3(n2026), 
            .O(n22_adj_4650));
    defparam i2_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i3_4_lut (.I0(n2007), .I1(n49), .I2(n2060), .I3(n2026), 
            .O(n23_adj_4649));
    defparam i3_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i1_2_lut (.I0(n15450), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4531));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_1617 (.I0(n2014), .I1(n43), .I2(n2067), .I3(n2026), 
            .O(n21_adj_4651));
    defparam i1_4_lut_adj_1617.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_23__I_0_i1369_3_lut (.I0(n2006), .I1(n2059), 
            .I2(n2026), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n15545), 
            .I3(GND_net), .O(n15_adj_4529));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_41_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[23]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4555));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1376_3_lut (.I0(n2013), .I1(n2066), 
            .I2(n2026), .I3(GND_net), .O(n23_adj_4617));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_4_lut (.I0(n2008), .I1(n27_adj_4618), .I2(n2061), .I3(n2026), 
            .O(n28_adj_4644));
    defparam i8_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i6_4_lut (.I0(n2004), .I1(n45), .I2(n2057), .I3(n2026), 
            .O(n26_adj_4646));
    defparam i6_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i7_4_lut (.I0(n2012), .I1(n13_adj_4616), .I2(n2065), .I3(n2026), 
            .O(n27_adj_4645));
    defparam i7_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i5_4_lut (.I0(n2017), .I1(n23_adj_4617), .I2(n2070), .I3(n2026), 
            .O(n25_adj_4647));
    defparam i5_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4554));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut (.I0(n2009), .I1(n39), .I2(n2062), .I3(n2026), 
            .O(n30_adj_4642));
    defparam i10_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i16_4_lut_adj_1618 (.I0(n21_adj_4651), .I1(n23_adj_4649), .I2(n22_adj_4650), 
            .I3(n24_adj_4648), .O(n36));
    defparam i16_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n2015), .I1(n37), .I2(n2068), .I3(n2026), 
            .O(n29_adj_4643));
    defparam i9_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i17_4_lut (.I0(n25_adj_4647), .I1(n27_adj_4645), .I2(n26_adj_4646), 
            .I3(n28_adj_4644), .O(n37_adj_4641));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28752_4_lut (.I0(n37_adj_4641), .I1(n29_adj_4643), .I2(n36), 
            .I3(n30_adj_4642), .O(n22055));
    defparam i28752_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4540), .I3(n25068), .O(displacement_23__N_50[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_41_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[8]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_41_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[9]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_41_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[10]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4553));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4552));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4551));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4550));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n25068), .I0(encoder1_position[15]), 
            .I1(n10_adj_4540), .CO(n25069));
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4541), .I3(n25067), .O(displacement_23__N_50[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_41_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[11]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_add_566_4_lut (.I0(GND_net), .I1(n836), 
            .I2(GND_net), .I3(n25153), .O(n889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_4 (.CI(n25153), .I0(n836), 
            .I1(GND_net), .CO(n25154));
    SB_LUT4 encoder0_position_23__I_0_add_566_3_lut (.I0(GND_net), .I1(n837), 
            .I2(VCC_net), .I3(n25152), .O(n890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_3 (.CI(n25152), .I0(n837), 
            .I1(VCC_net), .CO(n25153));
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_566_2_lut (.I0(GND_net), .I1(n430), 
            .I2(GND_net), .I3(VCC_net), .O(n891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_2 (.CI(VCC_net), .I0(n430), 
            .I1(GND_net), .CO(n25152));
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12790_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4216), .I3(GND_net), .O(n16899));   // verilog/coms.v(127[12] 300[6])
    defparam i12790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_513_9_lut (.I0(n34194), .I1(n752), 
            .I2(VCC_net), .I3(n25151), .O(n830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12907_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n29539), 
            .I3(GND_net), .O(n17016));   // verilog/coms.v(127[12] 300[6])
    defparam i12907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12791_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4216), .I3(GND_net), .O(n16900));   // verilog/coms.v(127[12] 300[6])
    defparam i12791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_513_8_lut (.I0(GND_net), .I1(n753), 
            .I2(VCC_net), .I3(n25150), .O(n806)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12908_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n29539), 
            .I3(GND_net), .O(n17017));   // verilog/coms.v(127[12] 300[6])
    defparam i12908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12909_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n29539), 
            .I3(GND_net), .O(n17018));   // verilog/coms.v(127[12] 300[6])
    defparam i12909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12910_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n29539), 
            .I3(GND_net), .O(n17019));   // verilog/coms.v(127[12] 300[6])
    defparam i12910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12911_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n29539), 
            .I3(GND_net), .O(n17020));   // verilog/coms.v(127[12] 300[6])
    defparam i12911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12912_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n29539), 
            .I3(GND_net), .O(n17021));   // verilog/coms.v(127[12] 300[6])
    defparam i12912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_41_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[12]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_23__I_0_add_513_8 (.CI(n25150), .I0(n753), 
            .I1(VCC_net), .CO(n25151));
    SB_LUT4 i12913_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n29539), 
            .I3(GND_net), .O(n17022));   // verilog/coms.v(127[12] 300[6])
    defparam i12913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12792_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4216), .I3(GND_net), .O(n16901));   // verilog/coms.v(127[12] 300[6])
    defparam i12792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_41_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[13]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12914_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n29539), 
            .I3(GND_net), .O(n17023));   // verilog/coms.v(127[12] 300[6])
    defparam i12914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut (.I0(pwm_counter[27]), .I1(pwm_counter[28]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4654));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1619 (.I0(pwm_counter[23]), .I1(pwm_counter[29]), 
            .I2(pwm_counter[25]), .I3(pwm_counter[26]), .O(n14_adj_4653));
    defparam i6_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1620 (.I0(pwm_counter[30]), .I1(n14_adj_4653), 
            .I2(n10_adj_4654), .I3(pwm_counter[24]), .O(n15453));
    defparam i7_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i12915_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n29542), 
            .I3(GND_net), .O(n17024));   // verilog/coms.v(127[12] 300[6])
    defparam i12915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12916_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n29542), 
            .I3(GND_net), .O(n17025));   // verilog/coms.v(127[12] 300[6])
    defparam i12916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12917_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n29542), 
            .I3(GND_net), .O(n17026));   // verilog/coms.v(127[12] 300[6])
    defparam i12917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12918_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n29542), 
            .I3(GND_net), .O(n17027));   // verilog/coms.v(127[12] 300[6])
    defparam i12918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4549));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12919_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n29542), 
            .I3(GND_net), .O(n17028));   // verilog/coms.v(127[12] 300[6])
    defparam i12919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4548));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4547));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_41_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[14]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12920_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n29542), 
            .I3(GND_net), .O(n17029));   // verilog/coms.v(127[12] 300[6])
    defparam i12920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12921_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n29542), 
            .I3(GND_net), .O(n17030));   // verilog/coms.v(127[12] 300[6])
    defparam i12921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4546));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1322_3_lut (.I0(n1934), .I1(n1987), 
            .I2(n1948), .I3(GND_net), .O(n2012));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1315_3_lut (.I0(n1927), .I1(n1980), 
            .I2(n1948), .I3(GND_net), .O(n2005));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12922_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n29542), 
            .I3(GND_net), .O(n17031));   // verilog/coms.v(127[12] 300[6])
    defparam i12922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4545));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1327_3_lut (.I0(n1939), .I1(n1992), 
            .I2(n1948), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1324_3_lut (.I0(n1936), .I1(n1989), 
            .I2(n1948), .I3(GND_net), .O(n2014));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1325_3_lut (.I0(n1937), .I1(n1990), 
            .I2(n1948), .I3(GND_net), .O(n2015));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1313_3_lut (.I0(n1925), .I1(n1978), 
            .I2(n1948), .I3(GND_net), .O(n2003));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1332_3_lut (.I0(n444), .I1(n1997), 
            .I2(n1948), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1331_3_lut (.I0(n1943), .I1(n1996), 
            .I2(n1948), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4503), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n445));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1317_3_lut (.I0(n1929), .I1(n1982), 
            .I2(n1948), .I3(GND_net), .O(n2007));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1323_3_lut (.I0(n1935), .I1(n1988), 
            .I2(n1948), .I3(GND_net), .O(n2013));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1314_3_lut (.I0(n1926), .I1(n1979), 
            .I2(n1948), .I3(GND_net), .O(n2004));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4532));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1319_3_lut (.I0(n1931), .I1(n1984), 
            .I2(n1948), .I3(GND_net), .O(n2009));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1316_3_lut (.I0(n1928), .I1(n1981), 
            .I2(n1948), .I3(GND_net), .O(n2006));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1320_3_lut (.I0(n1932), .I1(n1985), 
            .I2(n1948), .I3(GND_net), .O(n2010));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12798_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n29532), .I3(GND_net), .O(n16907));   // verilog/coms.v(127[12] 300[6])
    defparam i12798_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12799_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n29532), .I3(GND_net), .O(n16908));   // verilog/coms.v(127[12] 300[6])
    defparam i12799_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1326_3_lut (.I0(n1938), .I1(n1991), 
            .I2(n1948), .I3(GND_net), .O(n2016));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4544));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1310_3_lut (.I0(n1922), .I1(n1975), 
            .I2(n1948), .I3(GND_net), .O(n2000));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1330_3_lut (.I0(n1942), .I1(n1995), 
            .I2(n1948), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1328_3_lut (.I0(n1940), .I1(n1993), 
            .I2(n1948), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12800_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n29532), .I3(GND_net), .O(n16909));   // verilog/coms.v(127[12] 300[6])
    defparam i12800_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1329_3_lut (.I0(n1941), .I1(n1994), 
            .I2(n1948), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1311_3_lut (.I0(n1923), .I1(n1976), 
            .I2(n1948), .I3(GND_net), .O(n2001));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1318_3_lut (.I0(n1930), .I1(n1983), 
            .I2(n1948), .I3(GND_net), .O(n2008));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1321_3_lut (.I0(n1933), .I1(n1986), 
            .I2(n1948), .I3(GND_net), .O(n2011));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1312_3_lut (.I0(n1924), .I1(n1977), 
            .I2(n1948), .I3(GND_net), .O(n2002));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut (.I0(n2002), .I1(n2011), .I2(n2008), .I3(n2001), 
            .O(n30_adj_4565));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17887_3_lut (.I0(n445), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n21989));
    defparam i17887_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1621 (.I0(n2019), .I1(n2018), .I2(n21989), .I3(n2020), 
            .O(n30717));
    defparam i2_4_lut_adj_1621.LUT_INIT = 16'h8880;
    SB_LUT4 i15_4_lut (.I0(n2003), .I1(n30_adj_4565), .I2(n2015), .I3(n2014), 
            .O(n34_adj_4563));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2000), .I1(n2016), .I2(n2010), .I3(n2006), 
            .O(n32));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2009), .I1(n2004), .I2(n2013), .I3(n2007), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2017), .I1(n2005), .I2(n2012), .I3(n30717), 
            .O(n31_adj_4564));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(144[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12801_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n29532), .I3(GND_net), .O(n16910));   // verilog/coms.v(127[12] 300[6])
    defparam i12801_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1622 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n78), .I3(GND_net), .O(n63));
    defparam i2_3_lut_adj_1622.LUT_INIT = 16'hfdfd;
    SB_LUT4 i28748_4_lut (.I0(n31_adj_4564), .I1(n33), .I2(n32), .I3(n34_adj_4563), 
            .O(n2026));
    defparam i28748_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1494_3_lut (.I0(n2026), .I1(n4679), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[1]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1494_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1274_3_lut (.I0(n1861), .I1(n1914), 
            .I2(n1870), .I3(GND_net), .O(n1939));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1269_3_lut (.I0(n1856), .I1(n1909), 
            .I2(n1870), .I3(GND_net), .O(n1934));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12802_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n29532), .I3(GND_net), .O(n16911));   // verilog/coms.v(127[12] 300[6])
    defparam i12802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1275_3_lut (.I0(n1862), .I1(n1915), 
            .I2(n1870), .I3(GND_net), .O(n1940));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1278_3_lut (.I0(n443), .I1(n1918), 
            .I2(n1870), .I3(GND_net), .O(n1943));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1277_3_lut (.I0(n1864), .I1(n1917), 
            .I2(n1870), .I3(GND_net), .O(n1942));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1276_3_lut (.I0(n1863), .I1(n1916), 
            .I2(n1870), .I3(GND_net), .O(n1941));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4506), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n444));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_513_7_lut (.I0(GND_net), .I1(n754), 
            .I2(GND_net), .I3(n25149), .O(n807)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_7 (.CI(n25149), .I0(n754), 
            .I1(GND_net), .CO(n25150));
    SB_LUT4 encoder0_position_23__I_0_i1259_3_lut (.I0(n1846), .I1(n1899), 
            .I2(n1870), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_6_lut (.I0(GND_net), .I1(n755), 
            .I2(GND_net), .I3(n25148), .O(n808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1264_3_lut (.I0(n1851), .I1(n1904), 
            .I2(n1870), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1268_3_lut (.I0(n1855), .I1(n1908), 
            .I2(n1870), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1261_3_lut (.I0(n1848), .I1(n1901), 
            .I2(n1870), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1258_3_lut (.I0(n1845), .I1(n1898), 
            .I2(n1870), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_513_6 (.CI(n25148), .I0(n755), 
            .I1(GND_net), .CO(n25149));
    SB_LUT4 encoder0_position_23__I_0_i1262_3_lut (.I0(n1849), .I1(n1902), 
            .I2(n1870), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1267_3_lut (.I0(n1854), .I1(n1907), 
            .I2(n1870), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1272_3_lut (.I0(n1859), .I1(n1912), 
            .I2(n1870), .I3(GND_net), .O(n1937));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1273_3_lut (.I0(n1860), .I1(n1913), 
            .I2(n1870), .I3(GND_net), .O(n1938));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1273_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n25067), .I0(encoder1_position[14]), 
            .I1(n11_adj_4541), .CO(n25068));
    SB_LUT4 encoder0_position_23__I_0_i1260_3_lut (.I0(n1847), .I1(n1900), 
            .I2(n1870), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1271_3_lut (.I0(n1858), .I1(n1911), 
            .I2(n1870), .I3(GND_net), .O(n1936));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1257_3_lut (.I0(n1844), .I1(n1897), 
            .I2(n1870), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1265_3_lut (.I0(n1852), .I1(n1905), 
            .I2(n1870), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_5_lut (.I0(GND_net), .I1(n756), 
            .I2(VCC_net), .I3(n25147), .O(n809)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1266_3_lut (.I0(n1853), .I1(n1906), 
            .I2(n1870), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_513_5 (.CI(n25147), .I0(n756), 
            .I1(VCC_net), .CO(n25148));
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4542), .I3(n25066), .O(displacement_23__N_50[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1270_3_lut (.I0(n1857), .I1(n1910), 
            .I2(n1870), .I3(GND_net), .O(n1935));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1263_3_lut (.I0(n1850), .I1(n1903), 
            .I2(n1870), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_4_lut_adj_1623 (.I0(n1925), .I1(n1938), .I2(n1937), .I3(n1932), 
            .O(n28));
    defparam i10_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1624 (.I0(n1926), .I1(n1933), .I2(n1929), .I3(n1924), 
            .O(n31));
    defparam i13_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i17973_4_lut (.I0(n444), .I1(n1941), .I2(n1942), .I3(n1943), 
            .O(n22075));
    defparam i17973_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_2_lut (.I0(n1928), .I1(n1935), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4561));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1625 (.I0(n1931), .I1(n1930), .I2(n1922), .I3(n1936), 
            .O(n30));
    defparam i12_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1626 (.I0(n31), .I1(n1927), .I2(n28), .I3(n1923), 
            .O(n34));
    defparam i16_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i28381_1_lut (.I0(n700), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34057));
    defparam i28381_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_1627 (.I0(n1940), .I1(n1934), .I2(n1939), .I3(n22075), 
            .O(n21_adj_4562));
    defparam i3_4_lut_adj_1627.LUT_INIT = 16'heccc;
    SB_LUT4 i28723_4_lut (.I0(n21_adj_4562), .I1(n34), .I2(n30), .I3(n22_adj_4561), 
            .O(n1948));
    defparam i28723_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1493_3_lut (.I0(n1948), .I1(n4678), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[2]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1493_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1217_3_lut (.I0(n1779), .I1(n1832), 
            .I2(n1792), .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1215_3_lut (.I0(n1777), .I1(n1830), 
            .I2(n1792), .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1218_3_lut (.I0(n1780), .I1(n1833), 
            .I2(n1792), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1214_3_lut (.I0(n1776), .I1(n1829), 
            .I2(n1792), .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1207_3_lut (.I0(n1769), .I1(n1822), 
            .I2(n1792), .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1219_3_lut (.I0(n1781), .I1(n1834), 
            .I2(n1792), .I3(GND_net), .O(n1859));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1204_3_lut (.I0(n1766), .I1(n1819), 
            .I2(n1792), .I3(GND_net), .O(n1844));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1224_3_lut (.I0(n442), .I1(n1839), 
            .I2(n1792), .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1224_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1223_3_lut (.I0(n1785), .I1(n1838), 
            .I2(n1792), .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4507), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n443));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1208_3_lut (.I0(n1770), .I1(n1823), 
            .I2(n1792), .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1211_3_lut (.I0(n1773), .I1(n1826), 
            .I2(n1792), .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1213_3_lut (.I0(n1775), .I1(n1828), 
            .I2(n1792), .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1206_3_lut (.I0(n1768), .I1(n1821), 
            .I2(n1792), .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1209_3_lut (.I0(n1771), .I1(n1824), 
            .I2(n1792), .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1216_3_lut (.I0(n1778), .I1(n1831), 
            .I2(n1792), .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1210_3_lut (.I0(n1772), .I1(n1825), 
            .I2(n1792), .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1205_3_lut (.I0(n1767), .I1(n1820), 
            .I2(n1792), .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1212_3_lut (.I0(n1774), .I1(n1827), 
            .I2(n1792), .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_4_lut (.I0(GND_net), .I1(n757), 
            .I2(GND_net), .I3(n25146), .O(n810)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n25066), .I0(encoder1_position[13]), 
            .I1(n12_adj_4542), .CO(n25067));
    SB_LUT4 encoder0_position_23__I_0_i1222_3_lut (.I0(n1784), .I1(n1837), 
            .I2(n1792), .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1220_3_lut (.I0(n1782), .I1(n1835), 
            .I2(n1792), .I3(GND_net), .O(n1860));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1221_3_lut (.I0(n1783), .I1(n1836), 
            .I2(n1792), .I3(GND_net), .O(n1861));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1628 (.I0(n1851), .I1(n1848), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4634));
    defparam i1_2_lut_adj_1628.LUT_INIT = 16'heeee;
    SB_LUT4 i17899_3_lut (.I0(n443), .I1(n1863), .I2(n1864), .I3(GND_net), 
            .O(n22001));
    defparam i17899_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1629 (.I0(n1861), .I1(n1860), .I2(n22001), .I3(n1862), 
            .O(n31108));
    defparam i2_4_lut_adj_1629.LUT_INIT = 16'h8880;
    SB_LUT4 i13_4_lut_adj_1630 (.I0(n1844), .I1(n1859), .I2(n1847), .I3(n18_adj_4634), 
            .O(n30_adj_4630));
    defparam i13_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1631 (.I0(n1852), .I1(n31108), .I2(n1845), .I3(n1850), 
            .O(n28_adj_4632));
    defparam i11_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1632 (.I0(n1856), .I1(n1849), .I2(n1846), .I3(n1853), 
            .O(n29_adj_4631));
    defparam i12_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1633 (.I0(n1854), .I1(n1858), .I2(n1855), .I3(n1857), 
            .O(n27_adj_4633));
    defparam i10_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i28696_4_lut (.I0(n27_adj_4633), .I1(n29_adj_4631), .I2(n28_adj_4632), 
            .I3(n30_adj_4630), .O(n1870));
    defparam i28696_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1492_3_lut (.I0(n1870), .I1(n4677), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[3]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1492_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1165_3_lut (.I0(n1702), .I1(n1755), 
            .I2(n1714), .I3(GND_net), .O(n1780));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1165_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1154_3_lut (.I0(n1691), .I1(n1744), 
            .I2(n1714), .I3(GND_net), .O(n1769));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1161_3_lut (.I0(n1698), .I1(n1751), 
            .I2(n1714), .I3(GND_net), .O(n1776));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4543));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1164_3_lut (.I0(n1701), .I1(n1754), 
            .I2(n1714), .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1160_3_lut (.I0(n1697), .I1(n1750), 
            .I2(n1714), .I3(GND_net), .O(n1775));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1160_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4542));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1152_3_lut (.I0(n1689), .I1(n1742), 
            .I2(n1714), .I3(GND_net), .O(n1767));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1157_3_lut (.I0(n1694), .I1(n1747), 
            .I2(n1714), .I3(GND_net), .O(n1772));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1168_3_lut (.I0(n1705), .I1(n1758), 
            .I2(n1714), .I3(GND_net), .O(n1783));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1166_3_lut (.I0(n1703), .I1(n1756), 
            .I2(n1714), .I3(GND_net), .O(n1781));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1167_3_lut (.I0(n1704), .I1(n1757), 
            .I2(n1714), .I3(GND_net), .O(n1782));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1170_3_lut (.I0(n441), .I1(n1760), 
            .I2(n1714), .I3(GND_net), .O(n1785));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1169_3_lut (.I0(n1706), .I1(n1759), 
            .I2(n1714), .I3(GND_net), .O(n1784));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4508), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n442));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1153_3_lut (.I0(n1690), .I1(n1743), 
            .I2(n1714), .I3(GND_net), .O(n1768));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1159_3_lut (.I0(n1696), .I1(n1749), 
            .I2(n1714), .I3(GND_net), .O(n1774));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1162_3_lut (.I0(n1699), .I1(n1752), 
            .I2(n1714), .I3(GND_net), .O(n1777));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1162_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1163_3_lut (.I0(n1700), .I1(n1753), 
            .I2(n1714), .I3(GND_net), .O(n1778));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1163_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1156_3_lut (.I0(n1693), .I1(n1746), 
            .I2(n1714), .I3(GND_net), .O(n1771));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1151_3_lut (.I0(n1688), .I1(n1741), 
            .I2(n1714), .I3(GND_net), .O(n1766));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1158_3_lut (.I0(n1695), .I1(n1748), 
            .I2(n1714), .I3(GND_net), .O(n1773));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12743_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n28583), .I3(GND_net), .O(n16852));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12743_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1155_3_lut (.I0(n1692), .I1(n1745), 
            .I2(n1714), .I3(GND_net), .O(n1770));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17901_3_lut (.I0(n442), .I1(n1784), .I2(n1785), .I3(GND_net), 
            .O(n22003));
    defparam i17901_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i12744_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n4216), .I3(GND_net), .O(n16853));   // verilog/coms.v(127[12] 300[6])
    defparam i12744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1634 (.I0(n1782), .I1(n1781), .I2(n22003), .I3(n1783), 
            .O(n30832));
    defparam i2_4_lut_adj_1634.LUT_INIT = 16'h8880;
    SB_LUT4 i12_4_lut_adj_1635 (.I0(n1772), .I1(n1767), .I2(n1775), .I3(n1779), 
            .O(n28_adj_4626));
    defparam i12_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1636 (.I0(n1770), .I1(n1773), .I2(n1766), .I3(n1771), 
            .O(n26_adj_4628));
    defparam i10_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1637 (.I0(n1778), .I1(n1777), .I2(n1774), .I3(n1768), 
            .O(n27_adj_4627));
    defparam i11_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1638 (.I0(n30832), .I1(n1776), .I2(n1769), .I3(n1780), 
            .O(n25_adj_4629));
    defparam i9_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 i28670_4_lut (.I0(n25_adj_4629), .I1(n27_adj_4627), .I2(n26_adj_4628), 
            .I3(n28_adj_4626), .O(n1792));
    defparam i28670_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1491_3_lut (.I0(n1792), .I1(n4676), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[4]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1491_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i12746_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n21215), 
            .I3(n15595), .O(n16855));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12746_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_23__I_0_i1103_3_lut (.I0(n1615), .I1(n1668), 
            .I2(n1636), .I3(GND_net), .O(n1693));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1108_3_lut (.I0(n1620), .I1(n1673), 
            .I2(n1636), .I3(GND_net), .O(n1698));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1102_3_lut (.I0(n1614), .I1(n1667), 
            .I2(n1636), .I3(GND_net), .O(n1692));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12747_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n21215), 
            .I3(n15590), .O(n16856));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12747_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12748_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n15595), 
            .O(n16857));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12748_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i1105_3_lut (.I0(n1617), .I1(n1670), 
            .I2(n1636), .I3(GND_net), .O(n1695));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1110_3_lut (.I0(n1622), .I1(n1675), 
            .I2(n1636), .I3(GND_net), .O(n1700));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1101_3_lut (.I0(n1613), .I1(n1666), 
            .I2(n1636), .I3(GND_net), .O(n1691));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1114_3_lut (.I0(n1626), .I1(n1679), 
            .I2(n1636), .I3(GND_net), .O(n1704));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1112_3_lut (.I0(n1624), .I1(n1677), 
            .I2(n1636), .I3(GND_net), .O(n1702));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1113_3_lut (.I0(n1625), .I1(n1678), 
            .I2(n1636), .I3(GND_net), .O(n1703));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1104_3_lut (.I0(n1616), .I1(n1669), 
            .I2(n1636), .I3(GND_net), .O(n1694));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4543), .I3(n25065), .O(displacement_23__N_50[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12749_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n15590), 
            .O(n16858));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12749_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i1109_3_lut (.I0(n1621), .I1(n1674), 
            .I2(n1636), .I3(GND_net), .O(n1699));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1107_3_lut (.I0(n1619), .I1(n1672), 
            .I2(n1636), .I3(GND_net), .O(n1697));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1111_3_lut (.I0(n1623), .I1(n1676), 
            .I2(n1636), .I3(GND_net), .O(n1701));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1098_3_lut (.I0(n1610), .I1(n1663), 
            .I2(n1636), .I3(GND_net), .O(n1688));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28518_1_lut (.I0(n778), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34194));
    defparam i28518_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1106_3_lut (.I0(n1618), .I1(n1671), 
            .I2(n1636), .I3(GND_net), .O(n1696));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1099_3_lut (.I0(n1611), .I1(n1664), 
            .I2(n1636), .I3(GND_net), .O(n1689));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1099_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4520), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n430));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1100_3_lut (.I0(n1612), .I1(n1665), 
            .I2(n1636), .I3(GND_net), .O(n1690));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1116_3_lut (.I0(n440), .I1(n1681), 
            .I2(n1636), .I3(GND_net), .O(n1706));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i522_3_lut (.I0(n429), .I1(n812), 
            .I2(n778), .I3(GND_net), .O(n837));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1115_3_lut (.I0(n1627), .I1(n1680), 
            .I2(n1636), .I3(GND_net), .O(n1705));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4509), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n441));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17905_3_lut (.I0(n441), .I1(n1705), .I2(n1706), .I3(GND_net), 
            .O(n22007));
    defparam i17905_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1639 (.I0(n1703), .I1(n1702), .I2(n22007), .I3(n1704), 
            .O(n30808));
    defparam i2_4_lut_adj_1639.LUT_INIT = 16'h8880;
    SB_LUT4 i11_4_lut_adj_1640 (.I0(n1690), .I1(n1689), .I2(n1696), .I3(n1688), 
            .O(n26_adj_4586));
    defparam i11_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1641 (.I0(n1691), .I1(n30808), .I2(n1700), .I3(n1695), 
            .O(n24_adj_4588));
    defparam i9_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i521_3_lut (.I0(n758), .I1(n811), 
            .I2(n778), .I3(GND_net), .O(n836));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_4_lut_adj_1642 (.I0(n1701), .I1(n1697), .I2(n1699), .I3(n1694), 
            .O(n25_adj_4587));
    defparam i10_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut (.I0(n1692), .I1(n1698), .I2(n1693), .I3(GND_net), 
            .O(n23_adj_4589));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_23__I_0_add_513_4 (.CI(n25146), .I0(n757), 
            .I1(GND_net), .CO(n25147));
    SB_LUT4 i28642_4_lut (.I0(n23_adj_4589), .I1(n25_adj_4587), .I2(n24_adj_4588), 
            .I3(n26_adj_4586), .O(n1714));
    defparam i28642_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1490_3_lut (.I0(n1714), .I1(n4675), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[5]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1490_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_add_513_3_lut (.I0(GND_net), .I1(n758), 
            .I2(VCC_net), .I3(n25145), .O(n811)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4541));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1054_3_lut (.I0(n1541), .I1(n1594), 
            .I2(n1558), .I3(GND_net), .O(n1619));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1056_3_lut (.I0(n1543), .I1(n1596), 
            .I2(n1558), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1055_3_lut (.I0(n1542), .I1(n1595), 
            .I2(n1558), .I3(GND_net), .O(n1620));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1057_3_lut (.I0(n1544), .I1(n1597), 
            .I2(n1558), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1045_3_lut (.I0(n1532), .I1(n1585), 
            .I2(n1558), .I3(GND_net), .O(n1610));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1050_3_lut (.I0(n1537), .I1(n1590), 
            .I2(n1558), .I3(GND_net), .O(n1615));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1052_3_lut (.I0(n1539), .I1(n1592), 
            .I2(n1558), .I3(GND_net), .O(n1617));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1047_3_lut (.I0(n1534), .I1(n1587), 
            .I2(n1558), .I3(GND_net), .O(n1612));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12750_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4535), 
            .I3(n15595), .O(n16859));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12750_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i1049_3_lut (.I0(n1536), .I1(n1589), 
            .I2(n1558), .I3(GND_net), .O(n1614));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_513_3 (.CI(n25145), .I0(n758), 
            .I1(VCC_net), .CO(n25146));
    SB_LUT4 i12751_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4535), 
            .I3(n15590), .O(n16860));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12751_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12752_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4530), 
            .I3(n15595), .O(n16861));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12752_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i1060_3_lut (.I0(n1547), .I1(n1600), 
            .I2(n1558), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1058_3_lut (.I0(n1545), .I1(n1598), 
            .I2(n1558), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1059_3_lut (.I0(n1546), .I1(n1599), 
            .I2(n1558), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12753_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n16862));   // verilog/coms.v(127[12] 300[6])
    defparam i12753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1048_3_lut (.I0(n1535), .I1(n1588), 
            .I2(n1558), .I3(GND_net), .O(n1613));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12754_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n8868), 
            .I3(GND_net), .O(n16863));   // verilog/coms.v(127[12] 300[6])
    defparam i12754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1051_3_lut (.I0(n1538), .I1(n1591), 
            .I2(n1558), .I3(GND_net), .O(n1616));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1053_3_lut (.I0(n1540), .I1(n1593), 
            .I2(n1558), .I3(GND_net), .O(n1618));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12755_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n8868), 
            .I3(GND_net), .O(n16864));   // verilog/coms.v(127[12] 300[6])
    defparam i12755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_513_2_lut (.I0(GND_net), .I1(n429), 
            .I2(GND_net), .I3(VCC_net), .O(n812)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1046_3_lut (.I0(n1533), .I1(n1586), 
            .I2(n1558), .I3(GND_net), .O(n1611));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1062_3_lut (.I0(n439), .I1(n1602), 
            .I2(n1558), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12756_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n4218), .I3(GND_net), .O(n16865));   // verilog/coms.v(127[12] 300[6])
    defparam i12756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1061_3_lut (.I0(n1548), .I1(n1601), 
            .I2(n1558), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12970_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n4218), .I3(GND_net), .O(n17079));   // verilog/coms.v(127[12] 300[6])
    defparam i12970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2782_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4510), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n440));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17907_3_lut (.I0(n440), .I1(n1626), .I2(n1627), .I3(GND_net), 
            .O(n22009));
    defparam i17907_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1643 (.I0(n1624), .I1(n1623), .I2(n22009), .I3(n1625), 
            .O(n31395));
    defparam i2_4_lut_adj_1643.LUT_INIT = 16'h8880;
    SB_LUT4 i12971_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n4218), .I3(GND_net), .O(n17080));   // verilog/coms.v(127[12] 300[6])
    defparam i12971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_2_lut_adj_1644 (.I0(n1611), .I1(n1618), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4501));
    defparam i4_2_lut_adj_1644.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1645 (.I0(n1614), .I1(n1612), .I2(n1617), .I3(n1615), 
            .O(n24_adj_4499));
    defparam i10_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1646 (.I0(n1610), .I1(n1622), .I2(n1620), .I3(n31395), 
            .O(n22_adj_4500));
    defparam i8_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i12972_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n4218), .I3(GND_net), .O(n17081));   // verilog/coms.v(127[12] 300[6])
    defparam i12972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1647 (.I0(n1616), .I1(n24_adj_4499), .I2(n18_adj_4501), 
            .I3(n1613), .O(n26));
    defparam i12_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 i12973_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n4218), .I3(GND_net), .O(n17082));   // verilog/coms.v(127[12] 300[6])
    defparam i12973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28618_4_lut (.I0(n1621), .I1(n26), .I2(n22_adj_4500), .I3(n1619), 
            .O(n1636));
    defparam i28618_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1489_3_lut (.I0(n1636), .I1(n4674), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[6]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1489_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i12974_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n4218), .I3(GND_net), .O(n17083));   // verilog/coms.v(127[12] 300[6])
    defparam i12974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1001_3_lut (.I0(n1463), .I1(n1516), 
            .I2(n1480), .I3(GND_net), .O(n1541));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i995_3_lut (.I0(n1457), .I1(n1510), 
            .I2(n1480), .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12975_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n4218), .I3(GND_net), .O(n17084));   // verilog/coms.v(127[12] 300[6])
    defparam i12975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12976_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n4218), .I3(GND_net), .O(n17085));   // verilog/coms.v(127[12] 300[6])
    defparam i12976_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n25065), .I0(encoder1_position[12]), 
            .I1(n13_adj_4543), .CO(n25066));
    SB_LUT4 i12977_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n4218), .I3(GND_net), .O(n17086));   // verilog/coms.v(127[12] 300[6])
    defparam i12977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i992_3_lut (.I0(n1454), .I1(n1507), 
            .I2(n1480), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12978_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n4218), .I3(GND_net), .O(n17087));   // verilog/coms.v(127[12] 300[6])
    defparam i12978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i997_3_lut (.I0(n1459), .I1(n1512), 
            .I2(n1480), .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1004_3_lut (.I0(n1466), .I1(n1519), 
            .I2(n1480), .I3(GND_net), .O(n1544));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12979_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n4218), .I3(GND_net), .O(n17088));   // verilog/coms.v(127[12] 300[6])
    defparam i12979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i994_3_lut (.I0(n1456), .I1(n1509), 
            .I2(n1480), .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12980_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n4218), .I3(GND_net), .O(n17089));   // verilog/coms.v(127[12] 300[6])
    defparam i12980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12981_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n4218), .I3(GND_net), .O(n17090));   // verilog/coms.v(127[12] 300[6])
    defparam i12981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1005_3_lut (.I0(n1467), .I1(n1520), 
            .I2(n1480), .I3(GND_net), .O(n1545));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1003_3_lut (.I0(n1465), .I1(n1518), 
            .I2(n1480), .I3(GND_net), .O(n1543));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12982_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n4218), .I3(GND_net), .O(n17091));   // verilog/coms.v(127[12] 300[6])
    defparam i12982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12983_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n4218), .I3(GND_net), .O(n17092));   // verilog/coms.v(127[12] 300[6])
    defparam i12983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i996_3_lut (.I0(n1458), .I1(n1511), 
            .I2(n1480), .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i999_3_lut (.I0(n1461), .I1(n1514), 
            .I2(n1480), .I3(GND_net), .O(n1539));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1000_3_lut (.I0(n1462), .I1(n1515), 
            .I2(n1480), .I3(GND_net), .O(n1540));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i998_3_lut (.I0(n1460), .I1(n1513), 
            .I2(n1480), .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12984_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n4218), .I3(GND_net), .O(n17093));   // verilog/coms.v(127[12] 300[6])
    defparam i12984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1002_3_lut (.I0(n1464), .I1(n1517), 
            .I2(n1480), .I3(GND_net), .O(n1542));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i993_3_lut (.I0(n1455), .I1(n1508), 
            .I2(n1480), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12985_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n4218), .I3(GND_net), .O(n17094));   // verilog/coms.v(127[12] 300[6])
    defparam i12985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1008_3_lut (.I0(n438), .I1(n1523), 
            .I2(n1480), .I3(GND_net), .O(n1548));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1007_3_lut (.I0(n1469), .I1(n1522), 
            .I2(n1480), .I3(GND_net), .O(n1547));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1006_3_lut (.I0(n1468), .I1(n1521), 
            .I2(n1480), .I3(GND_net), .O(n1546));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1006_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12986_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n4218), .I3(GND_net), .O(n17095));   // verilog/coms.v(127[12] 300[6])
    defparam i12986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2782_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_4511), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n439));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4544), .I3(n25064), .O(displacement_23__N_50[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17993_4_lut (.I0(n439), .I1(n1546), .I2(n1547), .I3(n1548), 
            .O(n22095));
    defparam i17993_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut_adj_1648 (.I0(n1545), .I1(n1534), .I2(n1544), .I3(n22095), 
            .O(n17_adj_4493));
    defparam i4_4_lut_adj_1648.LUT_INIT = 16'heccc;
    SB_LUT4 i8_4_lut_adj_1649 (.I0(n1533), .I1(n1542), .I2(n1538), .I3(n1540), 
            .O(n21_adj_4491));
    defparam i8_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1539), .I1(n1536), .I2(n1543), .I3(GND_net), 
            .O(n20_adj_4492));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12987_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n4218), .I3(GND_net), .O(n17096));   // verilog/coms.v(127[12] 300[6])
    defparam i12987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1650 (.I0(n21_adj_4491), .I1(n17_adj_4493), .I2(n1537), 
            .I3(n1532), .O(n24_adj_4490));
    defparam i11_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i12988_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n4218), .I3(GND_net), .O(n17097));   // verilog/coms.v(127[12] 300[6])
    defparam i12988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12989_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n4218), .I3(GND_net), .O(n17098));   // verilog/coms.v(127[12] 300[6])
    defparam i12989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28595_4_lut (.I0(n1535), .I1(n24_adj_4490), .I2(n20_adj_4492), 
            .I3(n1541), .O(n1558));
    defparam i28595_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i12990_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n4218), .I3(GND_net), .O(n17099));   // verilog/coms.v(127[12] 300[6])
    defparam i12990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1488_3_lut (.I0(n1558), .I1(n4673), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[7]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1488_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i943_3_lut (.I0(n1380), .I1(n1433), 
            .I2(n1402), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12991_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n4218), .I3(GND_net), .O(n17100));   // verilog/coms.v(127[12] 300[6])
    defparam i12991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i944_3_lut (.I0(n1381), .I1(n1434), 
            .I2(n1402), .I3(GND_net), .O(n1459));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i946_3_lut (.I0(n1383), .I1(n1436), 
            .I2(n1402), .I3(GND_net), .O(n1461));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i942_3_lut (.I0(n1379), .I1(n1432), 
            .I2(n1402), .I3(GND_net), .O(n1457));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i941_3_lut (.I0(n1378), .I1(n1431), 
            .I2(n1402), .I3(GND_net), .O(n1456));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12992_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n4218), .I3(GND_net), .O(n17101));   // verilog/coms.v(127[12] 300[6])
    defparam i12992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i939_3_lut (.I0(n1376), .I1(n1429), 
            .I2(n1402), .I3(GND_net), .O(n1454));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i954_3_lut (.I0(n437), .I1(n1444), 
            .I2(n1402), .I3(GND_net), .O(n1469));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12993_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n12944), .I3(GND_net), .O(n17102));   // verilog/coms.v(127[12] 300[6])
    defparam i12993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12994_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n12944), .I3(GND_net), .O(n17103));   // verilog/coms.v(127[12] 300[6])
    defparam i12994_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n25064), .I0(encoder1_position[11]), 
            .I1(n14_adj_4544), .CO(n25065));
    SB_LUT4 encoder0_position_23__I_0_i953_3_lut (.I0(n1390), .I1(n1443), 
            .I2(n1402), .I3(GND_net), .O(n1468));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i952_3_lut (.I0(n1389), .I1(n1442), 
            .I2(n1402), .I3(GND_net), .O(n1467));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12995_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n12944), .I3(GND_net), .O(n17104));   // verilog/coms.v(127[12] 300[6])
    defparam i12995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12996_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n12944), .I3(GND_net), .O(n17105));   // verilog/coms.v(127[12] 300[6])
    defparam i12996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2782_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4512), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n438));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i940_3_lut (.I0(n1377), .I1(n1430), 
            .I2(n1402), .I3(GND_net), .O(n1455));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12997_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n12944), .I3(GND_net), .O(n17106));   // verilog/coms.v(127[12] 300[6])
    defparam i12997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i949_3_lut (.I0(n1386), .I1(n1439), 
            .I2(n1402), .I3(GND_net), .O(n1464));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i947_3_lut (.I0(n1384), .I1(n1437), 
            .I2(n1402), .I3(GND_net), .O(n1462));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i945_3_lut (.I0(n1382), .I1(n1435), 
            .I2(n1402), .I3(GND_net), .O(n1460));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i950_3_lut (.I0(n1387), .I1(n1440), 
            .I2(n1402), .I3(GND_net), .O(n1465));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i950_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12998_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n12944), .I3(GND_net), .O(n17107));   // verilog/coms.v(127[12] 300[6])
    defparam i12998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i948_3_lut (.I0(n1385), .I1(n1438), 
            .I2(n1402), .I3(GND_net), .O(n1463));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i948_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i951_3_lut (.I0(n1388), .I1(n1441), 
            .I2(n1402), .I3(GND_net), .O(n1466));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i951_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4545), .I3(n25063), .O(displacement_23__N_50[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17995_4_lut (.I0(n438), .I1(n1467), .I2(n1468), .I3(n1469), 
            .O(n22097));
    defparam i17995_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n1466), .I1(n1463), .I2(n1465), .I3(n22097), 
            .O(n5_adj_4498));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'heccc;
    SB_LUT4 i2_2_lut_adj_1652 (.I0(n1454), .I1(n1456), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4559));
    defparam i2_2_lut_adj_1652.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(n1457), .I1(n5_adj_4498), .I2(n1461), 
            .I3(n1459), .O(n7_adj_4560));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_DFF h1_26 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n25063), .I0(encoder1_position[10]), 
            .I1(n15_adj_4545), .CO(n25064));
    SB_LUT4 i12999_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n12944), .I3(GND_net), .O(n17108));   // verilog/coms.v(127[12] 300[6])
    defparam i12999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1654 (.I0(n1460), .I1(n1462), .I2(n1464), .I3(n1455), 
            .O(n31908));
    defparam i3_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i28809_4_lut (.I0(n31908), .I1(n7_adj_4560), .I2(n1458), .I3(n8_adj_4559), 
            .O(n1480));
    defparam i28809_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1487_3_lut (.I0(n1480), .I1(n4672), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[8]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1487_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i892_3_lut (.I0(n1304), .I1(n1357), 
            .I2(n1324), .I3(GND_net), .O(n1382));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i886_3_lut (.I0(n1298), .I1(n1351), 
            .I2(n1324), .I3(GND_net), .O(n1376));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i891_3_lut (.I0(n1303), .I1(n1356), 
            .I2(n1324), .I3(GND_net), .O(n1381));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i895_3_lut (.I0(n1307), .I1(n1360), 
            .I2(n1324), .I3(GND_net), .O(n1385));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i898_3_lut (.I0(n1310), .I1(n1363), 
            .I2(n1324), .I3(GND_net), .O(n1388));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i898_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i896_3_lut (.I0(n1308), .I1(n1361), 
            .I2(n1324), .I3(GND_net), .O(n1386));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i897_3_lut (.I0(n1309), .I1(n1362), 
            .I2(n1324), .I3(GND_net), .O(n1387));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i900_3_lut (.I0(n436), .I1(n1365), 
            .I2(n1324), .I3(GND_net), .O(n1390));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i899_3_lut (.I0(n1311), .I1(n1364), 
            .I2(n1324), .I3(GND_net), .O(n1389));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4513), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n437));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i888_3_lut (.I0(n1300), .I1(n1353), 
            .I2(n1324), .I3(GND_net), .O(n1378));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i894_3_lut (.I0(n1306), .I1(n1359), 
            .I2(n1324), .I3(GND_net), .O(n1384));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i894_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i889_3_lut (.I0(n1301), .I1(n1354), 
            .I2(n1324), .I3(GND_net), .O(n1379));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13000_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n12944), .I3(GND_net), .O(n17109));   // verilog/coms.v(127[12] 300[6])
    defparam i13000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i887_3_lut (.I0(n1299), .I1(n1352), 
            .I2(n1324), .I3(GND_net), .O(n1377));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i890_3_lut (.I0(n1302), .I1(n1355), 
            .I2(n1324), .I3(GND_net), .O(n1380));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i890_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i893_3_lut (.I0(n1305), .I1(n1358), 
            .I2(n1324), .I3(GND_net), .O(n1383));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17919_3_lut (.I0(n437), .I1(n1389), .I2(n1390), .I3(GND_net), 
            .O(n22021));
    defparam i17919_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1655 (.I0(n1387), .I1(n1386), .I2(n22021), .I3(n1388), 
            .O(n31590));
    defparam i2_4_lut_adj_1655.LUT_INIT = 16'h8880;
    SB_LUT4 i7_4_lut_adj_1656 (.I0(n1383), .I1(n1380), .I2(n1377), .I3(n31590), 
            .O(n18_adj_4557));
    defparam i7_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1385), .I1(n1381), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4558));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1657 (.I0(n1379), .I1(n18_adj_4557), .I2(n1384), 
            .I3(n1378), .O(n20_adj_4556));
    defparam i9_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 i28517_4_lut (.I0(n1376), .I1(n20_adj_4556), .I2(n16_adj_4558), 
            .I3(n1382), .O(n1402));
    defparam i28517_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1486_3_lut (.I0(n1402), .I1(n4671), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[9]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1486_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i834_3_lut (.I0(n1221), .I1(n1274), 
            .I2(n1246), .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i836_3_lut (.I0(n1223), .I1(n1276), 
            .I2(n1246), .I3(GND_net), .O(n1301));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i839_3_lut (.I0(n1226), .I1(n1279), 
            .I2(n1246), .I3(GND_net), .O(n1304));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i841_3_lut (.I0(n1228), .I1(n1281), 
            .I2(n1246), .I3(GND_net), .O(n1306));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i835_3_lut (.I0(n1222), .I1(n1275), 
            .I2(n1246), .I3(GND_net), .O(n1300));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i846_3_lut (.I0(n435), .I1(n1286), 
            .I2(n1246), .I3(GND_net), .O(n1311));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i845_3_lut (.I0(n1232), .I1(n1285), 
            .I2(n1246), .I3(GND_net), .O(n1310));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4514), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n436));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i840_3_lut (.I0(n1227), .I1(n1280), 
            .I2(n1246), .I3(GND_net), .O(n1305));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i833_3_lut (.I0(n1220), .I1(n1273), 
            .I2(n1246), .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i833_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i837_3_lut (.I0(n1224), .I1(n1277), 
            .I2(n1246), .I3(GND_net), .O(n1302));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i838_3_lut (.I0(n1225), .I1(n1278), 
            .I2(n1246), .I3(GND_net), .O(n1303));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i844_3_lut (.I0(n1231), .I1(n1284), 
            .I2(n1246), .I3(GND_net), .O(n1309));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i842_3_lut (.I0(n1229), .I1(n1282), 
            .I2(n1246), .I3(GND_net), .O(n1307));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i843_3_lut (.I0(n1230), .I1(n1283), 
            .I2(n1246), .I3(GND_net), .O(n1308));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4546), .I3(n25062), .O(displacement_23__N_50[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17921_3_lut (.I0(n436), .I1(n1310), .I2(n1311), .I3(GND_net), 
            .O(n22023));
    defparam i17921_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1658 (.I0(n1308), .I1(n1307), .I2(n22023), .I3(n1309), 
            .O(n31097));
    defparam i2_4_lut_adj_1658.LUT_INIT = 16'h8880;
    SB_LUT4 i6_4_lut_adj_1659 (.I0(n1300), .I1(n31097), .I2(n1306), .I3(n1304), 
            .O(n16_adj_4623));
    defparam i6_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n25062), .I0(encoder1_position[9]), 
            .I1(n16_adj_4546), .CO(n25063));
    SB_LUT4 i7_4_lut_adj_1660 (.I0(n1303), .I1(n1302), .I2(n1298), .I3(n1305), 
            .O(n17_adj_4622));
    defparam i7_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i28497_4_lut (.I0(n17_adj_4622), .I1(n1301), .I2(n16_adj_4623), 
            .I3(n1299), .O(n1324));
    defparam i28497_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1485_3_lut (.I0(n1324), .I1(n4670), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[10]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1485_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i780_3_lut (.I0(n1142), .I1(n1195), 
            .I2(n1168), .I3(GND_net), .O(n1220));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i786_3_lut (.I0(n1148), .I1(n1201), 
            .I2(n1168), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i788_3_lut (.I0(n1150), .I1(n1203), 
            .I2(n1168), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i782_3_lut (.I0(n1144), .I1(n1197), 
            .I2(n1168), .I3(GND_net), .O(n1222));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i789_3_lut (.I0(n1151), .I1(n1204), 
            .I2(n1168), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i781_3_lut (.I0(n1143), .I1(n1196), 
            .I2(n1168), .I3(GND_net), .O(n1221));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i787_3_lut (.I0(n1149), .I1(n1202), 
            .I2(n1168), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i785_3_lut (.I0(n1147), .I1(n1200), 
            .I2(n1168), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i784_3_lut (.I0(n1146), .I1(n1199), 
            .I2(n1168), .I3(GND_net), .O(n1224));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4547), .I3(n25061), .O(displacement_23__N_50[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i783_3_lut (.I0(n1145), .I1(n1198), 
            .I2(n1168), .I3(GND_net), .O(n1223));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i792_3_lut (.I0(n434), .I1(n1207), 
            .I2(n1168), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i791_3_lut (.I0(n1153), .I1(n1206), 
            .I2(n1168), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i790_3_lut (.I0(n1152), .I1(n1205), 
            .I2(n1168), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4515), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n435));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17933_4_lut (.I0(n435), .I1(n1230), .I2(n1231), .I3(n1232), 
            .O(n22035));
    defparam i17933_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1661 (.I0(n1223), .I1(n1224), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4637));
    defparam i1_2_lut_adj_1661.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1662 (.I0(n1229), .I1(n1222), .I2(n1228), .I3(n22035), 
            .O(n12_adj_4636));
    defparam i3_4_lut_adj_1662.LUT_INIT = 16'heccc;
    SB_CARRY encoder0_position_23__I_0_add_513_2 (.CI(VCC_net), .I0(n429), 
            .I1(GND_net), .CO(n25145));
    SB_LUT4 i7_4_lut_adj_1663 (.I0(n1225), .I1(n1227), .I2(n1221), .I3(n10_adj_4637), 
            .O(n16_adj_4635));
    defparam i7_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i28425_4_lut (.I0(n1226), .I1(n16_adj_4635), .I2(n12_adj_4636), 
            .I3(n1220), .O(n1246));
    defparam i28425_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1484_3_lut (.I0(n1246), .I1(n4669), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[11]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1484_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n25061), .I0(encoder1_position[8]), 
            .I1(n17_adj_4547), .CO(n25062));
    SB_LUT4 encoder0_position_23__I_0_i728_3_lut (.I0(n1065), .I1(n1118), 
            .I2(n1090), .I3(GND_net), .O(n1143));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i727_3_lut (.I0(n1064), .I1(n1117), 
            .I2(n1090), .I3(GND_net), .O(n1142));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i738_3_lut (.I0(n433), .I1(n1128), 
            .I2(n1090), .I3(GND_net), .O(n1153));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i737_3_lut (.I0(n1074), .I1(n1127), 
            .I2(n1090), .I3(GND_net), .O(n1152));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4548), .I3(n25060), .O(displacement_23__N_50[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i736_3_lut (.I0(n1073), .I1(n1126), 
            .I2(n1090), .I3(GND_net), .O(n1151));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i736_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n25060), .I0(encoder1_position[7]), 
            .I1(n18_adj_4548), .CO(n25061));
    SB_LUT4 mux_2782_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4516), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n434));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i734_3_lut (.I0(n1071), .I1(n1124), 
            .I2(n1090), .I3(GND_net), .O(n1149));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i730_3_lut (.I0(n1067), .I1(n1120), 
            .I2(n1090), .I3(GND_net), .O(n1145));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i730_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i735_3_lut (.I0(n1072), .I1(n1125), 
            .I2(n1090), .I3(GND_net), .O(n1150));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13001_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n12944), .I3(GND_net), .O(n17110));   // verilog/coms.v(127[12] 300[6])
    defparam i13001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i732_3_lut (.I0(n1069), .I1(n1122), 
            .I2(n1090), .I3(GND_net), .O(n1147));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i732_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i729_3_lut (.I0(n1066), .I1(n1119), 
            .I2(n1090), .I3(GND_net), .O(n1144));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1495_3_lut (.I0(n22055), .I1(n4680), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[0]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1495_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i733_3_lut (.I0(n1070), .I1(n1123), 
            .I2(n1090), .I3(GND_net), .O(n1148));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i733_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4549), .I3(n25059), .O(displacement_23__N_50[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i731_3_lut (.I0(n1068), .I1(n1121), 
            .I2(n1090), .I3(GND_net), .O(n1146));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17939_4_lut (.I0(n434), .I1(n1151), .I2(n1152), .I3(n1153), 
            .O(n22041));
    defparam i17939_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i6_4_lut_adj_1664 (.I0(n1146), .I1(n1148), .I2(n1144), .I3(n1147), 
            .O(n14_adj_4496));
    defparam i6_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[0]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 i1_4_lut_adj_1665 (.I0(n1150), .I1(n1145), .I2(n1149), .I3(n22041), 
            .O(n9_adj_4497));
    defparam i1_4_lut_adj_1665.LUT_INIT = 16'heccc;
    SB_LUT4 i28573_4_lut (.I0(n9_adj_4497), .I1(n14_adj_4496), .I2(n1142), 
            .I3(n1143), .O(n1168));
    defparam i28573_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1483_3_lut (.I0(n1168), .I1(n4668), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[12]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1483_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i679_3_lut (.I0(n991), .I1(n1044), 
            .I2(n1012), .I3(GND_net), .O(n1069));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i679_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i676_3_lut (.I0(n988), .I1(n1041), 
            .I2(n1012), .I3(GND_net), .O(n1066));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i677_3_lut (.I0(n989), .I1(n1042), 
            .I2(n1012), .I3(GND_net), .O(n1067));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i682_3_lut (.I0(n994), .I1(n1047), 
            .I2(n1012), .I3(GND_net), .O(n1072));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i682_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i680_3_lut (.I0(n992), .I1(n1045), 
            .I2(n1012), .I3(GND_net), .O(n1070));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i680_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i681_3_lut (.I0(n993), .I1(n1046), 
            .I2(n1012), .I3(GND_net), .O(n1071));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i678_3_lut (.I0(n990), .I1(n1043), 
            .I2(n1012), .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i674_3_lut (.I0(n986), .I1(n1039), 
            .I2(n1012), .I3(GND_net), .O(n1064));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i675_3_lut (.I0(n987), .I1(n1040), 
            .I2(n1012), .I3(GND_net), .O(n1065));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i684_3_lut (.I0(n432), .I1(n1049), 
            .I2(n1012), .I3(GND_net), .O(n1074));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i684_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i683_3_lut (.I0(n995), .I1(n1048), 
            .I2(n1012), .I3(GND_net), .O(n1073));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_2782_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4517), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n433));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17784_3_lut (.I0(n433), .I1(n1073), .I2(n1074), .I3(GND_net), 
            .O(n21885));
    defparam i17784_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1666 (.I0(n1071), .I1(n1070), .I2(n21885), .I3(n1072), 
            .O(n30785));
    defparam i2_4_lut_adj_1666.LUT_INIT = 16'h8880;
    SB_LUT4 i5_4_lut_adj_1667 (.I0(n1065), .I1(n1064), .I2(n30785), .I3(n1068), 
            .O(n12_adj_4655));
    defparam i5_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i28556_4_lut (.I0(n1067), .I1(n12_adj_4655), .I2(n1066), .I3(n1069), 
            .O(n1090));
    defparam i28556_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1482_3_lut (.I0(n1090), .I1(n4667), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[13]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1482_3_lut.LUT_INIT = 16'hc5c5;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_i622_3_lut (.I0(n909), .I1(n962), 
            .I2(n934), .I3(GND_net), .O(n987));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i622_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n25059), .I0(encoder1_position[6]), 
            .I1(n19_adj_4549), .CO(n25060));
    SB_LUT4 encoder0_position_23__I_0_i623_3_lut (.I0(n910), .I1(n963), 
            .I2(n934), .I3(GND_net), .O(n988));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i623_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i630_3_lut (.I0(n431), .I1(n970), 
            .I2(n934), .I3(GND_net), .O(n995));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i630_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4550), .I3(n25058), .O(displacement_23__N_50[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i629_3_lut (.I0(n916), .I1(n969), 
            .I2(n934), .I3(GND_net), .O(n994));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i629_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i628_3_lut (.I0(n915), .I1(n968), 
            .I2(n934), .I3(GND_net), .O(n993));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i628_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n25058), .I0(encoder1_position[5]), 
            .I1(n20_adj_4550), .CO(n25059));
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4551), .I3(n25057), .O(displacement_23__N_50[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n25057), .I0(encoder1_position[4]), 
            .I1(n21_adj_4551), .CO(n25058));
    SB_LUT4 mux_2782_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4518), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n432));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4552), .I3(n25056), .O(displacement_23__N_50[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i626_3_lut (.I0(n913), .I1(n966), 
            .I2(n934), .I3(GND_net), .O(n991));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i626_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n25056), .I0(encoder1_position[3]), 
            .I1(n22_adj_4552), .CO(n25057));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4553), .I3(n25055), .O(displacement_23__N_50[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i627_3_lut (.I0(n914), .I1(n967), 
            .I2(n934), .I3(GND_net), .O(n992));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i627_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i625_3_lut (.I0(n912), .I1(n965), 
            .I2(n934), .I3(GND_net), .O(n990));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i621_3_lut (.I0(n908), .I1(n961), 
            .I2(n934), .I3(GND_net), .O(n986));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i624_3_lut (.I0(n911), .I1(n964), 
            .I2(n934), .I3(GND_net), .O(n989));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i624_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n25055), .I0(encoder1_position[2]), 
            .I1(n23_adj_4553), .CO(n25056));
    SB_LUT4 i17951_4_lut (.I0(n432), .I1(n993), .I2(n994), .I3(n995), 
            .O(n22053));
    defparam i17951_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i13002_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n12944), .I3(GND_net), .O(n17111));   // verilog/coms.v(127[12] 300[6])
    defparam i13002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4554), .I3(n25054), .O(displacement_23__N_50[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n25054), .I0(encoder1_position[1]), 
            .I1(n24_adj_4554), .CO(n25055));
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4540));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i520_3_lut (.I0(n757), .I1(n810), 
            .I2(n778), .I3(GND_net), .O(n835));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13003_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n12944), .I3(GND_net), .O(n17112));   // verilog/coms.v(127[12] 300[6])
    defparam i13003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4555), .I3(VCC_net), .O(displacement_23__N_50[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4555), .CO(n25054));
    SB_LUT4 i2_2_lut_adj_1668 (.I0(n989), .I1(n986), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4620));
    defparam i2_2_lut_adj_1668.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1669 (.I0(n990), .I1(n992), .I2(n991), .I3(n22053), 
            .O(n7_adj_4621));
    defparam i1_4_lut_adj_1669.LUT_INIT = 16'heaaa;
    SB_LUT4 i28788_4_lut (.I0(n988), .I1(n7_adj_4621), .I2(n987), .I3(n8_adj_4620), 
            .O(n1012));
    defparam i28788_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1481_3_lut (.I0(n1012), .I1(n4666), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[14]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1481_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i570_3_lut (.I0(n832), .I1(n885), 
            .I2(n856), .I3(GND_net), .O(n910));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i569_3_lut (.I0(n831), .I1(n884), 
            .I2(n856), .I3(GND_net), .O(n909));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13004_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n12944), .I3(GND_net), .O(n17113));   // verilog/coms.v(127[12] 300[6])
    defparam i13004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i571_3_lut (.I0(n833), .I1(n886), 
            .I2(n856), .I3(GND_net), .O(n911));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i571_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i576_3_lut (.I0(n430), .I1(n891), 
            .I2(n856), .I3(GND_net), .O(n916));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i575_3_lut (.I0(n837), .I1(n890), 
            .I2(n856), .I3(GND_net), .O(n915));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13005_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n12944), .I3(GND_net), .O(n17114));   // verilog/coms.v(127[12] 300[6])
    defparam i13005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i574_3_lut (.I0(n836), .I1(n889), 
            .I2(n856), .I3(GND_net), .O(n914));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13006_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n12944), .I3(GND_net), .O(n17115));   // verilog/coms.v(127[12] 300[6])
    defparam i13006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2782_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4519), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n431));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4614));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i572_3_lut (.I0(n834), .I1(n887), 
            .I2(n856), .I3(GND_net), .O(n912));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4613));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13007_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n12944), .I3(GND_net), .O(n17116));   // verilog/coms.v(127[12] 300[6])
    defparam i13007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4612));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i568_3_lut (.I0(n830), .I1(n883), 
            .I2(n856), .I3(GND_net), .O(n908));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i573_3_lut (.I0(n835), .I1(n888), 
            .I2(n856), .I3(GND_net), .O(n913));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17955_4_lut (.I0(n431), .I1(n914), .I2(n915), .I3(n916), 
            .O(n22057));
    defparam i17955_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4611));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_adj_1670 (.I0(n913), .I1(n908), .I2(n912), .I3(n22057), 
            .O(n7_adj_4615));
    defparam i2_4_lut_adj_1670.LUT_INIT = 16'heccc;
    SB_LUT4 i28766_4_lut (.I0(n7_adj_4615), .I1(n911), .I2(n909), .I3(n910), 
            .O(n934));
    defparam i28766_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1480_3_lut (.I0(n934), .I1(n4665), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[15]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1480_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i516_3_lut (.I0(n753), .I1(n806), 
            .I2(n778), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i517_3_lut (.I0(n754), .I1(n807), 
            .I2(n778), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i518_3_lut (.I0(n755), .I1(n808), 
            .I2(n778), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17844_3_lut (.I0(n430), .I1(n836), .I2(n837), .I3(GND_net), 
            .O(n21945));
    defparam i17844_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1671 (.I0(n834), .I1(n833), .I2(n21945), .I3(n835), 
            .O(n31461));
    defparam i2_4_lut_adj_1671.LUT_INIT = 16'h8880;
    SB_LUT4 i28404_4_lut (.I0(n31461), .I1(n830), .I2(n832), .I3(n831), 
            .O(n856));
    defparam i28404_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1479_3_lut (.I0(n856), .I1(n4664), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[16]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1479_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1478_3_lut (.I0(n778), .I1(n4663), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[17]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1478_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1477_3_lut (.I0(n700), .I1(n4662), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[18]));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i1477_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4591));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13008_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n12944), .I3(GND_net), .O(n17117));   // verilog/coms.v(127[12] 300[6])
    defparam i13008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13009_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n12944), .I3(GND_net), .O(n17118));   // verilog/coms.v(127[12] 300[6])
    defparam i13009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12793_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4216), .I3(GND_net), .O(n16902));   // verilog/coms.v(127[12] 300[6])
    defparam i12793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13010_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n12944), .I3(GND_net), .O(n17119));   // verilog/coms.v(127[12] 300[6])
    defparam i13010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13011_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n12944), .I3(GND_net), .O(n17120));   // verilog/coms.v(127[12] 300[6])
    defparam i13011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13012_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n12944), .I3(GND_net), .O(n17121));   // verilog/coms.v(127[12] 300[6])
    defparam i13012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12794_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4216), .I3(GND_net), .O(n16903));   // verilog/coms.v(127[12] 300[6])
    defparam i12794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13013_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n12944), .I3(GND_net), .O(n17122));   // verilog/coms.v(127[12] 300[6])
    defparam i13013_3_lut.LUT_INIT = 16'hcaca;
    SB_IO SCL_pad (.PACKAGE_PIN(SCL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCL_pad.PIN_TYPE = 6'b011001;
    defparam SCL_pad.PULLUP = 1'b0;
    defparam SCL_pad.NEG_TRIGGER = 1'b0;
    defparam SCL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13014_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n12944), .I3(GND_net), .O(n17123));   // verilog/coms.v(127[12] 300[6])
    defparam i13014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13015_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n12944), .I3(GND_net), .O(n17124));   // verilog/coms.v(127[12] 300[6])
    defparam i13015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_41_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[15]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13016_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n12944), .I3(GND_net), .O(n17125));   // verilog/coms.v(127[12] 300[6])
    defparam i13016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13017_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n12944), .I3(GND_net), .O(n17126));   // verilog/coms.v(127[12] 300[6])
    defparam i13017_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13018_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n12944), .I3(GND_net), .O(n17127));   // verilog/coms.v(127[12] 300[6])
    defparam i13018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4488));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13019_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n12944), .I3(GND_net), .O(n17128));   // verilog/coms.v(127[12] 300[6])
    defparam i13019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12795_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n29532), .I3(GND_net), .O(n16904));   // verilog/coms.v(127[12] 300[6])
    defparam i12795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13020_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n12944), .I3(GND_net), .O(n17129));   // verilog/coms.v(127[12] 300[6])
    defparam i13020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1354_7_lut (.I0(GND_net), .I1(n509), .I2(GND_net), .I3(n24951), 
            .O(n4429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1354_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13021_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n12944), .I3(GND_net), .O(n17130));   // verilog/coms.v(127[12] 300[6])
    defparam i13021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13022_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n12944), .I3(GND_net), .O(n17131));   // verilog/coms.v(127[12] 300[6])
    defparam i13022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13023_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n12944), .I3(GND_net), .O(n17132));   // verilog/coms.v(127[12] 300[6])
    defparam i13023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13024_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n12944), .I3(GND_net), .O(n17133));   // verilog/coms.v(127[12] 300[6])
    defparam i13024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13025_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n12944), .I3(GND_net), .O(n17134));   // verilog/coms.v(127[12] 300[6])
    defparam i13025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13026_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n12944), .I3(GND_net), .O(n17135));   // verilog/coms.v(127[12] 300[6])
    defparam i13026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1354_6_lut (.I0(n32219), .I1(n510), .I2(GND_net), .I3(n24950), 
            .O(n33173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1354_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i13027_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n12944), .I3(GND_net), .O(n17136));   // verilog/coms.v(127[12] 300[6])
    defparam i13027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13028_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n12944), .I3(GND_net), .O(n17137));   // verilog/coms.v(127[12] 300[6])
    defparam i13028_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1354_6 (.CI(n24950), .I0(n510), .I1(GND_net), .CO(n24951));
    SB_LUT4 i13029_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n12944), .I3(GND_net), .O(n17138));   // verilog/coms.v(127[12] 300[6])
    defparam i13029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1354_5_lut (.I0(GND_net), .I1(n511), .I2(VCC_net), .I3(n24949), 
            .O(n4431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1354_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13030_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n12944), .I3(GND_net), .O(n17139));   // verilog/coms.v(127[12] 300[6])
    defparam i13030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13031_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n12944), .I3(GND_net), .O(n17140));   // verilog/coms.v(127[12] 300[6])
    defparam i13031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13032_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n12944), .I3(GND_net), .O(n17141));   // verilog/coms.v(127[12] 300[6])
    defparam i13032_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1354_5 (.CI(n24949), .I0(n511), .I1(VCC_net), .CO(n24950));
    SB_LUT4 add_1354_4_lut (.I0(GND_net), .I1(n425), .I2(GND_net), .I3(n24948), 
            .O(n4432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1354_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1354_4 (.CI(n24948), .I0(n425), .I1(GND_net), .CO(n24949));
    SB_LUT4 i13033_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n12944), .I3(GND_net), .O(n17142));   // verilog/coms.v(127[12] 300[6])
    defparam i13033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13034_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n12944), .I3(GND_net), .O(n17143));   // verilog/coms.v(127[12] 300[6])
    defparam i13034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13035_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n12944), .I3(GND_net), .O(n17144));   // verilog/coms.v(127[12] 300[6])
    defparam i13035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_41_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[16]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13036_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n12944), .I3(GND_net), .O(n17145));   // verilog/coms.v(127[12] 300[6])
    defparam i13036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13037_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n12944), .I3(GND_net), .O(n17146));   // verilog/coms.v(127[12] 300[6])
    defparam i13037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13038_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n12944), .I3(GND_net), .O(n17147));   // verilog/coms.v(127[12] 300[6])
    defparam i13038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12796_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n29532), .I3(GND_net), .O(n16905));   // verilog/coms.v(127[12] 300[6])
    defparam i12796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13039_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n12944), .I3(GND_net), .O(n17148));   // verilog/coms.v(127[12] 300[6])
    defparam i13039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13040_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n12944), .I3(GND_net), .O(n17149));   // verilog/coms.v(127[12] 300[6])
    defparam i13040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1354_3_lut (.I0(GND_net), .I1(n426), .I2(VCC_net), .I3(n24947), 
            .O(n4433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1354_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13041_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n12944), 
            .I3(GND_net), .O(n17150));   // verilog/coms.v(127[12] 300[6])
    defparam i13041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13042_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n12944), 
            .I3(GND_net), .O(n17151));   // verilog/coms.v(127[12] 300[6])
    defparam i13042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13043_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n12944), 
            .I3(GND_net), .O(n17152));   // verilog/coms.v(127[12] 300[6])
    defparam i13043_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1354_3 (.CI(n24947), .I0(n426), .I1(VCC_net), .CO(n24948));
    SB_LUT4 add_1354_2_lut (.I0(GND_net), .I1(n427), .I2(GND_net), .I3(VCC_net), 
            .O(n4434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1354_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13044_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n12944), 
            .I3(GND_net), .O(n17153));   // verilog/coms.v(127[12] 300[6])
    defparam i13044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13045_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n12944), 
            .I3(GND_net), .O(n17154));   // verilog/coms.v(127[12] 300[6])
    defparam i13045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13046_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n12944), 
            .I3(GND_net), .O(n17155));   // verilog/coms.v(127[12] 300[6])
    defparam i13046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13047_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n12944), 
            .I3(GND_net), .O(n17156));   // verilog/coms.v(127[12] 300[6])
    defparam i13047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13048_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n12944), 
            .I3(GND_net), .O(n17157));   // verilog/coms.v(127[12] 300[6])
    defparam i13048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13049_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n12944), 
            .I3(GND_net), .O(n17158));   // verilog/coms.v(127[12] 300[6])
    defparam i13049_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1354_2 (.CI(VCC_net), .I0(n427), .I1(GND_net), .CO(n24947));
    SB_LUT4 i13050_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n12944), 
            .I3(GND_net), .O(n17159));   // verilog/coms.v(127[12] 300[6])
    defparam i13050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i463_3_lut (.I0(n675), .I1(n728), 
            .I2(n700), .I3(GND_net), .O(n753));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i465_3_lut (.I0(n677), .I1(n730), 
            .I2(n700), .I3(GND_net), .O(n755));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i467_3_lut (.I0(n679), .I1(n732), 
            .I2(n700), .I3(GND_net), .O(n757));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i464_3_lut (.I0(n676), .I1(n729), 
            .I2(n700), .I3(GND_net), .O(n754));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_486_24_lut (.I0(duty[22]), .I1(n34501), .I2(n3), .I3(n24946), 
            .O(pwm_setpoint_22__N_3[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_24_lut.LUT_INIT = 16'h8BB8;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_50[23]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_LUT4 add_486_23_lut (.I0(duty[21]), .I1(n34501), .I2(n4_adj_4488), 
            .I3(n24945), .O(pwm_setpoint_22__N_3[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13051_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n12944), 
            .I3(GND_net), .O(n17160));   // verilog/coms.v(127[12] 300[6])
    defparam i13051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13052_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n12944), 
            .I3(GND_net), .O(n17161));   // verilog/coms.v(127[12] 300[6])
    defparam i13052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13053_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n12944), 
            .I3(GND_net), .O(n17162));   // verilog/coms.v(127[12] 300[6])
    defparam i13053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13054_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n12944), 
            .I3(GND_net), .O(n17163));   // verilog/coms.v(127[12] 300[6])
    defparam i13054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13055_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n12944), 
            .I3(GND_net), .O(n17164));   // verilog/coms.v(127[12] 300[6])
    defparam i13055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13056_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n12944), 
            .I3(GND_net), .O(n17165));   // verilog/coms.v(127[12] 300[6])
    defparam i13056_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_50[22]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_LUT4 i13057_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n12944), 
            .I3(GND_net), .O(n17166));   // verilog/coms.v(127[12] 300[6])
    defparam i13057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13058_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n12944), 
            .I3(GND_net), .O(n17167));   // verilog/coms.v(127[12] 300[6])
    defparam i13058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13059_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n12944), 
            .I3(GND_net), .O(n17168));   // verilog/coms.v(127[12] 300[6])
    defparam i13059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13060_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n12944), 
            .I3(GND_net), .O(n17169));   // verilog/coms.v(127[12] 300[6])
    defparam i13060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13061_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n12944), 
            .I3(GND_net), .O(n17170));   // verilog/coms.v(127[12] 300[6])
    defparam i13061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13062_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n12944), 
            .I3(GND_net), .O(n17171));   // verilog/coms.v(127[12] 300[6])
    defparam i13062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13063_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n12944), 
            .I3(GND_net), .O(n17172));   // verilog/coms.v(127[12] 300[6])
    defparam i13063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13064_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n12944), 
            .I3(GND_net), .O(n17173));   // verilog/coms.v(127[12] 300[6])
    defparam i13064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13065_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n12944), .I3(GND_net), .O(n17174));   // verilog/coms.v(127[12] 300[6])
    defparam i13065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13066_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n12944), .I3(GND_net), .O(n17175));   // verilog/coms.v(127[12] 300[6])
    defparam i13066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13067_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n12944), .I3(GND_net), .O(n17176));   // verilog/coms.v(127[12] 300[6])
    defparam i13067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13068_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n12944), .I3(GND_net), .O(n17177));   // verilog/coms.v(127[12] 300[6])
    defparam i13068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13069_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n12944), .I3(GND_net), .O(n17178));   // verilog/coms.v(127[12] 300[6])
    defparam i13069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13070_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n12944), .I3(GND_net), .O(n17179));   // verilog/coms.v(127[12] 300[6])
    defparam i13070_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_486_23 (.CI(n24945), .I0(n34501), .I1(n4_adj_4488), .CO(n24946));
    SB_LUT4 mux_2782_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4524), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n426));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13071_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n12944), .I3(GND_net), .O(n17180));   // verilog/coms.v(127[12] 300[6])
    defparam i13071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13072_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n12944), .I3(GND_net), .O(n17181));   // verilog/coms.v(127[12] 300[6])
    defparam i13072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_41_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[17]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13073_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n12944), .I3(GND_net), .O(n17182));   // verilog/coms.v(127[12] 300[6])
    defparam i13073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13074_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n12944), .I3(GND_net), .O(n17183));   // verilog/coms.v(127[12] 300[6])
    defparam i13074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13075_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n12944), .I3(GND_net), .O(n17184));   // verilog/coms.v(127[12] 300[6])
    defparam i13075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13076_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n12944), .I3(GND_net), .O(n17185));   // verilog/coms.v(127[12] 300[6])
    defparam i13076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13077_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n12944), .I3(GND_net), .O(n17186));   // verilog/coms.v(127[12] 300[6])
    defparam i13077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13078_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n12944), .I3(GND_net), .O(n17187));   // verilog/coms.v(127[12] 300[6])
    defparam i13078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13079_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n12944), .I3(GND_net), .O(n17188));   // verilog/coms.v(127[12] 300[6])
    defparam i13079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13080_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n12944), .I3(GND_net), .O(n17189));   // verilog/coms.v(127[12] 300[6])
    defparam i13080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13081_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n12944), .I3(GND_net), .O(n17190));   // verilog/coms.v(127[12] 300[6])
    defparam i13081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13082_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n12944), .I3(GND_net), .O(n17191));   // verilog/coms.v(127[12] 300[6])
    defparam i13082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13083_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n12944), .I3(GND_net), .O(n17192));   // verilog/coms.v(127[12] 300[6])
    defparam i13083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13084_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n12944), .I3(GND_net), .O(n17193));   // verilog/coms.v(127[12] 300[6])
    defparam i13084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13085_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n12944), .I3(GND_net), .O(n17194));   // verilog/coms.v(127[12] 300[6])
    defparam i13085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13086_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n12944), .I3(GND_net), .O(n17195));   // verilog/coms.v(127[12] 300[6])
    defparam i13086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13087_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n12944), .I3(GND_net), .O(n17196));   // verilog/coms.v(127[12] 300[6])
    defparam i13087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13088_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n12944), .I3(GND_net), .O(n17197));   // verilog/coms.v(127[12] 300[6])
    defparam i13088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13089_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n12944), .I3(GND_net), .O(n17198));   // verilog/coms.v(127[12] 300[6])
    defparam i13089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13090_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n12944), .I3(GND_net), .O(n17199));   // verilog/coms.v(127[12] 300[6])
    defparam i13090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13091_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n12944), .I3(GND_net), .O(n17200));   // verilog/coms.v(127[12] 300[6])
    defparam i13091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13092_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n12944), .I3(GND_net), .O(n17201));   // verilog/coms.v(127[12] 300[6])
    defparam i13092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13093_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n12944), .I3(GND_net), .O(n17202));   // verilog/coms.v(127[12] 300[6])
    defparam i13093_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_50[21]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_50[20]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_50[19]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_50[18]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_50[17]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_50[16]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_50[15]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_50[14]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_50[13]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_50[12]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_50[11]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_50[10]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_50[9]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_50[8]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_50[7]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_50[6]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_50[5]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_50[4]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_50[3]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_50[2]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_50[1]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFFSR encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
            .C(clk32MHz), .D(n4659), .R(n2_adj_4591));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFFSR encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
            .C(clk32MHz), .D(n4660), .R(n2_adj_4591));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[19]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[18]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[17]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[16]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[15]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[14]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[13]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[12]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[11]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[10]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[9]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[8]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[7]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[6]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[5]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[4]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[3]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[2]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[1]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[22]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[21]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[20]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[19]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[18]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[17]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[16]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[15]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[14]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[13]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[12]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[11]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[10]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[9]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[8]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[7]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[6]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[5]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[4]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[3]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[2]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[1]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 mux_2782_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4525), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n425));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13094_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n12944), .I3(GND_net), .O(n17203));   // verilog/coms.v(127[12] 300[6])
    defparam i13094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13095_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n12944), .I3(GND_net), .O(n17204));   // verilog/coms.v(127[12] 300[6])
    defparam i13095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_486_22_lut (.I0(duty[20]), .I1(n34501), .I2(n5), .I3(n24944), 
            .O(pwm_setpoint_22__N_3[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13096_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n12944), .I3(GND_net), .O(n17205));   // verilog/coms.v(127[12] 300[6])
    defparam i13096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13097_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n12944), .I3(GND_net), .O(n17206));   // verilog/coms.v(127[12] 300[6])
    defparam i13097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13098_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n12944), .I3(GND_net), .O(n17207));   // verilog/coms.v(127[12] 300[6])
    defparam i13098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13099_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n12944), .I3(GND_net), .O(n17208));   // verilog/coms.v(127[12] 300[6])
    defparam i13099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13100_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n12944), .I3(GND_net), .O(n17209));   // verilog/coms.v(127[12] 300[6])
    defparam i13100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13101_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n12944), .I3(GND_net), .O(n17210));   // verilog/coms.v(127[12] 300[6])
    defparam i13101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13102_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n12944), .I3(GND_net), .O(n17211));   // verilog/coms.v(127[12] 300[6])
    defparam i13102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13103_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n12944), .I3(GND_net), .O(n17212));   // verilog/coms.v(127[12] 300[6])
    defparam i13103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2782_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4526), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_41_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[18]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13104_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n12944), .I3(GND_net), .O(n17213));   // verilog/coms.v(127[12] 300[6])
    defparam i13104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13105_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n12944), .I3(GND_net), .O(n17214));   // verilog/coms.v(127[12] 300[6])
    defparam i13105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13106_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n12944), .I3(GND_net), .O(n17215));   // verilog/coms.v(127[12] 300[6])
    defparam i13106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26546_1_lut (.I0(n4_adj_4625), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n32219));
    defparam i26546_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_2782_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4527), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n510));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13107_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n12944), .I3(GND_net), .O(n17216));   // verilog/coms.v(127[12] 300[6])
    defparam i13107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3383_2_lut (.I0(n2), .I1(encoder0_position[23]), .I2(GND_net), 
            .I3(GND_net), .O(n509));
    defparam i3383_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24632_4_lut (.I0(encoder0_position[22]), .I1(n33173), .I2(encoder0_position[23]), 
            .I3(n3_adj_4527), .O(n675));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam i24632_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY add_486_22 (.CI(n24944), .I0(n34501), .I1(n5), .CO(n24945));
    SB_LUT4 mux_41_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[19]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i24630_3_lut (.I0(encoder0_position[21]), .I1(n30290), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n676));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam i24630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13108_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n12944), .I3(GND_net), .O(n17217));   // verilog/coms.v(127[12] 300[6])
    defparam i13108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13109_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n12944), .I3(GND_net), .O(n17218));   // verilog/coms.v(127[12] 300[6])
    defparam i13109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_41_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[20]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13110_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n12944), .I3(GND_net), .O(n17219));   // verilog/coms.v(127[12] 300[6])
    defparam i13110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12797_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n29532), .I3(GND_net), .O(n16906));   // verilog/coms.v(127[12] 300[6])
    defparam i12797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13111_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n12944), .I3(GND_net), .O(n17220));   // verilog/coms.v(127[12] 300[6])
    defparam i13111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13112_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n12944), .I3(GND_net), .O(n17221));   // verilog/coms.v(127[12] 300[6])
    defparam i13112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13113_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n12944), .I3(GND_net), .O(n17222));   // verilog/coms.v(127[12] 300[6])
    defparam i13113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13114_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n12944), .I3(GND_net), .O(n17223));   // verilog/coms.v(127[12] 300[6])
    defparam i13114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13115_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n12944), .I3(GND_net), .O(n17224));   // verilog/coms.v(127[12] 300[6])
    defparam i13115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13116_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n12944), .I3(GND_net), .O(n17225));   // verilog/coms.v(127[12] 300[6])
    defparam i13116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13117_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n12944), .I3(GND_net), .O(n17226));   // verilog/coms.v(127[12] 300[6])
    defparam i13117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2782_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4523), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n427));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13118_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n12944), .I3(GND_net), .O(n17227));   // verilog/coms.v(127[12] 300[6])
    defparam i13118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13119_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n12944), .I3(GND_net), .O(n17228));   // verilog/coms.v(127[12] 300[6])
    defparam i13119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13120_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n12944), .I3(GND_net), .O(n17229));   // verilog/coms.v(127[12] 300[6])
    defparam i13120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13121_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n12944), .I3(GND_net), .O(n17230));   // verilog/coms.v(127[12] 300[6])
    defparam i13121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13122_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n12944), .I3(GND_net), .O(n17231));   // verilog/coms.v(127[12] 300[6])
    defparam i13122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13123_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n12944), .I3(GND_net), .O(n17232));   // verilog/coms.v(127[12] 300[6])
    defparam i13123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13124_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n12944), .I3(GND_net), .O(n17233));   // verilog/coms.v(127[12] 300[6])
    defparam i13124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13125_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n12944), .I3(GND_net), .O(n17234));   // verilog/coms.v(127[12] 300[6])
    defparam i13125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13126_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n12944), .I3(GND_net), .O(n17235));   // verilog/coms.v(127[12] 300[6])
    defparam i13126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13127_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n12944), .I3(GND_net), .O(n17236));   // verilog/coms.v(127[12] 300[6])
    defparam i13127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13128_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n12944), .I3(GND_net), .O(n17237));   // verilog/coms.v(127[12] 300[6])
    defparam i13128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13129_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[22]), 
            .I2(n12944), .I3(GND_net), .O(n17238));   // verilog/coms.v(127[12] 300[6])
    defparam i13129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13130_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n12944), .I3(GND_net), .O(n17239));   // verilog/coms.v(127[12] 300[6])
    defparam i13130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13131_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[22]), 
            .I2(n12944), .I3(GND_net), .O(n17240));   // verilog/coms.v(127[12] 300[6])
    defparam i13131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13132_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n12944), .I3(GND_net), .O(n17241));   // verilog/coms.v(127[12] 300[6])
    defparam i13132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13133_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n12944), .I3(GND_net), .O(n17242));   // verilog/coms.v(127[12] 300[6])
    defparam i13133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13134_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n12944), .I3(GND_net), .O(n17243));   // verilog/coms.v(127[12] 300[6])
    defparam i13134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13135_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n12944), .I3(GND_net), .O(n17244));   // verilog/coms.v(127[12] 300[6])
    defparam i13135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13136_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n12944), .I3(GND_net), .O(n17245));   // verilog/coms.v(127[12] 300[6])
    defparam i13136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13137_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n12944), .I3(GND_net), .O(n17246));   // verilog/coms.v(127[12] 300[6])
    defparam i13137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13138_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n12944), .I3(GND_net), .O(n17247));   // verilog/coms.v(127[12] 300[6])
    defparam i13138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13139_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n12944), .I3(GND_net), .O(n17248));   // verilog/coms.v(127[12] 300[6])
    defparam i13139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13140_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n12944), .I3(GND_net), .O(n17249));   // verilog/coms.v(127[12] 300[6])
    defparam i13140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13141_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n12944), .I3(GND_net), .O(n17250));   // verilog/coms.v(127[12] 300[6])
    defparam i13141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13142_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n12944), .I3(GND_net), .O(n17251));   // verilog/coms.v(127[12] 300[6])
    defparam i13142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13143_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n12944), .I3(GND_net), .O(n17252));   // verilog/coms.v(127[12] 300[6])
    defparam i13143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13144_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n12944), .I3(GND_net), .O(n17253));   // verilog/coms.v(127[12] 300[6])
    defparam i13144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13145_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n8868), 
            .I3(GND_net), .O(n17254));   // verilog/coms.v(127[12] 300[6])
    defparam i13145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_41_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[21]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13146_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n8868), 
            .I3(GND_net), .O(n17255));   // verilog/coms.v(127[12] 300[6])
    defparam i13146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13147_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n8868), 
            .I3(GND_net), .O(n17256));   // verilog/coms.v(127[12] 300[6])
    defparam i13147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1672 (.I0(n427), .I1(n6_adj_4524), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4502));
    defparam i1_2_lut_adj_1672.LUT_INIT = 16'heeee;
    SB_LUT4 i13148_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n8868), 
            .I3(GND_net), .O(n17257));   // verilog/coms.v(127[12] 300[6])
    defparam i13148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13149_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n8868), 
            .I3(GND_net), .O(n17258));   // verilog/coms.v(127[12] 300[6])
    defparam i13149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_486_21_lut (.I0(duty[19]), .I1(n34501), .I2(n6), .I3(n24943), 
            .O(pwm_setpoint_22__N_3[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_486_21 (.CI(n24943), .I0(n34501), .I1(n6), .CO(n24944));
    SB_LUT4 add_486_20_lut (.I0(duty[18]), .I1(n34501), .I2(n7), .I3(n24942), 
            .O(pwm_setpoint_22__N_3[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_486_20 (.CI(n24942), .I0(n34501), .I1(n7), .CO(n24943));
    SB_LUT4 i13150_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n8868), 
            .I3(GND_net), .O(n17259));   // verilog/coms.v(127[12] 300[6])
    defparam i13150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13151_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n8868), 
            .I3(GND_net), .O(n17260));   // verilog/coms.v(127[12] 300[6])
    defparam i13151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_486_19_lut (.I0(duty[17]), .I1(n34501), .I2(n8), .I3(n24941), 
            .O(pwm_setpoint_22__N_3[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_19_lut.LUT_INIT = 16'h8BB8;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13152_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n8868), 
            .I3(GND_net), .O(n17261));   // verilog/coms.v(127[12] 300[6])
    defparam i13152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(n4_adj_4526), .I1(n2), .I2(n5_adj_4525), 
            .I3(n7_adj_4502), .O(n4_adj_4625));
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'hc888;
    SB_LUT4 i13153_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n8868), 
            .I3(GND_net), .O(n17262));   // verilog/coms.v(127[12] 300[6])
    defparam i13153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13154_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n8868), 
            .I3(GND_net), .O(n17263));   // verilog/coms.v(127[12] 300[6])
    defparam i13154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13155_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n8868), 
            .I3(GND_net), .O(n17264));   // verilog/coms.v(127[12] 300[6])
    defparam i13155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_26_lut (.I0(GND_net), .I1(n2000), 
            .I2(VCC_net), .I3(n25421), .O(n2053)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_558_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4568));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13156_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n8868), 
            .I3(GND_net), .O(n17265));   // verilog/coms.v(127[12] 300[6])
    defparam i13156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13157_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n8868), 
            .I3(GND_net), .O(n17266));   // verilog/coms.v(127[12] 300[6])
    defparam i13157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_25_lut (.I0(GND_net), .I1(n2001), 
            .I2(VCC_net), .I3(n25420), .O(n2054)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_25 (.CI(n25420), .I0(n2001), 
            .I1(VCC_net), .CO(n25421));
    SB_LUT4 encoder0_position_23__I_0_add_1361_24_lut (.I0(GND_net), .I1(n2002), 
            .I2(VCC_net), .I3(n25419), .O(n2055)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_558_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4572));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_1361_24 (.CI(n25419), .I0(n2002), 
            .I1(VCC_net), .CO(n25420));
    SB_LUT4 i13158_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n8868), 
            .I3(GND_net), .O(n17267));   // verilog/coms.v(127[12] 300[6])
    defparam i13158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_23_lut (.I0(GND_net), .I1(n2003), 
            .I2(VCC_net), .I3(n25418), .O(n2056)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_23 (.CI(n25418), .I0(n2003), 
            .I1(VCC_net), .CO(n25419));
    SB_LUT4 i27559_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n33233));
    defparam i27559_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_558_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4574));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13159_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n8868), 
            .I3(GND_net), .O(n17268));   // verilog/coms.v(127[12] 300[6])
    defparam i13159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_558_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4570));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i27573_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n33247));
    defparam i27573_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.i_31__N_2364 ), .I1(n63_adj_4566), 
            .I2(n771), .I3(n2_adj_4638), .O(n5_adj_4639));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hcc08;
    SB_LUT4 encoder0_position_23__I_0_add_1361_22_lut (.I0(GND_net), .I1(n2004), 
            .I2(VCC_net), .I3(n25417), .O(n2057)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_22 (.CI(n25417), .I0(n2004), 
            .I1(VCC_net), .CO(n25418));
    SB_LUT4 encoder0_position_23__I_0_add_1361_21_lut (.I0(GND_net), .I1(n2005), 
            .I2(VCC_net), .I3(n25416), .O(n2058)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_21 (.CI(n25416), .I0(n2005), 
            .I1(VCC_net), .CO(n25417));
    SB_LUT4 i13160_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n8868), 
            .I3(GND_net), .O(n17269));   // verilog/coms.v(127[12] 300[6])
    defparam i13160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24624_3_lut (.I0(encoder0_position[18]), .I1(n30284), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n679));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam i24624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_20_lut (.I0(GND_net), .I1(n2006), 
            .I2(VCC_net), .I3(n25415), .O(n2059)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13161_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n8868), 
            .I3(GND_net), .O(n17270));   // verilog/coms.v(127[12] 300[6])
    defparam i13161_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_20 (.CI(n25415), .I0(n2006), 
            .I1(VCC_net), .CO(n25416));
    SB_LUT4 encoder0_position_23__I_0_add_1361_19_lut (.I0(GND_net), .I1(n2007), 
            .I2(VCC_net), .I3(n25414), .O(n2060)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_19 (.CI(n25414), .I0(n2007), 
            .I1(VCC_net), .CO(n25415));
    SB_LUT4 encoder0_position_23__I_0_add_1361_18_lut (.I0(GND_net), .I1(n2008), 
            .I2(VCC_net), .I3(n25413), .O(n2061)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_18 (.CI(n25413), .I0(n2008), 
            .I1(VCC_net), .CO(n25414));
    SB_LUT4 encoder0_position_23__I_0_add_1361_17_lut (.I0(GND_net), .I1(n2009), 
            .I2(VCC_net), .I3(n25412), .O(n2062)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_17 (.CI(n25412), .I0(n2009), 
            .I1(VCC_net), .CO(n25413));
    SB_LUT4 i13162_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n8868), 
            .I3(GND_net), .O(n17271));   // verilog/coms.v(127[12] 300[6])
    defparam i13162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_16_lut (.I0(GND_net), .I1(n2010), 
            .I2(VCC_net), .I3(n25411), .O(n2063)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_16 (.CI(n25411), .I0(n2010), 
            .I1(VCC_net), .CO(n25412));
    SB_LUT4 encoder0_position_23__I_0_add_1361_15_lut (.I0(GND_net), .I1(n2011), 
            .I2(VCC_net), .I3(n25410), .O(n2064)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_15 (.CI(n25410), .I0(n2011), 
            .I1(VCC_net), .CO(n25411));
    SB_LUT4 encoder0_position_23__I_0_add_1361_14_lut (.I0(GND_net), .I1(n2012), 
            .I2(VCC_net), .I3(n25409), .O(n2065)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_14 (.CI(n25409), .I0(n2012), 
            .I1(VCC_net), .CO(n25410));
    SB_LUT4 i13163_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n8868), 
            .I3(GND_net), .O(n17272));   // verilog/coms.v(127[12] 300[6])
    defparam i13163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24626_3_lut (.I0(encoder0_position[19]), .I1(n30286), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n678));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam i24626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13164_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n8868), 
            .I3(GND_net), .O(n17273));   // verilog/coms.v(127[12] 300[6])
    defparam i13164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13165_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n8868), 
            .I3(GND_net), .O(n17274));   // verilog/coms.v(127[12] 300[6])
    defparam i13165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_13_lut (.I0(GND_net), .I1(n2013), 
            .I2(VCC_net), .I3(n25408), .O(n2066)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_13 (.CI(n25408), .I0(n2013), 
            .I1(VCC_net), .CO(n25409));
    SB_LUT4 encoder0_position_23__I_0_add_1361_12_lut (.I0(GND_net), .I1(n2014), 
            .I2(VCC_net), .I3(n25407), .O(n2067)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_12 (.CI(n25407), .I0(n2014), 
            .I1(VCC_net), .CO(n25408));
    SB_LUT4 i13166_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n8868), 
            .I3(GND_net), .O(n17275));   // verilog/coms.v(127[12] 300[6])
    defparam i13166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13167_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n8868), 
            .I3(GND_net), .O(n17276));   // verilog/coms.v(127[12] 300[6])
    defparam i13167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_11_lut (.I0(GND_net), .I1(n2015), 
            .I2(VCC_net), .I3(n25406), .O(n2068)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24628_3_lut (.I0(encoder0_position[20]), .I1(n30288), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n677));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam i24628_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_486_19 (.CI(n24941), .I0(n34501), .I1(n8), .CO(n24942));
    SB_LUT4 i17981_4_lut (.I0(n428), .I1(n677), .I2(n678), .I3(n679), 
            .O(n22083));
    defparam i17981_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_23__I_0_add_1361_11 (.CI(n25406), .I0(n2015), 
            .I1(VCC_net), .CO(n25407));
    SB_LUT4 encoder0_position_23__I_0_add_1361_10_lut (.I0(GND_net), .I1(n2016), 
            .I2(VCC_net), .I3(n25405), .O(n2069)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_10 (.CI(n25405), .I0(n2016), 
            .I1(VCC_net), .CO(n25406));
    SB_LUT4 encoder0_position_23__I_0_add_1361_9_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n25404), .O(n2070)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_9 (.CI(n25404), .I0(n2017), 
            .I1(VCC_net), .CO(n25405));
    SB_LUT4 encoder0_position_23__I_0_add_1361_8_lut (.I0(GND_net), .I1(n2018), 
            .I2(GND_net), .I3(n25403), .O(n2071)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_8 (.CI(n25403), .I0(n2018), 
            .I1(GND_net), .CO(n25404));
    SB_LUT4 encoder0_position_23__I_0_add_1361_7_lut (.I0(n2073), .I1(n2019), 
            .I2(GND_net), .I3(n25402), .O(n33199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_23__I_0_add_1361_7 (.CI(n25402), .I0(n2019), 
            .I1(GND_net), .CO(n25403));
    SB_LUT4 i13168_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n8868), 
            .I3(GND_net), .O(n17277));   // verilog/coms.v(127[12] 300[6])
    defparam i13168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_6_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n25401), .O(n2073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13169_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n8868), 
            .I3(GND_net), .O(n17278));   // verilog/coms.v(127[12] 300[6])
    defparam i13169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28391_4_lut (.I0(n676), .I1(n674), .I2(n675), .I3(n22083), 
            .O(n700));
    defparam i28391_4_lut.LUT_INIT = 16'h1333;
    SB_LUT4 i13170_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n8868), 
            .I3(GND_net), .O(n17279));   // verilog/coms.v(127[12] 300[6])
    defparam i13170_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_6 (.CI(n25401), .I0(n2020), 
            .I1(VCC_net), .CO(n25402));
    SB_LUT4 i13171_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n8868), 
            .I3(GND_net), .O(n17280));   // verilog/coms.v(127[12] 300[6])
    defparam i13171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_5_lut (.I0(n6_adj_4657), .I1(n2021), 
            .I2(GND_net), .I3(n25400), .O(n33155)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_5_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mux_40_i1_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_23__I_0_add_1361_5 (.CI(n25400), .I0(n2021), 
            .I1(GND_net), .CO(n25401));
    SB_LUT4 i13172_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n8868), 
            .I3(GND_net), .O(n17281));   // verilog/coms.v(127[12] 300[6])
    defparam i13172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_4_lut (.I0(n2076), .I1(n2022), 
            .I2(VCC_net), .I3(n25399), .O(n6_adj_4657)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_23__I_0_add_1361_4 (.CI(n25399), .I0(n2022), 
            .I1(VCC_net), .CO(n25400));
    SB_LUT4 i13173_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n8868), 
            .I3(GND_net), .O(n17282));   // verilog/coms.v(127[12] 300[6])
    defparam i13173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_40_i2_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_add_1361_3_lut (.I0(GND_net), .I1(n445), 
            .I2(GND_net), .I3(n25398), .O(n2076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_3 (.CI(n25398), .I0(n445), 
            .I1(GND_net), .CO(n25399));
    SB_CARRY encoder0_position_23__I_0_add_1361_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n25398));
    SB_LUT4 add_1400_23_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n25397), .O(n4659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_2782_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4522), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n428));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1400_22_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n25396), .O(n4660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i468_3_lut (.I0(n428), .I1(n733), 
            .I2(n700), .I3(GND_net), .O(n758));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i468_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1400_22 (.CI(n25396), .I0(GND_net), .I1(VCC_net), .CO(n25397));
    SB_LUT4 add_1400_21_lut (.I0(encoder0_position[23]), .I1(GND_net), .I2(n619), 
            .I3(n25395), .O(encoder0_position_scaled_23__N_26[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13174_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n8868), 
            .I3(GND_net), .O(n17283));   // verilog/coms.v(127[12] 300[6])
    defparam i13174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13175_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17284));   // verilog/coms.v(127[12] 300[6])
    defparam i13175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_486_18_lut (.I0(duty[16]), .I1(n34501), .I2(n9), .I3(n24940), 
            .O(pwm_setpoint_22__N_3[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1400_21 (.CI(n25395), .I0(GND_net), .I1(n619), .CO(n25396));
    SB_LUT4 mux_2782_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4521), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n429));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam mux_2782_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1400_20_lut (.I0(GND_net), .I1(GND_net), .I2(n700), .I3(n25394), 
            .O(n4662)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_20 (.CI(n25394), .I0(GND_net), .I1(n700), .CO(n25395));
    SB_LUT4 i17696_2_lut (.I0(n429), .I1(n758), .I2(GND_net), .I3(GND_net), 
            .O(n21796));
    defparam i17696_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_1400_19_lut (.I0(GND_net), .I1(GND_net), .I2(n778), .I3(n25393), 
            .O(n4663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13176_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17285));   // verilog/coms.v(127[12] 300[6])
    defparam i13176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(n754), .I1(n21796), .I2(n756), .I3(n757), 
            .O(n4_adj_4640));
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'ha8a0;
    SB_CARRY add_1400_19 (.CI(n25393), .I0(GND_net), .I1(n778), .CO(n25394));
    SB_LUT4 i13177_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17286));   // verilog/coms.v(127[12] 300[6])
    defparam i13177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13178_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17287));   // verilog/coms.v(127[12] 300[6])
    defparam i13178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13179_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17288));   // verilog/coms.v(127[12] 300[6])
    defparam i13179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_40_i3_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 add_1400_18_lut (.I0(GND_net), .I1(GND_net), .I2(n856), .I3(n25392), 
            .O(n4664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_18 (.CI(n25392), .I0(GND_net), .I1(n856), .CO(n25393));
    SB_LUT4 add_1400_17_lut (.I0(GND_net), .I1(GND_net), .I2(n934), .I3(n25391), 
            .O(n4665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_17 (.CI(n25391), .I0(GND_net), .I1(n934), .CO(n25392));
    SB_LUT4 add_1400_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1012), .I3(n25390), 
            .O(n4666)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13180_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17289));   // verilog/coms.v(127[12] 300[6])
    defparam i13180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13181_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17290));   // verilog/coms.v(127[12] 300[6])
    defparam i13181_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1400_16 (.CI(n25390), .I0(GND_net), .I1(n1012), .CO(n25391));
    SB_LUT4 i13182_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17291));   // verilog/coms.v(127[12] 300[6])
    defparam i13182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_40_i4_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_40_i5_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 add_1400_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1090), .I3(n25389), 
            .O(n4667)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13183_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17292));   // verilog/coms.v(127[12] 300[6])
    defparam i13183_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1400_15 (.CI(n25389), .I0(GND_net), .I1(n1090), .CO(n25390));
    SB_LUT4 mux_40_i6_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 add_1400_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1168), .I3(n25388), 
            .O(n4668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_40_i7_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY add_1400_14 (.CI(n25388), .I0(GND_net), .I1(n1168), .CO(n25389));
    SB_LUT4 add_1400_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1246), .I3(n25387), 
            .O(n4669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_13 (.CI(n25387), .I0(GND_net), .I1(n1246), .CO(n25388));
    SB_LUT4 i13184_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17293));   // verilog/coms.v(127[12] 300[6])
    defparam i13184_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_486_18 (.CI(n24940), .I0(n34501), .I1(n9), .CO(n24941));
    SB_LUT4 i13185_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17294));   // verilog/coms.v(127[12] 300[6])
    defparam i13185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1400_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1324), .I3(n25386), 
            .O(n4670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_12 (.CI(n25386), .I0(GND_net), .I1(n1324), .CO(n25387));
    SB_LUT4 add_1400_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1402), .I3(n25385), 
            .O(n4671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13186_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17295));   // verilog/coms.v(127[12] 300[6])
    defparam i13186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13187_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17296));   // verilog/coms.v(127[12] 300[6])
    defparam i13187_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1400_11 (.CI(n25385), .I0(GND_net), .I1(n1402), .CO(n25386));
    SB_LUT4 add_1400_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1480), .I3(n25384), 
            .O(n4672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_486_17_lut (.I0(duty[15]), .I1(n34501), .I2(n10), .I3(n24939), 
            .O(pwm_setpoint_22__N_3[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1400_10 (.CI(n25384), .I0(GND_net), .I1(n1480), .CO(n25385));
    SB_LUT4 add_1400_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1558), .I3(n25383), 
            .O(n4673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_9 (.CI(n25383), .I0(GND_net), .I1(n1558), .CO(n25384));
    SB_LUT4 i13188_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17297));   // verilog/coms.v(127[12] 300[6])
    defparam i13188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1400_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1636), .I3(n25382), 
            .O(n4674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13189_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17298));   // verilog/coms.v(127[12] 300[6])
    defparam i13189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13190_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17299));   // verilog/coms.v(127[12] 300[6])
    defparam i13190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_40_i8_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i13191_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17300));   // verilog/coms.v(127[12] 300[6])
    defparam i13191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13192_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17301));   // verilog/coms.v(127[12] 300[6])
    defparam i13192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13193_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17302));   // verilog/coms.v(127[12] 300[6])
    defparam i13193_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1400_8 (.CI(n25382), .I0(GND_net), .I1(n1636), .CO(n25383));
    SB_LUT4 add_1400_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1714), .I3(n25381), 
            .O(n4675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13194_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17303));   // verilog/coms.v(127[12] 300[6])
    defparam i13194_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1400_7 (.CI(n25381), .I0(GND_net), .I1(n1714), .CO(n25382));
    SB_LUT4 add_1400_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1792), .I3(n25380), 
            .O(n4676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_6 (.CI(n25380), .I0(GND_net), .I1(n1792), .CO(n25381));
    SB_LUT4 i28529_4_lut (.I0(n752), .I1(n755), .I2(n753), .I3(n4_adj_4640), 
            .O(n778));
    defparam i28529_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 add_1400_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1870), .I3(n25379), 
            .O(n4677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i466_3_lut (.I0(n678), .I1(n731), 
            .I2(n700), .I3(GND_net), .O(n756));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13195_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17304));   // verilog/coms.v(127[12] 300[6])
    defparam i13195_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1400_5 (.CI(n25379), .I0(GND_net), .I1(n1870), .CO(n25380));
    SB_LUT4 i13196_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17305));   // verilog/coms.v(127[12] 300[6])
    defparam i13196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i519_3_lut (.I0(n756), .I1(n809), 
            .I2(n778), .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_i519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13197_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17306));   // verilog/coms.v(127[12] 300[6])
    defparam i13197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1400_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1948), .I3(n25378), 
            .O(n4678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_4 (.CI(n25378), .I0(GND_net), .I1(n1948), .CO(n25379));
    SB_LUT4 add_1400_3_lut (.I0(GND_net), .I1(GND_net), .I2(n2026), .I3(n25377), 
            .O(n4679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_3 (.CI(n25377), .I0(GND_net), .I1(n2026), .CO(n25378));
    SB_LUT4 add_1400_2_lut (.I0(GND_net), .I1(GND_net), .I2(n22055), .I3(VCC_net), 
            .O(n4680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1400_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1400_2 (.CI(VCC_net), .I0(GND_net), .I1(n22055), .CO(n25377));
    SB_LUT4 encoder0_position_23__I_0_add_1308_24_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n25376), .O(n1975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13198_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17307));   // verilog/coms.v(127[12] 300[6])
    defparam i13198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13199_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17308));   // verilog/coms.v(127[12] 300[6])
    defparam i13199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1308_23_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n25375), .O(n1976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13200_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17309));   // verilog/coms.v(127[12] 300[6])
    defparam i13200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13201_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17310));   // verilog/coms.v(127[12] 300[6])
    defparam i13201_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1308_23 (.CI(n25375), .I0(n1923), 
            .I1(VCC_net), .CO(n25376));
    SB_LUT4 i13202_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17311));   // verilog/coms.v(127[12] 300[6])
    defparam i13202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1308_22_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n25374), .O(n1977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_22 (.CI(n25374), .I0(n1924), 
            .I1(VCC_net), .CO(n25375));
    SB_LUT4 encoder0_position_23__I_0_add_1308_21_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n25373), .O(n1978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_21 (.CI(n25373), .I0(n1925), 
            .I1(VCC_net), .CO(n25374));
    SB_LUT4 mux_40_i9_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i13203_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17312));   // verilog/coms.v(127[12] 300[6])
    defparam i13203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13204_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17313));   // verilog/coms.v(127[12] 300[6])
    defparam i13204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1308_20_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n25372), .O(n1979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_20 (.CI(n25372), .I0(n1926), 
            .I1(VCC_net), .CO(n25373));
    SB_LUT4 encoder0_position_23__I_0_add_1308_19_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n25371), .O(n1980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_19 (.CI(n25371), .I0(n1927), 
            .I1(VCC_net), .CO(n25372));
    SB_LUT4 i13205_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17314));   // verilog/coms.v(127[12] 300[6])
    defparam i13205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_40_i10_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[9]), 
            .I3(encoder0_position_scaled[9]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_add_1308_18_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n25370), .O(n1981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13207_4_lut (.I0(n30267), .I1(state[1]), .I2(state_3__N_272[1]), 
            .I3(n16698), .O(n17316));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13207_4_lut.LUT_INIT = 16'hfaee;
    SB_CARRY encoder0_position_23__I_0_add_1308_18 (.CI(n25370), .I0(n1928), 
            .I1(VCC_net), .CO(n25371));
    SB_LUT4 encoder0_position_23__I_0_add_1308_17_lut (.I0(GND_net), .I1(n1929), 
            .I2(VCC_net), .I3(n25369), .O(n1982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_40_i11_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[10]), 
            .I3(encoder0_position_scaled[10]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_23__I_0_add_1308_17 (.CI(n25369), .I0(n1929), 
            .I1(VCC_net), .CO(n25370));
    SB_LUT4 encoder0_position_23__I_0_add_1308_16_lut (.I0(GND_net), .I1(n1930), 
            .I2(VCC_net), .I3(n25368), .O(n1983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_16 (.CI(n25368), .I0(n1930), 
            .I1(VCC_net), .CO(n25369));
    SB_LUT4 i13211_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n4216), .I3(GND_net), .O(n17320));   // verilog/coms.v(127[12] 300[6])
    defparam i13211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1308_15_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n25367), .O(n1984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13212_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n4216), .I3(GND_net), .O(n17321));   // verilog/coms.v(127[12] 300[6])
    defparam i13212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13213_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n4216), .I3(GND_net), .O(n17322));   // verilog/coms.v(127[12] 300[6])
    defparam i13213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13214_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n4216), .I3(GND_net), .O(n17323));   // verilog/coms.v(127[12] 300[6])
    defparam i13214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13215_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n4216), .I3(GND_net), .O(n17324));   // verilog/coms.v(127[12] 300[6])
    defparam i13215_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1308_15 (.CI(n25367), .I0(n1931), 
            .I1(VCC_net), .CO(n25368));
    SB_LUT4 encoder0_position_23__I_0_add_1308_14_lut (.I0(GND_net), .I1(n1932), 
            .I2(VCC_net), .I3(n25366), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_14 (.CI(n25366), .I0(n1932), 
            .I1(VCC_net), .CO(n25367));
    SB_LUT4 encoder0_position_23__I_0_add_1308_13_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n25365), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13216_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n4216), .I3(GND_net), .O(n17325));   // verilog/coms.v(127[12] 300[6])
    defparam i13216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13217_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n4216), .I3(GND_net), .O(n17326));   // verilog/coms.v(127[12] 300[6])
    defparam i13217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13218_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n4216), .I3(GND_net), .O(n17327));   // verilog/coms.v(127[12] 300[6])
    defparam i13218_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1308_13 (.CI(n25365), .I0(n1933), 
            .I1(VCC_net), .CO(n25366));
    SB_LUT4 encoder0_position_23__I_0_add_1308_12_lut (.I0(GND_net), .I1(n1934), 
            .I2(VCC_net), .I3(n25364), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13219_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n4216), .I3(GND_net), .O(n17328));   // verilog/coms.v(127[12] 300[6])
    defparam i13219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13220_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n4216), .I3(GND_net), .O(n17329));   // verilog/coms.v(127[12] 300[6])
    defparam i13220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13221_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n4216), .I3(GND_net), .O(n17330));   // verilog/coms.v(127[12] 300[6])
    defparam i13221_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1308_12 (.CI(n25364), .I0(n1934), 
            .I1(VCC_net), .CO(n25365));
    SB_LUT4 i13222_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n4216), .I3(GND_net), .O(n17331));   // verilog/coms.v(127[12] 300[6])
    defparam i13222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13223_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n4216), .I3(GND_net), .O(n17332));   // verilog/coms.v(127[12] 300[6])
    defparam i13223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13224_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n4216), .I3(GND_net), .O(n17333));   // verilog/coms.v(127[12] 300[6])
    defparam i13224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1308_11_lut (.I0(GND_net), .I1(n1935), 
            .I2(VCC_net), .I3(n25363), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_11 (.CI(n25363), .I0(n1935), 
            .I1(VCC_net), .CO(n25364));
    SB_LUT4 encoder0_position_23__I_0_add_1308_10_lut (.I0(GND_net), .I1(n1936), 
            .I2(VCC_net), .I3(n25362), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_10 (.CI(n25362), .I0(n1936), 
            .I1(VCC_net), .CO(n25363));
    SB_LUT4 encoder0_position_23__I_0_add_1308_9_lut (.I0(GND_net), .I1(n1937), 
            .I2(VCC_net), .I3(n25361), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_40_i12_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[11]), 
            .I3(encoder0_position_scaled[11]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_23__I_0_add_1308_9 (.CI(n25361), .I0(n1937), 
            .I1(VCC_net), .CO(n25362));
    SB_LUT4 i13225_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n4216), .I3(GND_net), .O(n17334));   // verilog/coms.v(127[12] 300[6])
    defparam i13225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13226_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n4216), .I3(GND_net), .O(n17335));   // verilog/coms.v(127[12] 300[6])
    defparam i13226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_40_i13_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[12]), 
            .I3(encoder0_position_scaled[12]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i13227_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n28583), .I3(GND_net), .O(n17336));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13227_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_8_lut (.I0(GND_net), .I1(n1938), 
            .I2(VCC_net), .I3(n25360), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_8 (.CI(n25360), .I0(n1938), 
            .I1(VCC_net), .CO(n25361));
    SB_LUT4 encoder0_position_23__I_0_add_1308_7_lut (.I0(GND_net), .I1(n1939), 
            .I2(GND_net), .I3(n25359), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_7 (.CI(n25359), .I0(n1939), 
            .I1(GND_net), .CO(n25360));
    SB_LUT4 encoder0_position_23__I_0_add_1308_6_lut (.I0(GND_net), .I1(n1940), 
            .I2(GND_net), .I3(n25358), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_6 (.CI(n25358), .I0(n1940), 
            .I1(GND_net), .CO(n25359));
    SB_LUT4 encoder0_position_23__I_0_add_1308_5_lut (.I0(GND_net), .I1(n1941), 
            .I2(VCC_net), .I3(n25357), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_5 (.CI(n25357), .I0(n1941), 
            .I1(VCC_net), .CO(n25358));
    SB_LUT4 encoder0_position_23__I_0_add_1308_4_lut (.I0(GND_net), .I1(n1942), 
            .I2(GND_net), .I3(n25356), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_4591), .I3(n25729), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_4592), .I3(n25728), .O(n3_adj_4527)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_4 (.CI(n25356), .I0(n1942), 
            .I1(GND_net), .CO(n25357));
    SB_LUT4 encoder0_position_23__I_0_add_1308_3_lut (.I0(GND_net), .I1(n1943), 
            .I2(VCC_net), .I3(n25355), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_3 (.CI(n25355), .I0(n1943), 
            .I1(VCC_net), .CO(n25356));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_25 (.CI(n25728), 
            .I0(GND_net), .I1(n3_adj_4592), .CO(n25729));
    SB_LUT4 encoder0_position_23__I_0_add_1308_2_lut (.I0(GND_net), .I1(n444), 
            .I2(GND_net), .I3(VCC_net), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_2 (.CI(VCC_net), .I0(n444), 
            .I1(GND_net), .CO(n25355));
    SB_CARRY add_486_17 (.CI(n24939), .I0(n34501), .I1(n10), .CO(n24940));
    SB_LUT4 encoder0_position_23__I_0_add_1255_23_lut (.I0(GND_net), .I1(n1844), 
            .I2(VCC_net), .I3(n25354), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_486_16_lut (.I0(duty[14]), .I1(n34501), .I2(n11), .I3(n24938), 
            .O(pwm_setpoint_22__N_3[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1255_22_lut (.I0(GND_net), .I1(n1845), 
            .I2(VCC_net), .I3(n25353), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13228_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n28583), .I3(GND_net), .O(n17337));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13228_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13229_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n28583), .I3(GND_net), .O(n17338));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13229_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1255_22 (.CI(n25353), .I0(n1845), 
            .I1(VCC_net), .CO(n25354));
    SB_LUT4 i13230_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n28583), .I3(GND_net), .O(n17339));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13230_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1255_21_lut (.I0(GND_net), .I1(n1846), 
            .I2(VCC_net), .I3(n25352), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_4593), .I3(n25727), .O(n4_adj_4526)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13231_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n28583), .I3(GND_net), .O(n17340));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13231_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4610));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_24 (.CI(n25727), 
            .I0(GND_net), .I1(n4_adj_4593), .CO(n25728));
    SB_CARRY encoder0_position_23__I_0_add_1255_21 (.CI(n25352), .I0(n1846), 
            .I1(VCC_net), .CO(n25353));
    SB_LUT4 encoder0_position_23__I_0_add_1255_20_lut (.I0(GND_net), .I1(n1847), 
            .I2(VCC_net), .I3(n25351), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_486_16 (.CI(n24938), .I0(n34501), .I1(n11), .CO(n24939));
    SB_CARRY encoder0_position_23__I_0_add_1255_20 (.CI(n25351), .I0(n1847), 
            .I1(VCC_net), .CO(n25352));
    SB_LUT4 encoder0_position_23__I_0_add_1255_19_lut (.I0(GND_net), .I1(n1848), 
            .I2(VCC_net), .I3(n25350), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_19 (.CI(n25350), .I0(n1848), 
            .I1(VCC_net), .CO(n25351));
    SB_LUT4 encoder0_position_23__I_0_add_1255_18_lut (.I0(GND_net), .I1(n1849), 
            .I2(VCC_net), .I3(n25349), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_18 (.CI(n25349), .I0(n1849), 
            .I1(VCC_net), .CO(n25350));
    SB_LUT4 encoder0_position_23__I_0_add_1255_17_lut (.I0(GND_net), .I1(n1850), 
            .I2(VCC_net), .I3(n25348), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_17 (.CI(n25348), .I0(n1850), 
            .I1(VCC_net), .CO(n25349));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_4594), .I3(n25726), .O(n5_adj_4525)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13232_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n28583), .I3(GND_net), .O(n17341));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13232_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_40_i14_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[13]), 
            .I3(encoder0_position_scaled[13]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_add_1255_16_lut (.I0(GND_net), .I1(n1851), 
            .I2(VCC_net), .I3(n25347), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_16 (.CI(n25347), .I0(n1851), 
            .I1(VCC_net), .CO(n25348));
    SB_LUT4 add_486_15_lut (.I0(duty[13]), .I1(n34501), .I2(n12), .I3(n24937), 
            .O(pwm_setpoint_22__N_3[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1255_15_lut (.I0(GND_net), .I1(n1852), 
            .I2(VCC_net), .I3(n25346), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_15 (.CI(n25346), .I0(n1852), 
            .I1(VCC_net), .CO(n25347));
    SB_LUT4 encoder0_position_23__I_0_add_1255_14_lut (.I0(GND_net), .I1(n1853), 
            .I2(VCC_net), .I3(n25345), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_14 (.CI(n25345), .I0(n1853), 
            .I1(VCC_net), .CO(n25346));
    SB_LUT4 encoder0_position_23__I_0_add_1255_13_lut (.I0(GND_net), .I1(n1854), 
            .I2(VCC_net), .I3(n25344), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_23 (.CI(n25726), 
            .I0(GND_net), .I1(n5_adj_4594), .CO(n25727));
    SB_CARRY encoder0_position_23__I_0_add_1255_13 (.CI(n25344), .I0(n1854), 
            .I1(VCC_net), .CO(n25345));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_4595), .I3(n25725), .O(n6_adj_4524)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_22 (.CI(n25725), 
            .I0(GND_net), .I1(n6_adj_4595), .CO(n25726));
    SB_LUT4 i13233_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n28583), .I3(GND_net), .O(n17342));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13233_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1255_12_lut (.I0(GND_net), .I1(n1855), 
            .I2(VCC_net), .I3(n25343), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_4596), .I3(n25724), .O(n7_adj_4523)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13234_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n28583), .I3(GND_net), .O(n17343));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13234_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_21 (.CI(n25724), 
            .I0(GND_net), .I1(n7_adj_4596), .CO(n25725));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_4597), .I3(n25723), .O(n8_adj_4522)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_12 (.CI(n25343), .I0(n1855), 
            .I1(VCC_net), .CO(n25344));
    SB_LUT4 encoder0_position_23__I_0_add_1255_11_lut (.I0(GND_net), .I1(n1856), 
            .I2(VCC_net), .I3(n25342), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_11 (.CI(n25342), .I0(n1856), 
            .I1(VCC_net), .CO(n25343));
    SB_LUT4 i13235_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n28583), .I3(GND_net), .O(n17344));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13235_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_486_15 (.CI(n24937), .I0(n34501), .I1(n12), .CO(n24938));
    SB_LUT4 encoder0_position_23__I_0_add_1255_10_lut (.I0(GND_net), .I1(n1857), 
            .I2(VCC_net), .I3(n25341), .O(n1910)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_10 (.CI(n25341), .I0(n1857), 
            .I1(VCC_net), .CO(n25342));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_20 (.CI(n25723), 
            .I0(GND_net), .I1(n8_adj_4597), .CO(n25724));
    SB_LUT4 add_486_14_lut (.I0(duty[12]), .I1(n34501), .I2(n13), .I3(n24936), 
            .O(pwm_setpoint_22__N_3[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1255_9_lut (.I0(GND_net), .I1(n1858), 
            .I2(VCC_net), .I3(n25340), .O(n1911)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13236_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n28583), .I3(GND_net), .O(n17345));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13236_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_486_14 (.CI(n24936), .I0(n34501), .I1(n13), .CO(n24937));
    SB_CARRY encoder0_position_23__I_0_add_1255_9 (.CI(n25340), .I0(n1858), 
            .I1(VCC_net), .CO(n25341));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_4598), .I3(n25722), .O(n9_adj_4521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_19 (.CI(n25722), 
            .I0(GND_net), .I1(n9_adj_4598), .CO(n25723));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_4599), .I3(n25721), .O(n10_adj_4520)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_8_lut (.I0(GND_net), .I1(n1859), 
            .I2(VCC_net), .I3(n25339), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_486_13_lut (.I0(duty[11]), .I1(n34501), .I2(n14), .I3(n24935), 
            .O(pwm_setpoint_22__N_3[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_18 (.CI(n25721), 
            .I0(GND_net), .I1(n10_adj_4599), .CO(n25722));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_4600), .I3(n25720), .O(n11_adj_4519)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_8 (.CI(n25339), .I0(n1859), 
            .I1(VCC_net), .CO(n25340));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_17 (.CI(n25720), 
            .I0(GND_net), .I1(n11_adj_4600), .CO(n25721));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_4601), .I3(n25719), .O(n12_adj_4518)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_7_lut (.I0(GND_net), .I1(n1860), 
            .I2(GND_net), .I3(n25338), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_16 (.CI(n25719), 
            .I0(GND_net), .I1(n12_adj_4601), .CO(n25720));
    SB_CARRY add_486_13 (.CI(n24935), .I0(n34501), .I1(n14), .CO(n24936));
    SB_LUT4 i13237_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n28583), .I3(GND_net), .O(n17346));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13237_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1255_7 (.CI(n25338), .I0(n1860), 
            .I1(GND_net), .CO(n25339));
    SB_LUT4 encoder0_position_23__I_0_add_1255_6_lut (.I0(GND_net), .I1(n1861), 
            .I2(GND_net), .I3(n25337), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_6 (.CI(n25337), .I0(n1861), 
            .I1(GND_net), .CO(n25338));
    SB_LUT4 encoder0_position_23__I_0_add_1255_5_lut (.I0(GND_net), .I1(n1862), 
            .I2(VCC_net), .I3(n25336), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_5 (.CI(n25336), .I0(n1862), 
            .I1(VCC_net), .CO(n25337));
    SB_LUT4 add_486_12_lut (.I0(duty[10]), .I1(n34501), .I2(n15), .I3(n24934), 
            .O(pwm_setpoint_22__N_3[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_4602), .I3(n25718), .O(n13_adj_4517)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_4_lut (.I0(GND_net), .I1(n1863), 
            .I2(GND_net), .I3(n25335), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_486_12 (.CI(n24934), .I0(n34501), .I1(n15), .CO(n24935));
    SB_CARRY encoder0_position_23__I_0_add_1255_4 (.CI(n25335), .I0(n1863), 
            .I1(GND_net), .CO(n25336));
    SB_LUT4 encoder0_position_23__I_0_add_1255_3_lut (.I0(GND_net), .I1(n1864), 
            .I2(VCC_net), .I3(n25334), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_3 (.CI(n25334), .I0(n1864), 
            .I1(VCC_net), .CO(n25335));
    SB_LUT4 encoder0_position_23__I_0_add_1255_2_lut (.I0(GND_net), .I1(n443), 
            .I2(GND_net), .I3(VCC_net), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_2 (.CI(VCC_net), .I0(n443), 
            .I1(GND_net), .CO(n25334));
    SB_LUT4 encoder0_position_23__I_0_add_1202_22_lut (.I0(GND_net), .I1(n1766), 
            .I2(VCC_net), .I3(n25333), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_486_11_lut (.I0(duty[9]), .I1(n34501), .I2(n16), .I3(n24933), 
            .O(pwm_setpoint_22__N_3[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_486_11 (.CI(n24933), .I0(n34501), .I1(n16), .CO(n24934));
    SB_LUT4 add_486_10_lut (.I0(duty[8]), .I1(n34501), .I2(n17), .I3(n24932), 
            .O(pwm_setpoint_22__N_3[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1202_21_lut (.I0(GND_net), .I1(n1767), 
            .I2(VCC_net), .I3(n25332), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_21 (.CI(n25332), .I0(n1767), 
            .I1(VCC_net), .CO(n25333));
    SB_LUT4 i13238_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n28583), .I3(GND_net), .O(n17347));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13238_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_15 (.CI(n25718), 
            .I0(GND_net), .I1(n13_adj_4602), .CO(n25719));
    SB_LUT4 encoder0_position_23__I_0_add_1202_20_lut (.I0(GND_net), .I1(n1768), 
            .I2(VCC_net), .I3(n25331), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_486_10 (.CI(n24932), .I0(n34501), .I1(n17), .CO(n24933));
    SB_LUT4 i13239_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n28583), .I3(GND_net), .O(n17348));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_40_i15_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[14]), 
            .I3(encoder0_position_scaled[14]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i13240_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n28583), .I3(GND_net), .O(n17349));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13240_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1202_20 (.CI(n25331), .I0(n1768), 
            .I1(VCC_net), .CO(n25332));
    SB_LUT4 encoder0_position_23__I_0_add_1202_19_lut (.I0(GND_net), .I1(n1769), 
            .I2(VCC_net), .I3(n25330), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13241_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n28583), .I3(GND_net), .O(n17350));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28429_2_lut_3_lut (.I0(n3_adj_4527), .I1(n4_adj_4625), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n619));
    defparam i28429_2_lut_3_lut.LUT_INIT = 16'h7f7f;
    SB_CARRY encoder0_position_23__I_0_add_1202_19 (.CI(n25330), .I0(n1769), 
            .I1(VCC_net), .CO(n25331));
    SB_LUT4 encoder0_position_23__I_0_add_1202_18_lut (.I0(GND_net), .I1(n1770), 
            .I2(VCC_net), .I3(n25329), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_18 (.CI(n25329), .I0(n1770), 
            .I1(VCC_net), .CO(n25330));
    SB_LUT4 i24629_3_lut_4_lut (.I0(n3_adj_4527), .I1(n4_adj_4625), .I2(n4431), 
            .I3(n4_adj_4526), .O(n30290));
    defparam i24629_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_23__I_0_add_1202_17_lut (.I0(GND_net), .I1(n1771), 
            .I2(VCC_net), .I3(n25328), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24623_3_lut_4_lut (.I0(n3_adj_4527), .I1(n4_adj_4625), .I2(n4434), 
            .I3(n7_adj_4523), .O(n30284));
    defparam i24623_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13242_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n28583), .I3(GND_net), .O(n17351));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24625_3_lut_4_lut (.I0(n3_adj_4527), .I1(n4_adj_4625), .I2(n4433), 
            .I3(n6_adj_4524), .O(n30286));
    defparam i24625_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i24627_3_lut_4_lut (.I0(n3_adj_4527), .I1(n4_adj_4625), .I2(n4432), 
            .I3(n5_adj_4525), .O(n30288));
    defparam i24627_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY encoder0_position_23__I_0_add_1202_17 (.CI(n25328), .I0(n1771), 
            .I1(VCC_net), .CO(n25329));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_4603), .I3(n25717), .O(n14_adj_4516)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13243_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n28583), .I3(GND_net), .O(n17352));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13244_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n28583), .I3(GND_net), .O(n17353));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1202_16_lut (.I0(GND_net), .I1(n1772), 
            .I2(VCC_net), .I3(n25327), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_16 (.CI(n25327), .I0(n1772), 
            .I1(VCC_net), .CO(n25328));
    SB_LUT4 add_486_9_lut (.I0(duty[7]), .I1(n34501), .I2(n18), .I3(n24931), 
            .O(pwm_setpoint_22__N_3[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_486_9 (.CI(n24931), .I0(n34501), .I1(n18), .CO(n24932));
    SB_LUT4 encoder0_position_23__I_0_add_1202_15_lut (.I0(GND_net), .I1(n1773), 
            .I2(VCC_net), .I3(n25326), .O(n1826)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_15 (.CI(n25326), .I0(n1773), 
            .I1(VCC_net), .CO(n25327));
    SB_LUT4 add_486_8_lut (.I0(duty[6]), .I1(n34501), .I2(n19), .I3(n24930), 
            .O(pwm_setpoint_22__N_3[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_486_8 (.CI(n24930), .I0(n34501), .I1(n19), .CO(n24931));
    SB_LUT4 mux_40_i16_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[15]), 
            .I3(encoder0_position_scaled[15]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_14 (.CI(n25717), 
            .I0(GND_net), .I1(n14_adj_4603), .CO(n25718));
    SB_LUT4 encoder0_position_23__I_0_add_1202_14_lut (.I0(GND_net), .I1(n1774), 
            .I2(VCC_net), .I3(n25325), .O(n1827)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_486_7_lut (.I0(duty[5]), .I1(n34501), .I2(n20), .I3(n24929), 
            .O(pwm_setpoint_22__N_3[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_486_7 (.CI(n24929), .I0(n34501), .I1(n20), .CO(n24930));
    SB_CARRY encoder0_position_23__I_0_add_1202_14 (.CI(n25325), .I0(n1774), 
            .I1(VCC_net), .CO(n25326));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_4604), .I3(n25716), .O(n15_adj_4515)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_486_6_lut (.I0(duty[4]), .I1(n34501), .I2(n21), .I3(n24928), 
            .O(pwm_setpoint_22__N_3[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_13 (.CI(n25716), 
            .I0(GND_net), .I1(n15_adj_4604), .CO(n25717));
    SB_CARRY add_486_6 (.CI(n24928), .I0(n34501), .I1(n21), .CO(n24929));
    SB_LUT4 encoder0_position_23__I_0_add_1202_13_lut (.I0(GND_net), .I1(n1775), 
            .I2(VCC_net), .I3(n25324), .O(n1828)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13245_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n28583), .I3(GND_net), .O(n17354));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13245_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1202_13 (.CI(n25324), .I0(n1775), 
            .I1(VCC_net), .CO(n25325));
    SB_LUT4 encoder0_position_23__I_0_add_1202_12_lut (.I0(GND_net), .I1(n1776), 
            .I2(VCC_net), .I3(n25323), .O(n1829)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13246_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n28583), .I3(GND_net), .O(n17355));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13246_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1202_12 (.CI(n25323), .I0(n1776), 
            .I1(VCC_net), .CO(n25324));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_4605), .I3(n25715), .O(n16_adj_4514)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1202_11_lut (.I0(GND_net), .I1(n1777), 
            .I2(VCC_net), .I3(n25322), .O(n1830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_11 (.CI(n25322), .I0(n1777), 
            .I1(VCC_net), .CO(n25323));
    SB_LUT4 encoder0_position_23__I_0_add_1202_10_lut (.I0(GND_net), .I1(n1778), 
            .I2(VCC_net), .I3(n25321), .O(n1831)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_10 (.CI(n25321), .I0(n1778), 
            .I1(VCC_net), .CO(n25322));
    SB_LUT4 encoder0_position_23__I_0_add_1202_9_lut (.I0(GND_net), .I1(n1779), 
            .I2(VCC_net), .I3(n25320), .O(n1832)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_9 (.CI(n25320), .I0(n1779), 
            .I1(VCC_net), .CO(n25321));
    SB_LUT4 encoder0_position_23__I_0_add_1202_8_lut (.I0(GND_net), .I1(n1780), 
            .I2(VCC_net), .I3(n25319), .O(n1833)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_8 (.CI(n25319), .I0(n1780), 
            .I1(VCC_net), .CO(n25320));
    SB_LUT4 encoder0_position_23__I_0_add_1202_7_lut (.I0(GND_net), .I1(n1781), 
            .I2(GND_net), .I3(n25318), .O(n1834)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_7 (.CI(n25318), .I0(n1781), 
            .I1(GND_net), .CO(n25319));
    SB_LUT4 encoder0_position_23__I_0_add_1202_6_lut (.I0(GND_net), .I1(n1782), 
            .I2(GND_net), .I3(n25317), .O(n1835)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_6 (.CI(n25317), .I0(n1782), 
            .I1(GND_net), .CO(n25318));
    SB_LUT4 encoder0_position_23__I_0_add_1202_5_lut (.I0(GND_net), .I1(n1783), 
            .I2(VCC_net), .I3(n25316), .O(n1836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_5 (.CI(n25316), .I0(n1783), 
            .I1(VCC_net), .CO(n25317));
    SB_LUT4 mux_40_i17_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[16]), 
            .I3(encoder0_position_scaled[16]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i13247_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n28583), .I3(GND_net), .O(n17356));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13248_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n28583), .I3(GND_net), .O(n17357));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13248_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_12 (.CI(n25715), 
            .I0(GND_net), .I1(n16_adj_4605), .CO(n25716));
    SB_LUT4 encoder0_position_23__I_0_add_1202_4_lut (.I0(GND_net), .I1(n1784), 
            .I2(GND_net), .I3(n25315), .O(n1837)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_486_5_lut (.I0(duty[3]), .I1(n34501), .I2(n22), .I3(n24927), 
            .O(pwm_setpoint_22__N_3[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_1202_4 (.CI(n25315), .I0(n1784), 
            .I1(GND_net), .CO(n25316));
    SB_LUT4 encoder0_position_23__I_0_add_1202_3_lut (.I0(GND_net), .I1(n1785), 
            .I2(VCC_net), .I3(n25314), .O(n1838)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_3 (.CI(n25314), .I0(n1785), 
            .I1(VCC_net), .CO(n25315));
    SB_LUT4 encoder0_position_23__I_0_add_1202_2_lut (.I0(GND_net), .I1(n442), 
            .I2(GND_net), .I3(VCC_net), .O(n1839)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_4606), .I3(n25714), .O(n17_adj_4513)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_2 (.CI(VCC_net), .I0(n442), 
            .I1(GND_net), .CO(n25314));
    SB_CARRY add_486_5 (.CI(n24927), .I0(n34501), .I1(n22), .CO(n24928));
    SB_LUT4 add_486_4_lut (.I0(duty[2]), .I1(n34501), .I2(n23), .I3(n24926), 
            .O(pwm_setpoint_22__N_3[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_11 (.CI(n25714), 
            .I0(GND_net), .I1(n17_adj_4606), .CO(n25715));
    SB_LUT4 encoder0_position_23__I_0_add_1149_21_lut (.I0(GND_net), .I1(n1688), 
            .I2(VCC_net), .I3(n25313), .O(n1741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13249_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n28583), .I3(GND_net), .O(n17358));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13250_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n28583), .I3(GND_net), .O(n17359));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1149_20_lut (.I0(GND_net), .I1(n1689), 
            .I2(VCC_net), .I3(n25312), .O(n1742)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_20 (.CI(n25312), .I0(n1689), 
            .I1(VCC_net), .CO(n25313));
    SB_LUT4 encoder0_position_23__I_0_add_1149_19_lut (.I0(GND_net), .I1(n1690), 
            .I2(VCC_net), .I3(n25311), .O(n1743)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13251_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n28583), .I3(GND_net), .O(n17360));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13251_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1149_19 (.CI(n25311), .I0(n1690), 
            .I1(VCC_net), .CO(n25312));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_4607), .I3(n25713), .O(n18_adj_4512)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1149_18_lut (.I0(GND_net), .I1(n1691), 
            .I2(VCC_net), .I3(n25310), .O(n1744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_18 (.CI(n25310), .I0(n1691), 
            .I1(VCC_net), .CO(n25311));
    SB_LUT4 encoder0_position_23__I_0_add_1149_17_lut (.I0(GND_net), .I1(n1692), 
            .I2(VCC_net), .I3(n25309), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_10 (.CI(n25713), 
            .I0(GND_net), .I1(n18_adj_4607), .CO(n25714));
    SB_CARRY encoder0_position_23__I_0_add_1149_17 (.CI(n25309), .I0(n1692), 
            .I1(VCC_net), .CO(n25310));
    SB_LUT4 encoder0_position_23__I_0_add_1149_16_lut (.I0(GND_net), .I1(n1693), 
            .I2(VCC_net), .I3(n25308), .O(n1746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_16 (.CI(n25308), .I0(n1693), 
            .I1(VCC_net), .CO(n25309));
    SB_LUT4 encoder0_position_23__I_0_add_1149_15_lut (.I0(GND_net), .I1(n1694), 
            .I2(VCC_net), .I3(n25307), .O(n1747)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_15 (.CI(n25307), .I0(n1694), 
            .I1(VCC_net), .CO(n25308));
    SB_LUT4 encoder0_position_23__I_0_add_1149_14_lut (.I0(GND_net), .I1(n1695), 
            .I2(VCC_net), .I3(n25306), .O(n1748)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_14 (.CI(n25306), .I0(n1695), 
            .I1(VCC_net), .CO(n25307));
    SB_LUT4 encoder0_position_23__I_0_add_1149_13_lut (.I0(GND_net), .I1(n1696), 
            .I2(VCC_net), .I3(n25305), .O(n1749)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_13 (.CI(n25305), .I0(n1696), 
            .I1(VCC_net), .CO(n25306));
    SB_LUT4 i13252_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n28583), .I3(GND_net), .O(n17361));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1149_12_lut (.I0(GND_net), .I1(n1697), 
            .I2(VCC_net), .I3(n25304), .O(n1750)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_12 (.CI(n25304), .I0(n1697), 
            .I1(VCC_net), .CO(n25305));
    SB_LUT4 encoder0_position_23__I_0_add_1149_11_lut (.I0(GND_net), .I1(n1698), 
            .I2(VCC_net), .I3(n25303), .O(n1751)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_11 (.CI(n25303), .I0(n1698), 
            .I1(VCC_net), .CO(n25304));
    SB_LUT4 encoder0_position_23__I_0_add_1149_10_lut (.I0(GND_net), .I1(n1699), 
            .I2(VCC_net), .I3(n25302), .O(n1752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_10 (.CI(n25302), .I0(n1699), 
            .I1(VCC_net), .CO(n25303));
    SB_LUT4 encoder0_position_23__I_0_add_1149_9_lut (.I0(GND_net), .I1(n1700), 
            .I2(VCC_net), .I3(n25301), .O(n1753)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_9 (.CI(n25301), .I0(n1700), 
            .I1(VCC_net), .CO(n25302));
    SB_LUT4 i13253_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n28583), .I3(GND_net), .O(n17362));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13254_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n28583), .I3(GND_net), .O(n17363));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13254_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13255_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n28583), .I3(GND_net), .O(n17364));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13255_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13256_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n28583), .I3(GND_net), .O(n17365));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13256_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i409_3_lut_4_lut (.I0(n2), .I1(encoder0_position[23]), 
            .I2(n619), .I3(n4429), .O(n674));
    defparam encoder0_position_23__I_0_i409_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_LUT4 i13257_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n28583), .I3(GND_net), .O(n17366));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13258_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n4216), .I3(GND_net), .O(n17367));   // verilog/coms.v(127[12] 300[6])
    defparam i13258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13259_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n4216), .I3(GND_net), .O(n17368));   // verilog/coms.v(127[12] 300[6])
    defparam i13259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13260_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n4216), .I3(GND_net), .O(n17369));   // verilog/coms.v(127[12] 300[6])
    defparam i13260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13261_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n4216), .I3(GND_net), .O(n17370));   // verilog/coms.v(127[12] 300[6])
    defparam i13261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13262_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n4216), .I3(GND_net), .O(n17371));   // verilog/coms.v(127[12] 300[6])
    defparam i13262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13263_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n4216), .I3(GND_net), .O(n17372));   // verilog/coms.v(127[12] 300[6])
    defparam i13263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13264_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n4216), .I3(GND_net), .O(n17373));   // verilog/coms.v(127[12] 300[6])
    defparam i13264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13271_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4530), 
            .I3(n15590), .O(n17380));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13271_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13272_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n31883), 
            .I3(GND_net), .O(n17381));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13273_3_lut (.I0(quadA_debounced_adj_4504), .I1(reg_B_adj_4715[1]), 
            .I2(n32056), .I3(GND_net), .O(n17382));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_40_i18_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[17]), 
            .I3(encoder0_position_scaled[17]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i13267_3_lut (.I0(n16802), .I1(r_Bit_Index[0]), .I2(n16710), 
            .I3(GND_net), .O(n17376));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13267_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4609));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1149_8_lut (.I0(GND_net), .I1(n1701), 
            .I2(VCC_net), .I3(n25300), .O(n1754)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_8 (.CI(n25300), .I0(n1701), 
            .I1(VCC_net), .CO(n25301));
    SB_LUT4 encoder0_position_23__I_0_add_1149_7_lut (.I0(GND_net), .I1(n1702), 
            .I2(GND_net), .I3(n25299), .O(n1755)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_7 (.CI(n25299), .I0(n1702), 
            .I1(GND_net), .CO(n25300));
    SB_LUT4 encoder0_position_23__I_0_add_1149_6_lut (.I0(GND_net), .I1(n1703), 
            .I2(GND_net), .I3(n25298), .O(n1756)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_6 (.CI(n25298), .I0(n1703), 
            .I1(GND_net), .CO(n25299));
    SB_LUT4 encoder0_position_23__I_0_add_1149_5_lut (.I0(GND_net), .I1(n1704), 
            .I2(VCC_net), .I3(n25297), .O(n1757)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_5 (.CI(n25297), .I0(n1704), 
            .I1(VCC_net), .CO(n25298));
    SB_LUT4 encoder0_position_23__I_0_add_1149_4_lut (.I0(GND_net), .I1(n1705), 
            .I2(GND_net), .I3(n25296), .O(n1758)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_4 (.CI(n25296), .I0(n1705), 
            .I1(GND_net), .CO(n25297));
    SB_LUT4 encoder0_position_23__I_0_add_1149_3_lut (.I0(GND_net), .I1(n1706), 
            .I2(VCC_net), .I3(n25295), .O(n1759)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_3 (.CI(n25295), .I0(n1706), 
            .I1(VCC_net), .CO(n25296));
    SB_LUT4 encoder0_position_23__I_0_add_1149_2_lut (.I0(GND_net), .I1(n441), 
            .I2(GND_net), .I3(VCC_net), .O(n1760)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_2 (.CI(VCC_net), .I0(n441), 
            .I1(GND_net), .CO(n25295));
    SB_LUT4 encoder0_position_23__I_0_add_1096_20_lut (.I0(GND_net), .I1(n1610), 
            .I2(VCC_net), .I3(n25294), .O(n1663)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_19_lut (.I0(GND_net), .I1(n1611), 
            .I2(VCC_net), .I3(n25293), .O(n1664)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_19 (.CI(n25293), .I0(n1611), 
            .I1(VCC_net), .CO(n25294));
    SB_LUT4 encoder0_position_23__I_0_add_1096_18_lut (.I0(GND_net), .I1(n1612), 
            .I2(VCC_net), .I3(n25292), .O(n1665)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_18 (.CI(n25292), .I0(n1612), 
            .I1(VCC_net), .CO(n25293));
    SB_LUT4 encoder0_position_23__I_0_add_1096_17_lut (.I0(GND_net), .I1(n1613), 
            .I2(VCC_net), .I3(n25291), .O(n1666)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_17 (.CI(n25291), .I0(n1613), 
            .I1(VCC_net), .CO(n25292));
    SB_LUT4 encoder0_position_23__I_0_add_1096_16_lut (.I0(GND_net), .I1(n1614), 
            .I2(VCC_net), .I3(n25290), .O(n1667)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_16 (.CI(n25290), .I0(n1614), 
            .I1(VCC_net), .CO(n25291));
    SB_LUT4 encoder0_position_23__I_0_add_1096_15_lut (.I0(GND_net), .I1(n1615), 
            .I2(VCC_net), .I3(n25289), .O(n1668)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_15 (.CI(n25289), .I0(n1615), 
            .I1(VCC_net), .CO(n25290));
    SB_LUT4 encoder0_position_23__I_0_add_1096_14_lut (.I0(GND_net), .I1(n1616), 
            .I2(VCC_net), .I3(n25288), .O(n1669)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_14 (.CI(n25288), .I0(n1616), 
            .I1(VCC_net), .CO(n25289));
    SB_LUT4 encoder0_position_23__I_0_add_1096_13_lut (.I0(GND_net), .I1(n1617), 
            .I2(VCC_net), .I3(n25287), .O(n1670)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_13 (.CI(n25287), .I0(n1617), 
            .I1(VCC_net), .CO(n25288));
    SB_LUT4 encoder0_position_23__I_0_add_1096_12_lut (.I0(GND_net), .I1(n1618), 
            .I2(VCC_net), .I3(n25286), .O(n1671)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_12 (.CI(n25286), .I0(n1618), 
            .I1(VCC_net), .CO(n25287));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_4608), .I3(n25712), .O(n19_adj_4511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_11_lut (.I0(GND_net), .I1(n1619), 
            .I2(VCC_net), .I3(n25285), .O(n1672)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_11 (.CI(n25285), .I0(n1619), 
            .I1(VCC_net), .CO(n25286));
    SB_LUT4 encoder0_position_23__I_0_add_1096_10_lut (.I0(GND_net), .I1(n1620), 
            .I2(VCC_net), .I3(n25284), .O(n1673)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_10 (.CI(n25284), .I0(n1620), 
            .I1(VCC_net), .CO(n25285));
    SB_LUT4 encoder0_position_23__I_0_add_1096_9_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n25283), .O(n1674)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_9 (.CI(n25283), .I0(n1621), 
            .I1(VCC_net), .CO(n25284));
    SB_LUT4 encoder0_position_23__I_0_add_1096_8_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n25282), .O(n1675)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_8 (.CI(n25282), .I0(n1622), 
            .I1(VCC_net), .CO(n25283));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_9 (.CI(n25712), 
            .I0(GND_net), .I1(n19_adj_4608), .CO(n25713));
    SB_LUT4 encoder0_position_23__I_0_add_1096_7_lut (.I0(GND_net), .I1(n1623), 
            .I2(GND_net), .I3(n25281), .O(n1676)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_7 (.CI(n25281), .I0(n1623), 
            .I1(GND_net), .CO(n25282));
    SB_LUT4 encoder0_position_23__I_0_add_1096_6_lut (.I0(GND_net), .I1(n1624), 
            .I2(GND_net), .I3(n25280), .O(n1677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_6 (.CI(n25280), .I0(n1624), 
            .I1(GND_net), .CO(n25281));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_4609), .I3(n25711), .O(n20_adj_4510)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_5_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n25279), .O(n1678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_5 (.CI(n25279), .I0(n1625), 
            .I1(VCC_net), .CO(n25280));
    SB_LUT4 mux_40_i19_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[18]), 
            .I3(encoder0_position_scaled[18]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_add_1096_4_lut (.I0(GND_net), .I1(n1626), 
            .I2(GND_net), .I3(n25278), .O(n1679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_4 (.CI(n25278), .I0(n1626), 
            .I1(GND_net), .CO(n25279));
    SB_LUT4 mux_40_i20_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[19]), 
            .I3(encoder0_position_scaled[19]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_add_1096_3_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n25277), .O(n1680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_3 (.CI(n25277), .I0(n1627), 
            .I1(VCC_net), .CO(n25278));
    SB_LUT4 encoder0_position_23__I_0_add_1096_2_lut (.I0(GND_net), .I1(n440), 
            .I2(GND_net), .I3(VCC_net), .O(n1681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_2 (.CI(VCC_net), .I0(n440), 
            .I1(GND_net), .CO(n25277));
    SB_LUT4 encoder0_position_23__I_0_add_1043_19_lut (.I0(GND_net), .I1(n1532), 
            .I2(VCC_net), .I3(n25276), .O(n1585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_8 (.CI(n25711), 
            .I0(GND_net), .I1(n20_adj_4609), .CO(n25712));
    SB_LUT4 encoder0_position_23__I_0_add_1043_18_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n25275), .O(n1586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_18 (.CI(n25275), .I0(n1533), 
            .I1(VCC_net), .CO(n25276));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_4610), .I3(n25710), .O(n21_adj_4509)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1043_17_lut (.I0(GND_net), .I1(n1534), 
            .I2(VCC_net), .I3(n25274), .O(n1587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_17 (.CI(n25274), .I0(n1534), 
            .I1(VCC_net), .CO(n25275));
    SB_LUT4 mux_40_i21_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[20]), 
            .I3(encoder0_position_scaled[20]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_40_i22_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[21]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_40_i23_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[22]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4608));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_7 (.CI(n25710), 
            .I0(GND_net), .I1(n21_adj_4610), .CO(n25711));
    SB_LUT4 encoder0_position_23__I_0_add_1043_16_lut (.I0(GND_net), .I1(n1535), 
            .I2(VCC_net), .I3(n25273), .O(n1588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27821_4_lut (.I0(state[0]), .I1(start), .I2(n21971), .I3(\neo_pixel_transmitter.done ), 
            .O(n33118));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27821_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 i27773_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n33120));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27773_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i18_4_lut (.I0(n33120), .I1(n33118), .I2(state[1]), .I3(n22115), 
            .O(n28495));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i12758_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4216), .I3(GND_net), .O(n16867));   // verilog/coms.v(127[12] 300[6])
    defparam i12758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1675 (.I0(\FRAME_MATCHER.i_31__N_2364 ), .I1(n6_adj_4624), 
            .I2(n29497), .I3(n771), .O(n31065));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1675.LUT_INIT = 16'hfcfe;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n63), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n31065), .I3(n12869), .O(n28937));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'hd5f5;
    SB_LUT4 i12761_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n31883), 
            .I3(GND_net), .O(n16870));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12761_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12762_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_4704[1]), .I2(n8947), 
            .I3(n4_adj_4494), .O(n16871));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12762_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i12763_3_lut (.I0(quadB_debounced_adj_4505), .I1(reg_B_adj_4715[0]), 
            .I2(n32056), .I3(GND_net), .O(n16872));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12763_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1677 (.I0(n5_adj_4590), .I1(n122), .I2(n2329), 
            .I3(n63_adj_4566), .O(n6_adj_4656));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1677.LUT_INIT = 16'heaaa;
    SB_LUT4 mux_40_i24_3_lut_4_lut (.I0(n15450), .I1(control_mode[1]), .I2(motor_state_23__N_74[23]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam mux_40_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_23__I_0_add_1043_16 (.CI(n25273), .I0(n1535), 
            .I1(VCC_net), .CO(n25274));
    SB_LUT4 encoder0_position_23__I_0_add_1043_15_lut (.I0(GND_net), .I1(n1536), 
            .I2(VCC_net), .I3(n25272), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_15 (.CI(n25272), .I0(n1536), 
            .I1(VCC_net), .CO(n25273));
    SB_LUT4 i3_4_lut_adj_1678 (.I0(n35368), .I1(n6_adj_4656), .I2(\FRAME_MATCHER.i_31__N_2370 ), 
            .I3(n4452), .O(n8_adj_4489));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1678.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut_adj_1679 (.I0(n122), .I1(n8_adj_4489), .I2(n63), 
            .I3(n5_adj_4639), .O(n35073));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1679.LUT_INIT = 16'hefcf;
    SB_LUT4 encoder0_position_23__I_0_add_1043_14_lut (.I0(GND_net), .I1(n1537), 
            .I2(VCC_net), .I3(n25271), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_14 (.CI(n25271), .I0(n1537), 
            .I1(VCC_net), .CO(n25272));
    SB_LUT4 encoder0_position_23__I_0_add_1043_13_lut (.I0(GND_net), .I1(n1538), 
            .I2(VCC_net), .I3(n25270), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_13 (.CI(n25270), .I0(n1538), 
            .I1(VCC_net), .CO(n25271));
    SB_LUT4 i12765_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n4216), .I3(GND_net), .O(n16874));   // verilog/coms.v(127[12] 300[6])
    defparam i12765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_12_lut (.I0(GND_net), .I1(n1539), 
            .I2(VCC_net), .I3(n25269), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_12 (.CI(n25269), .I0(n1539), 
            .I1(VCC_net), .CO(n25270));
    SB_LUT4 encoder0_position_23__I_0_add_1043_11_lut (.I0(GND_net), .I1(n1540), 
            .I2(VCC_net), .I3(n25268), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1680 (.I0(n15453), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n15455));
    defparam i1_2_lut_adj_1680.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_23__I_0_add_1043_11 (.CI(n25268), .I0(n1540), 
            .I1(VCC_net), .CO(n25269));
    SB_LUT4 i27565_4_lut (.I0(n27), .I1(n15_adj_4576), .I2(n13_adj_4575), 
            .I3(n11_adj_4573), .O(n33239));
    defparam i27565_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_23__I_0_add_1043_10_lut (.I0(GND_net), .I1(n1541), 
            .I2(VCC_net), .I3(n25267), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27864_4_lut (.I0(n9_adj_4571), .I1(n7_adj_4569), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n33540));
    defparam i27864_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i28049_4_lut (.I0(n15_adj_4576), .I1(n13_adj_4575), .I2(n11_adj_4573), 
            .I3(n33540), .O(n33725));
    defparam i28049_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY encoder0_position_23__I_0_add_1043_10 (.CI(n25267), .I0(n1541), 
            .I1(VCC_net), .CO(n25268));
    SB_LUT4 i12766_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n4216), .I3(GND_net), .O(n16875));   // verilog/coms.v(127[12] 300[6])
    defparam i12766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_9_lut (.I0(GND_net), .I1(n1542), 
            .I2(VCC_net), .I3(n25266), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_9 (.CI(n25266), .I0(n1542), 
            .I1(VCC_net), .CO(n25267));
    SB_LUT4 encoder0_position_23__I_0_add_1043_8_lut (.I0(GND_net), .I1(n1543), 
            .I2(VCC_net), .I3(n25265), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_8 (.CI(n25265), .I0(n1543), 
            .I1(VCC_net), .CO(n25266));
    SB_LUT4 encoder0_position_23__I_0_add_1043_7_lut (.I0(GND_net), .I1(n1544), 
            .I2(GND_net), .I3(n25264), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28047_4_lut (.I0(n21_adj_4579), .I1(n19_adj_4578), .I2(n17_adj_4577), 
            .I3(n33725), .O(n33723));
    defparam i28047_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY encoder0_position_23__I_0_add_1043_7 (.CI(n25264), .I0(n1544), 
            .I1(GND_net), .CO(n25265));
    SB_LUT4 i27567_4_lut (.I0(n27), .I1(n25_adj_4581), .I2(n23_adj_4580), 
            .I3(n33723), .O(n33241));
    defparam i27567_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_558_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4567));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 encoder0_position_23__I_0_add_1043_6_lut (.I0(GND_net), .I1(n1545), 
            .I2(GND_net), .I3(n25263), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28197_3_lut (.I0(n4_adj_4567), .I1(pwm_setpoint[13]), .I2(n27), 
            .I3(GND_net), .O(n33873));   // verilog/pwm.v(21[8:24])
    defparam i28197_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1043_6 (.CI(n25263), .I0(n1545), 
            .I1(GND_net), .CO(n25264));
    SB_LUT4 encoder0_position_23__I_0_add_1043_5_lut (.I0(GND_net), .I1(n1546), 
            .I2(VCC_net), .I3(n25262), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_5 (.CI(n25262), .I0(n1546), 
            .I1(VCC_net), .CO(n25263));
    SB_LUT4 encoder0_position_23__I_0_add_1043_4_lut (.I0(GND_net), .I1(n1547), 
            .I2(GND_net), .I3(n25261), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_4 (.CI(n25261), .I0(n1547), 
            .I1(GND_net), .CO(n25262));
    SB_LUT4 encoder0_position_23__I_0_add_1043_3_lut (.I0(GND_net), .I1(n1548), 
            .I2(VCC_net), .I3(n25260), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_558_i30_3_lut (.I0(n12_adj_4574), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30_adj_4583));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28198_3_lut (.I0(n33873), .I1(pwm_setpoint[14]), .I2(n29_adj_4582), 
            .I3(GND_net), .O(n33874));   // verilog/pwm.v(21[8:24])
    defparam i28198_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1043_3 (.CI(n25260), .I0(n1548), 
            .I1(VCC_net), .CO(n25261));
    SB_LUT4 i27561_4_lut (.I0(n33_adj_4585), .I1(n31_adj_4584), .I2(n29_adj_4582), 
            .I3(n33239), .O(n33235));
    defparam i27561_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_23__I_0_add_1043_2_lut (.I0(GND_net), .I1(n439), 
            .I2(GND_net), .I3(VCC_net), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_2 (.CI(VCC_net), .I0(n439), 
            .I1(GND_net), .CO(n25260));
    SB_LUT4 encoder0_position_23__I_0_add_990_18_lut (.I0(GND_net), .I1(n1454), 
            .I2(VCC_net), .I3(n25259), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_990_17_lut (.I0(GND_net), .I1(n1455), 
            .I2(VCC_net), .I3(n25258), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28300_4_lut (.I0(n30_adj_4583), .I1(n10_adj_4572), .I2(n35), 
            .I3(n33233), .O(n33976));   // verilog/pwm.v(21[8:24])
    defparam i28300_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28174_3_lut (.I0(n33874), .I1(pwm_setpoint[15]), .I2(n31_adj_4584), 
            .I3(GND_net), .O(n33850));   // verilog/pwm.v(21[8:24])
    defparam i28174_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_17 (.CI(n25258), .I0(n1455), 
            .I1(VCC_net), .CO(n25259));
    SB_LUT4 encoder0_position_23__I_0_add_990_16_lut (.I0(GND_net), .I1(n1456), 
            .I2(VCC_net), .I3(n25257), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28199_3_lut (.I0(n6_adj_4568), .I1(pwm_setpoint[10]), .I2(n21_adj_4579), 
            .I3(GND_net), .O(n33875));   // verilog/pwm.v(21[8:24])
    defparam i28199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28200_3_lut (.I0(n33875), .I1(pwm_setpoint[11]), .I2(n23_adj_4580), 
            .I3(GND_net), .O(n33876));   // verilog/pwm.v(21[8:24])
    defparam i28200_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_16 (.CI(n25257), .I0(n1456), 
            .I1(VCC_net), .CO(n25258));
    SB_LUT4 i27854_4_lut (.I0(n23_adj_4580), .I1(n21_adj_4579), .I2(n19_adj_4578), 
            .I3(n33247), .O(n33530));
    defparam i27854_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 encoder0_position_23__I_0_add_990_15_lut (.I0(GND_net), .I1(n1457), 
            .I2(VCC_net), .I3(n25256), .O(n1510)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28097_3_lut (.I0(n8_adj_4570), .I1(pwm_setpoint[9]), .I2(n19_adj_4578), 
            .I3(GND_net), .O(n33773));   // verilog/pwm.v(21[8:24])
    defparam i28097_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_15 (.CI(n25256), .I0(n1457), 
            .I1(VCC_net), .CO(n25257));
    SB_LUT4 encoder0_position_23__I_0_add_990_14_lut (.I0(GND_net), .I1(n1458), 
            .I2(VCC_net), .I3(n25255), .O(n1511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_14 (.CI(n25255), .I0(n1458), 
            .I1(VCC_net), .CO(n25256));
    SB_LUT4 i28172_3_lut (.I0(n33876), .I1(pwm_setpoint[12]), .I2(n25_adj_4581), 
            .I3(GND_net), .O(n33848));   // verilog/pwm.v(21[8:24])
    defparam i28172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_990_13_lut (.I0(GND_net), .I1(n1459), 
            .I2(VCC_net), .I3(n25254), .O(n1512)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_13 (.CI(n25254), .I0(n1459), 
            .I1(VCC_net), .CO(n25255));
    SB_LUT4 i28131_4_lut (.I0(n33_adj_4585), .I1(n31_adj_4584), .I2(n29_adj_4582), 
            .I3(n33241), .O(n33807));
    defparam i28131_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_990_12_lut (.I0(GND_net), .I1(n1460), 
            .I2(VCC_net), .I3(n25253), .O(n1513)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28349_4_lut (.I0(n33850), .I1(n33976), .I2(n35), .I3(n33235), 
            .O(n34025));   // verilog/pwm.v(21[8:24])
    defparam i28349_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28193_4_lut (.I0(n33848), .I1(n33773), .I2(n25_adj_4581), 
            .I3(n33530), .O(n33869));   // verilog/pwm.v(21[8:24])
    defparam i28193_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28353_4_lut (.I0(n33869), .I1(n34025), .I2(n35), .I3(n33807), 
            .O(n34029));   // verilog/pwm.v(21[8:24])
    defparam i28353_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_23__I_0_add_990_12 (.CI(n25253), .I0(n1460), 
            .I1(VCC_net), .CO(n25254));
    SB_LUT4 i28354_3_lut (.I0(n34029), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n34030));   // verilog/pwm.v(21[8:24])
    defparam i28354_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_add_990_11_lut (.I0(GND_net), .I1(n1461), 
            .I2(VCC_net), .I3(n25252), .O(n1514)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_11 (.CI(n25252), .I0(n1461), 
            .I1(VCC_net), .CO(n25253));
    SB_LUT4 encoder0_position_23__I_0_add_990_10_lut (.I0(GND_net), .I1(n1462), 
            .I2(VCC_net), .I3(n25251), .O(n1515)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28352_3_lut (.I0(n34030), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n34028));   // verilog/pwm.v(21[8:24])
    defparam i28352_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_990_10 (.CI(n25251), .I0(n1462), 
            .I1(VCC_net), .CO(n25252));
    SB_LUT4 encoder0_position_23__I_0_add_990_9_lut (.I0(GND_net), .I1(n1463), 
            .I2(VCC_net), .I3(n25250), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_9 (.CI(n25250), .I0(n1463), 
            .I1(VCC_net), .CO(n25251));
    SB_LUT4 encoder0_position_23__I_0_add_990_8_lut (.I0(GND_net), .I1(n1464), 
            .I2(VCC_net), .I3(n25249), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_8 (.CI(n25249), .I0(n1464), 
            .I1(VCC_net), .CO(n25250));
    SB_LUT4 encoder0_position_23__I_0_add_990_7_lut (.I0(GND_net), .I1(n1465), 
            .I2(GND_net), .I3(n25248), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_7 (.CI(n25248), .I0(n1465), 
            .I1(GND_net), .CO(n25249));
    SB_LUT4 encoder0_position_23__I_0_add_990_6_lut (.I0(GND_net), .I1(n1466), 
            .I2(GND_net), .I3(n25247), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28280_3_lut (.I0(n34028), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n33956));   // verilog/pwm.v(21[8:24])
    defparam i28280_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_990_6 (.CI(n25247), .I0(n1466), 
            .I1(GND_net), .CO(n25248));
    SB_LUT4 encoder0_position_23__I_0_add_990_5_lut (.I0(GND_net), .I1(n1467), 
            .I2(VCC_net), .I3(n25246), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_5 (.CI(n25246), .I0(n1467), 
            .I1(VCC_net), .CO(n25247));
    SB_LUT4 encoder0_position_23__I_0_add_990_4_lut (.I0(GND_net), .I1(n1468), 
            .I2(GND_net), .I3(n25245), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12767_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n4216), .I3(GND_net), .O(n16876));   // verilog/coms.v(127[12] 300[6])
    defparam i12767_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_4 (.CI(n25245), .I0(n1468), 
            .I1(GND_net), .CO(n25246));
    SB_LUT4 encoder0_position_23__I_0_add_990_3_lut (.I0(GND_net), .I1(n1469), 
            .I2(VCC_net), .I3(n25244), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_3 (.CI(n25244), .I0(n1469), 
            .I1(VCC_net), .CO(n25245));
    SB_LUT4 encoder0_position_23__I_0_add_990_2_lut (.I0(GND_net), .I1(n438), 
            .I2(GND_net), .I3(VCC_net), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_2 (.CI(VCC_net), .I0(n438), 
            .I1(GND_net), .CO(n25244));
    SB_LUT4 encoder0_position_23__I_0_add_937_17_lut (.I0(GND_net), .I1(n1376), 
            .I2(VCC_net), .I3(n25243), .O(n1429)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_937_16_lut (.I0(GND_net), .I1(n1377), 
            .I2(VCC_net), .I3(n25242), .O(n1430)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_16 (.CI(n25242), .I0(n1377), 
            .I1(VCC_net), .CO(n25243));
    SB_LUT4 encoder0_position_23__I_0_add_937_15_lut (.I0(GND_net), .I1(n1378), 
            .I2(VCC_net), .I3(n25241), .O(n1431)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_15 (.CI(n25241), .I0(n1378), 
            .I1(VCC_net), .CO(n25242));
    SB_LUT4 encoder0_position_23__I_0_add_937_14_lut (.I0(GND_net), .I1(n1379), 
            .I2(VCC_net), .I3(n25240), .O(n1432)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_14 (.CI(n25240), .I0(n1379), 
            .I1(VCC_net), .CO(n25241));
    SB_LUT4 encoder0_position_23__I_0_add_937_13_lut (.I0(GND_net), .I1(n1380), 
            .I2(VCC_net), .I3(n25239), .O(n1433)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_13 (.CI(n25239), .I0(n1380), 
            .I1(VCC_net), .CO(n25240));
    SB_LUT4 encoder0_position_23__I_0_add_937_12_lut (.I0(GND_net), .I1(n1381), 
            .I2(VCC_net), .I3(n25238), .O(n1434)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_12 (.CI(n25238), .I0(n1381), 
            .I1(VCC_net), .CO(n25239));
    SB_LUT4 encoder0_position_23__I_0_add_937_11_lut (.I0(GND_net), .I1(n1382), 
            .I2(VCC_net), .I3(n25237), .O(n1435)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_11 (.CI(n25237), .I0(n1382), 
            .I1(VCC_net), .CO(n25238));
    SB_LUT4 i12768_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n4216), .I3(GND_net), .O(n16877));   // verilog/coms.v(127[12] 300[6])
    defparam i12768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_937_10_lut (.I0(GND_net), .I1(n1383), 
            .I2(VCC_net), .I3(n25236), .O(n1436)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_4611), .I3(n25709), .O(n22_adj_4508)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_6 (.CI(n25709), 
            .I0(GND_net), .I1(n22_adj_4611), .CO(n25710));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_4612), .I3(n25708), .O(n23_adj_4507)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_10 (.CI(n25236), .I0(n1383), 
            .I1(VCC_net), .CO(n25237));
    SB_LUT4 encoder0_position_23__I_0_add_937_9_lut (.I0(GND_net), .I1(n1384), 
            .I2(VCC_net), .I3(n25235), .O(n1437)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12769_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n4216), .I3(GND_net), .O(n16878));   // verilog/coms.v(127[12] 300[6])
    defparam i12769_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_937_9 (.CI(n25235), .I0(n1384), 
            .I1(VCC_net), .CO(n25236));
    SB_LUT4 encoder0_position_23__I_0_add_937_8_lut (.I0(GND_net), .I1(n1385), 
            .I2(VCC_net), .I3(n25234), .O(n1438)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_8 (.CI(n25234), .I0(n1385), 
            .I1(VCC_net), .CO(n25235));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_5 (.CI(n25708), 
            .I0(GND_net), .I1(n23_adj_4612), .CO(n25709));
    SB_LUT4 encoder0_position_23__I_0_add_937_7_lut (.I0(GND_net), .I1(n1386), 
            .I2(GND_net), .I3(n25233), .O(n1439)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_7 (.CI(n25233), .I0(n1386), 
            .I1(GND_net), .CO(n25234));
    SB_LUT4 encoder0_position_23__I_0_add_937_6_lut (.I0(GND_net), .I1(n1387), 
            .I2(GND_net), .I3(n25232), .O(n1440)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_6 (.CI(n25232), .I0(n1387), 
            .I1(GND_net), .CO(n25233));
    SB_LUT4 encoder0_position_23__I_0_add_937_5_lut (.I0(GND_net), .I1(n1388), 
            .I2(VCC_net), .I3(n25231), .O(n1441)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_5 (.CI(n25231), .I0(n1388), 
            .I1(VCC_net), .CO(n25232));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_4613), .I3(n25707), .O(n24_adj_4506)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_937_4_lut (.I0(GND_net), .I1(n1389), 
            .I2(GND_net), .I3(n25230), .O(n1442)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12770_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n4216), .I3(GND_net), .O(n16879));   // verilog/coms.v(127[12] 300[6])
    defparam i12770_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_937_4 (.CI(n25230), .I0(n1389), 
            .I1(GND_net), .CO(n25231));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_4 (.CI(n25707), 
            .I0(GND_net), .I1(n24_adj_4613), .CO(n25708));
    SB_LUT4 encoder0_position_23__I_0_add_937_3_lut (.I0(GND_net), .I1(n1390), 
            .I2(VCC_net), .I3(n25229), .O(n1443)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12771_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n4216), .I3(GND_net), .O(n16880));   // verilog/coms.v(127[12] 300[6])
    defparam i12771_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_937_3 (.CI(n25229), .I0(n1390), 
            .I1(VCC_net), .CO(n25230));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_4614), .I3(n25706), .O(n25_adj_4503)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_937_2_lut (.I0(GND_net), .I1(n437), 
            .I2(GND_net), .I3(VCC_net), .O(n1444)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12772_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n4216), .I3(GND_net), .O(n16881));   // verilog/coms.v(127[12] 300[6])
    defparam i12772_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_937_2 (.CI(VCC_net), .I0(n437), 
            .I1(GND_net), .CO(n25229));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_3 (.CI(n25706), 
            .I0(GND_net), .I1(n25_adj_4614), .CO(n25707));
    SB_LUT4 i12773_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n4216), .I3(GND_net), .O(n16882));   // verilog/coms.v(127[12] 300[6])
    defparam i12773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_884_16_lut (.I0(GND_net), .I1(n1298), 
            .I2(VCC_net), .I3(n25228), .O(n1351)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_884_15_lut (.I0(GND_net), .I1(n1299), 
            .I2(VCC_net), .I3(n25227), .O(n1352)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_15 (.CI(n25227), .I0(n1299), 
            .I1(VCC_net), .CO(n25228));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n25706));
    SB_CARRY add_486_4 (.CI(n24926), .I0(n34501), .I1(n23), .CO(n24927));
    SB_LUT4 i12775_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n4216), .I3(GND_net), .O(n16884));   // verilog/coms.v(127[12] 300[6])
    defparam i12775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_486_3_lut (.I0(duty[1]), .I1(n34501), .I2(n24), .I3(n24925), 
            .O(pwm_setpoint_22__N_3[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12776_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n4216), .I3(GND_net), .O(n16885));   // verilog/coms.v(127[12] 300[6])
    defparam i12776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12777_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n4216), .I3(GND_net), .O(n16886));   // verilog/coms.v(127[12] 300[6])
    defparam i12777_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[0]));   // verilog/TinyFPGA_B.v(201[10] 204[6])
    SB_LUT4 encoder0_position_23__I_0_add_884_14_lut (.I0(GND_net), .I1(n1300), 
            .I2(VCC_net), .I3(n25226), .O(n1353)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12778_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n4216), .I3(GND_net), .O(n16887));   // verilog/coms.v(127[12] 300[6])
    defparam i12778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12779_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n4216), .I3(GND_net), .O(n16888));   // verilog/coms.v(127[12] 300[6])
    defparam i12779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12780_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n4216), .I3(GND_net), .O(n16889));   // verilog/coms.v(127[12] 300[6])
    defparam i12780_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_14 (.CI(n25226), .I0(n1300), 
            .I1(VCC_net), .CO(n25227));
    SB_LUT4 encoder0_position_23__I_0_add_884_13_lut (.I0(GND_net), .I1(n1301), 
            .I2(VCC_net), .I3(n25225), .O(n1354)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12781_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n4216), .I3(GND_net), .O(n16890));   // verilog/coms.v(127[12] 300[6])
    defparam i12781_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_13 (.CI(n25225), .I0(n1301), 
            .I1(VCC_net), .CO(n25226));
    SB_CARRY add_486_3 (.CI(n24925), .I0(n34501), .I1(n24), .CO(n24926));
    SB_LUT4 encoder0_position_23__I_0_add_884_12_lut (.I0(GND_net), .I1(n1302), 
            .I2(VCC_net), .I3(n25224), .O(n1355)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12782_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n4216), .I3(GND_net), .O(n16891));   // verilog/coms.v(127[12] 300[6])
    defparam i12782_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_12 (.CI(n25224), .I0(n1302), 
            .I1(VCC_net), .CO(n25225));
    SB_LUT4 add_486_2_lut (.I0(duty[0]), .I1(n34501), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_3[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_486_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_884_11_lut (.I0(GND_net), .I1(n1303), 
            .I2(VCC_net), .I3(n25223), .O(n1356)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_11 (.CI(n25223), .I0(n1303), 
            .I1(VCC_net), .CO(n25224));
    SB_LUT4 encoder0_position_23__I_0_add_884_10_lut (.I0(GND_net), .I1(n1304), 
            .I2(VCC_net), .I3(n25222), .O(n1357)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_10 (.CI(n25222), .I0(n1304), 
            .I1(VCC_net), .CO(n25223));
    SB_LUT4 i12783_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n4216), .I3(GND_net), .O(n16892));   // verilog/coms.v(127[12] 300[6])
    defparam i12783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_884_9_lut (.I0(GND_net), .I1(n1305), 
            .I2(VCC_net), .I3(n25221), .O(n1358)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_9 (.CI(n25221), .I0(n1305), 
            .I1(VCC_net), .CO(n25222));
    SB_LUT4 encoder0_position_23__I_0_add_884_8_lut (.I0(GND_net), .I1(n1306), 
            .I2(VCC_net), .I3(n25220), .O(n1359)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_8 (.CI(n25220), .I0(n1306), 
            .I1(VCC_net), .CO(n25221));
    SB_LUT4 encoder0_position_23__I_0_add_884_7_lut (.I0(GND_net), .I1(n1307), 
            .I2(GND_net), .I3(n25219), .O(n1360)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_7 (.CI(n25219), .I0(n1307), 
            .I1(GND_net), .CO(n25220));
    SB_CARRY add_486_2 (.CI(VCC_net), .I0(n34501), .I1(n25), .CO(n24925));
    SB_LUT4 encoder0_position_23__I_0_add_884_6_lut (.I0(GND_net), .I1(n1308), 
            .I2(GND_net), .I3(n25218), .O(n1361)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_6 (.CI(n25218), .I0(n1308), 
            .I1(GND_net), .CO(n25219));
    SB_LUT4 encoder0_position_23__I_0_add_884_5_lut (.I0(GND_net), .I1(n1309), 
            .I2(VCC_net), .I3(n25217), .O(n1362)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_5 (.CI(n25217), .I0(n1309), 
            .I1(VCC_net), .CO(n25218));
    SB_LUT4 encoder0_position_23__I_0_add_884_4_lut (.I0(GND_net), .I1(n1310), 
            .I2(GND_net), .I3(n25216), .O(n1363)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_4 (.CI(n25216), .I0(n1310), 
            .I1(GND_net), .CO(n25217));
    SB_LUT4 encoder0_position_23__I_0_add_884_3_lut (.I0(GND_net), .I1(n1311), 
            .I2(VCC_net), .I3(n25215), .O(n1364)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12784_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n4216), .I3(GND_net), .O(n16893));   // verilog/coms.v(127[12] 300[6])
    defparam i12784_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_3 (.CI(n25215), .I0(n1311), 
            .I1(VCC_net), .CO(n25216));
    SB_LUT4 encoder0_position_23__I_0_add_884_2_lut (.I0(GND_net), .I1(n436), 
            .I2(GND_net), .I3(VCC_net), .O(n1365)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_2 (.CI(VCC_net), .I0(n436), 
            .I1(GND_net), .CO(n25215));
    SB_LUT4 encoder0_position_23__I_0_add_831_15_lut (.I0(GND_net), .I1(n1220), 
            .I2(VCC_net), .I3(n25214), .O(n1273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12785_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n4216), .I3(GND_net), .O(n16894));   // verilog/coms.v(127[12] 300[6])
    defparam i12785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_14_lut (.I0(GND_net), .I1(n1221), 
            .I2(VCC_net), .I3(n25213), .O(n1274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_14 (.CI(n25213), .I0(n1221), 
            .I1(VCC_net), .CO(n25214));
    SB_LUT4 encoder0_position_23__I_0_add_831_13_lut (.I0(GND_net), .I1(n1222), 
            .I2(VCC_net), .I3(n25212), .O(n1275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_13 (.CI(n25212), .I0(n1222), 
            .I1(VCC_net), .CO(n25213));
    SB_LUT4 encoder0_position_23__I_0_add_831_12_lut (.I0(GND_net), .I1(n1223), 
            .I2(VCC_net), .I3(n25211), .O(n1276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12787_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n4216), .I3(GND_net), .O(n16896));   // verilog/coms.v(127[12] 300[6])
    defparam i12787_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_831_12 (.CI(n25211), .I0(n1223), 
            .I1(VCC_net), .CO(n25212));
    SB_LUT4 encoder0_position_23__I_0_add_831_11_lut (.I0(GND_net), .I1(n1224), 
            .I2(VCC_net), .I3(n25210), .O(n1277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_11 (.CI(n25210), .I0(n1224), 
            .I1(VCC_net), .CO(n25211));
    SB_LUT4 encoder0_position_23__I_0_add_831_10_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n25209), .O(n1278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_10 (.CI(n25209), .I0(n1225), 
            .I1(VCC_net), .CO(n25210));
    SB_LUT4 encoder0_position_23__I_0_add_831_9_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n25208), .O(n1279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_9 (.CI(n25208), .I0(n1226), 
            .I1(VCC_net), .CO(n25209));
    SB_LUT4 i12788_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4216), .I3(GND_net), .O(n16897));   // verilog/coms.v(127[12] 300[6])
    defparam i12788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_8_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n25207), .O(n1280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_8 (.CI(n25207), .I0(n1227), 
            .I1(VCC_net), .CO(n25208));
    SB_LUT4 encoder0_position_23__I_0_add_831_7_lut (.I0(GND_net), .I1(n1228), 
            .I2(GND_net), .I3(n25206), .O(n1281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_7 (.CI(n25206), .I0(n1228), 
            .I1(GND_net), .CO(n25207));
    SB_LUT4 encoder0_position_23__I_0_add_831_6_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n25205), .O(n1282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_6 (.CI(n25205), .I0(n1229), 
            .I1(GND_net), .CO(n25206));
    SB_LUT4 encoder0_position_23__I_0_add_831_5_lut (.I0(GND_net), .I1(n1230), 
            .I2(VCC_net), .I3(n25204), .O(n1283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_5 (.CI(n25204), .I0(n1230), 
            .I1(VCC_net), .CO(n25205));
    SB_LUT4 encoder0_position_23__I_0_add_831_4_lut (.I0(GND_net), .I1(n1231), 
            .I2(GND_net), .I3(n25203), .O(n1284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_4 (.CI(n25203), .I0(n1231), 
            .I1(GND_net), .CO(n25204));
    SB_LUT4 encoder0_position_23__I_0_add_831_3_lut (.I0(GND_net), .I1(n1232), 
            .I2(VCC_net), .I3(n25202), .O(n1285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_3 (.CI(n25202), .I0(n1232), 
            .I1(VCC_net), .CO(n25203));
    SB_LUT4 encoder0_position_23__I_0_add_831_2_lut (.I0(GND_net), .I1(n435), 
            .I2(GND_net), .I3(VCC_net), .O(n1286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_2 (.CI(VCC_net), .I0(n435), 
            .I1(GND_net), .CO(n25202));
    SB_LUT4 encoder0_position_23__I_0_add_778_14_lut (.I0(GND_net), .I1(n1142), 
            .I2(VCC_net), .I3(n25201), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_778_13_lut (.I0(GND_net), .I1(n1143), 
            .I2(VCC_net), .I3(n25200), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_13 (.CI(n25200), .I0(n1143), 
            .I1(VCC_net), .CO(n25201));
    SB_LUT4 encoder0_position_23__I_0_add_778_12_lut (.I0(GND_net), .I1(n1144), 
            .I2(VCC_net), .I3(n25199), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4607));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 encoder0_position_23__I_0_add_460_8_lut (.I0(n34057), .I1(n674), 
            .I2(VCC_net), .I3(n25907), .O(n752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_add_460_7_lut (.I0(GND_net), .I1(n675), 
            .I2(GND_net), .I3(n25906), .O(n728)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_12 (.CI(n25199), .I0(n1144), 
            .I1(VCC_net), .CO(n25200));
    SB_LUT4 encoder0_position_23__I_0_add_778_11_lut (.I0(GND_net), .I1(n1145), 
            .I2(VCC_net), .I3(n25198), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_11 (.CI(n25198), .I0(n1145), 
            .I1(VCC_net), .CO(n25199));
    SB_LUT4 encoder0_position_23__I_0_add_778_10_lut (.I0(GND_net), .I1(n1146), 
            .I2(VCC_net), .I3(n25197), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_7 (.CI(n25906), .I0(n675), 
            .I1(GND_net), .CO(n25907));
    SB_LUT4 encoder0_position_23__I_0_add_460_6_lut (.I0(GND_net), .I1(n676), 
            .I2(GND_net), .I3(n25905), .O(n729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_10 (.CI(n25197), .I0(n1146), 
            .I1(VCC_net), .CO(n25198));
    SB_CARRY encoder0_position_23__I_0_add_460_6 (.CI(n25905), .I0(n676), 
            .I1(GND_net), .CO(n25906));
    SB_LUT4 encoder0_position_23__I_0_add_460_5_lut (.I0(GND_net), .I1(n677), 
            .I2(VCC_net), .I3(n25904), .O(n730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_5 (.CI(n25904), .I0(n677), 
            .I1(VCC_net), .CO(n25905));
    SB_LUT4 encoder0_position_23__I_0_add_460_4_lut (.I0(GND_net), .I1(n678), 
            .I2(GND_net), .I3(n25903), .O(n731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_4 (.CI(n25903), .I0(n678), 
            .I1(GND_net), .CO(n25904));
    SB_LUT4 encoder0_position_23__I_0_add_460_3_lut (.I0(GND_net), .I1(n679), 
            .I2(VCC_net), .I3(n25902), .O(n732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_3 (.CI(n25902), .I0(n679), 
            .I1(VCC_net), .CO(n25903));
    SB_LUT4 encoder0_position_23__I_0_add_460_2_lut (.I0(GND_net), .I1(n428), 
            .I2(GND_net), .I3(VCC_net), .O(n733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_2 (.CI(VCC_net), .I0(n428), 
            .I1(GND_net), .CO(n25902));
    SB_LUT4 encoder0_position_23__I_0_add_778_9_lut (.I0(GND_net), .I1(n1147), 
            .I2(VCC_net), .I3(n25196), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n3_adj_4532), .I3(n25076), .O(displacement_23__N_50[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_9 (.CI(n25196), .I0(n1147), 
            .I1(VCC_net), .CO(n25197));
    SB_LUT4 encoder0_position_23__I_0_add_778_8_lut (.I0(GND_net), .I1(n1148), 
            .I2(VCC_net), .I3(n25195), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_8 (.CI(n25195), .I0(n1148), 
            .I1(VCC_net), .CO(n25196));
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_778_7_lut (.I0(GND_net), .I1(n1149), 
            .I2(GND_net), .I3(n25194), .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_7 (.CI(n25194), .I0(n1149), 
            .I1(GND_net), .CO(n25195));
    SB_LUT4 encoder0_position_23__I_0_add_778_6_lut (.I0(GND_net), .I1(n1150), 
            .I2(GND_net), .I3(n25193), .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_6 (.CI(n25193), .I0(n1150), 
            .I1(GND_net), .CO(n25194));
    SB_LUT4 encoder0_position_23__I_0_add_778_5_lut (.I0(GND_net), .I1(n1151), 
            .I2(VCC_net), .I3(n25192), .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_5 (.CI(n25192), .I0(n1151), 
            .I1(VCC_net), .CO(n25193));
    SB_LUT4 encoder0_position_23__I_0_add_778_4_lut (.I0(GND_net), .I1(n1152), 
            .I2(GND_net), .I3(n25191), .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_4 (.CI(n25191), .I0(n1152), 
            .I1(GND_net), .CO(n25192));
    SB_LUT4 encoder0_position_23__I_0_add_778_3_lut (.I0(GND_net), .I1(n1153), 
            .I2(VCC_net), .I3(n25190), .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4532), .I3(n25075), .O(displacement_23__N_50[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n25075), .I0(encoder1_position[22]), 
            .I1(n3_adj_4532), .CO(n25076));
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n3_adj_4532), .I3(n25074), .O(displacement_23__N_50[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_3 (.CI(n25190), .I0(n1153), 
            .I1(VCC_net), .CO(n25191));
    SB_LUT4 encoder0_position_23__I_0_add_778_2_lut (.I0(GND_net), .I1(n434), 
            .I2(GND_net), .I3(VCC_net), .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_2 (.CI(VCC_net), .I0(n434), 
            .I1(GND_net), .CO(n25190));
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n25074), .I0(encoder1_position[21]), 
            .I1(n3_adj_4532), .CO(n25075));
    SB_LUT4 encoder0_position_23__I_0_add_725_13_lut (.I0(GND_net), .I1(n1064), 
            .I2(VCC_net), .I3(n25189), .O(n1117)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_12_lut (.I0(GND_net), .I1(n1065), 
            .I2(VCC_net), .I3(n25188), .O(n1118)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_12 (.CI(n25188), .I0(n1065), 
            .I1(VCC_net), .CO(n25189));
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4528), .I3(n25073), .O(displacement_23__N_50[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_11_lut (.I0(GND_net), .I1(n1066), 
            .I2(VCC_net), .I3(n25187), .O(n1119)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n25073), .I0(encoder1_position[20]), 
            .I1(n5_adj_4528), .CO(n25074));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4536), .I3(n25072), .O(displacement_23__N_50[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_11 (.CI(n25187), .I0(n1066), 
            .I1(VCC_net), .CO(n25188));
    SB_LUT4 encoder0_position_23__I_0_add_725_10_lut (.I0(GND_net), .I1(n1067), 
            .I2(VCC_net), .I3(n25186), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_10 (.CI(n25186), .I0(n1067), 
            .I1(VCC_net), .CO(n25187));
    SB_LUT4 encoder0_position_23__I_0_add_725_9_lut (.I0(GND_net), .I1(n1068), 
            .I2(VCC_net), .I3(n25185), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_9 (.CI(n25185), .I0(n1068), 
            .I1(VCC_net), .CO(n25186));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4606));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n25072), .I0(encoder1_position[19]), 
            .I1(n6_adj_4536), .CO(n25073));
    SB_LUT4 encoder0_position_23__I_0_add_725_8_lut (.I0(GND_net), .I1(n1069), 
            .I2(VCC_net), .I3(n25184), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_8 (.CI(n25184), .I0(n1069), 
            .I1(VCC_net), .CO(n25185));
    SB_LUT4 encoder0_position_23__I_0_add_725_7_lut (.I0(GND_net), .I1(n1070), 
            .I2(GND_net), .I3(n25183), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_7 (.CI(n25183), .I0(n1070), 
            .I1(GND_net), .CO(n25184));
    SB_LUT4 encoder0_position_23__I_0_add_725_6_lut (.I0(GND_net), .I1(n1071), 
            .I2(GND_net), .I3(n25182), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_6 (.CI(n25182), .I0(n1071), 
            .I1(GND_net), .CO(n25183));
    SB_LUT4 encoder0_position_23__I_0_add_725_5_lut (.I0(GND_net), .I1(n1072), 
            .I2(VCC_net), .I3(n25181), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_5 (.CI(n25181), .I0(n1072), 
            .I1(VCC_net), .CO(n25182));
    SB_LUT4 encoder0_position_23__I_0_add_725_4_lut (.I0(GND_net), .I1(n1073), 
            .I2(GND_net), .I3(n25180), .O(n1126)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_4 (.CI(n25180), .I0(n1073), 
            .I1(GND_net), .CO(n25181));
    SB_LUT4 encoder0_position_23__I_0_add_725_3_lut (.I0(GND_net), .I1(n1074), 
            .I2(VCC_net), .I3(n25179), .O(n1127)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_3 (.CI(n25179), .I0(n1074), 
            .I1(VCC_net), .CO(n25180));
    SB_LUT4 encoder0_position_23__I_0_add_725_2_lut (.I0(GND_net), .I1(n433), 
            .I2(GND_net), .I3(VCC_net), .O(n1128)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4537), .I3(n25071), .O(displacement_23__N_50[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n25071), .I0(encoder1_position[18]), 
            .I1(n7_adj_4537), .CO(n25072));
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4538), .I3(n25070), .O(displacement_23__N_50[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_2 (.CI(VCC_net), .I0(n433), 
            .I1(GND_net), .CO(n25179));
    SB_LUT4 encoder0_position_23__I_0_add_672_12_lut (.I0(GND_net), .I1(n986), 
            .I2(VCC_net), .I3(n25178), .O(n1039)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_672_11_lut (.I0(GND_net), .I1(n987), 
            .I2(VCC_net), .I3(n25177), .O(n1040)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_11 (.CI(n25177), .I0(n987), 
            .I1(VCC_net), .CO(n25178));
    SB_LUT4 encoder0_position_23__I_0_add_672_10_lut (.I0(GND_net), .I1(n988), 
            .I2(VCC_net), .I3(n25176), .O(n1041)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_10 (.CI(n25176), .I0(n988), 
            .I1(VCC_net), .CO(n25177));
    SB_LUT4 encoder0_position_23__I_0_add_672_9_lut (.I0(GND_net), .I1(n989), 
            .I2(VCC_net), .I3(n25175), .O(n1042)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_9 (.CI(n25175), .I0(n989), 
            .I1(VCC_net), .CO(n25176));
    SB_LUT4 encoder0_position_23__I_0_add_672_8_lut (.I0(GND_net), .I1(n990), 
            .I2(VCC_net), .I3(n25174), .O(n1043)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n25070), .I0(encoder1_position[17]), 
            .I1(n8_adj_4538), .CO(n25071));
    SB_CARRY encoder0_position_23__I_0_add_672_8 (.CI(n25174), .I0(n990), 
            .I1(VCC_net), .CO(n25175));
    SB_LUT4 encoder0_position_23__I_0_add_672_7_lut (.I0(GND_net), .I1(n991), 
            .I2(GND_net), .I3(n25173), .O(n1044)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_7 (.CI(n25173), .I0(n991), 
            .I1(GND_net), .CO(n25174));
    SB_LUT4 encoder0_position_23__I_0_add_672_6_lut (.I0(GND_net), .I1(n992), 
            .I2(GND_net), .I3(n25172), .O(n1045)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_6 (.CI(n25172), .I0(n992), 
            .I1(GND_net), .CO(n25173));
    SB_LUT4 encoder0_position_23__I_0_add_672_5_lut (.I0(GND_net), .I1(n993), 
            .I2(VCC_net), .I3(n25171), .O(n1046)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_5 (.CI(n25171), .I0(n993), 
            .I1(VCC_net), .CO(n25172));
    SB_LUT4 encoder0_position_23__I_0_add_672_4_lut (.I0(GND_net), .I1(n994), 
            .I2(GND_net), .I3(n25170), .O(n1047)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_4 (.CI(n25170), .I0(n994), 
            .I1(GND_net), .CO(n25171));
    SB_LUT4 encoder0_position_23__I_0_add_672_3_lut (.I0(GND_net), .I1(n995), 
            .I2(VCC_net), .I3(n25169), .O(n1048)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_3 (.CI(n25169), .I0(n995), 
            .I1(VCC_net), .CO(n25170));
    SB_LUT4 encoder0_position_23__I_0_add_672_2_lut (.I0(GND_net), .I1(n432), 
            .I2(GND_net), .I3(VCC_net), .O(n1049)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_2 (.CI(VCC_net), .I0(n432), 
            .I1(GND_net), .CO(n25169));
    SB_LUT4 encoder0_position_23__I_0_add_619_11_lut (.I0(GND_net), .I1(n908), 
            .I2(VCC_net), .I3(n25168), .O(n961)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_619_10_lut (.I0(GND_net), .I1(n909), 
            .I2(VCC_net), .I3(n25167), .O(n962)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_10 (.CI(n25167), .I0(n909), 
            .I1(VCC_net), .CO(n25168));
    SB_LUT4 encoder0_position_23__I_0_add_619_9_lut (.I0(GND_net), .I1(n910), 
            .I2(VCC_net), .I3(n25166), .O(n963)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_9 (.CI(n25166), .I0(n910), 
            .I1(VCC_net), .CO(n25167));
    SB_LUT4 encoder0_position_23__I_0_add_619_8_lut (.I0(GND_net), .I1(n911), 
            .I2(VCC_net), .I3(n25165), .O(n964)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_8 (.CI(n25165), .I0(n911), 
            .I1(VCC_net), .CO(n25166));
    SB_LUT4 encoder0_position_23__I_0_add_619_7_lut (.I0(GND_net), .I1(n912), 
            .I2(GND_net), .I3(n25164), .O(n965)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_7 (.CI(n25164), .I0(n912), 
            .I1(GND_net), .CO(n25165));
    SB_LUT4 encoder0_position_23__I_0_add_619_6_lut (.I0(GND_net), .I1(n913), 
            .I2(GND_net), .I3(n25163), .O(n966)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_6 (.CI(n25163), .I0(n913), 
            .I1(GND_net), .CO(n25164));
    SB_LUT4 encoder0_position_23__I_0_add_619_5_lut (.I0(GND_net), .I1(n914), 
            .I2(VCC_net), .I3(n25162), .O(n967)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_5 (.CI(n25162), .I0(n914), 
            .I1(VCC_net), .CO(n25163));
    SB_LUT4 encoder0_position_23__I_0_add_619_4_lut (.I0(GND_net), .I1(n915), 
            .I2(GND_net), .I3(n25161), .O(n968)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_4 (.CI(n25161), .I0(n915), 
            .I1(GND_net), .CO(n25162));
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4539), .I3(n25069), .O(displacement_23__N_50[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_619_3_lut (.I0(GND_net), .I1(n916), 
            .I2(VCC_net), .I3(n25160), .O(n969)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_3 (.CI(n25160), .I0(n916), 
            .I1(VCC_net), .CO(n25161));
    SB_LUT4 encoder0_position_23__I_0_add_619_2_lut (.I0(GND_net), .I1(n431), 
            .I2(GND_net), .I3(VCC_net), .O(n970)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n25069), .I0(encoder1_position[16]), 
            .I1(n9_adj_4539), .CO(n25070));
    SB_CARRY encoder0_position_23__I_0_add_619_2 (.CI(VCC_net), .I0(n431), 
            .I1(GND_net), .CO(n25160));
    SB_LUT4 encoder0_position_23__I_0_add_566_10_lut (.I0(GND_net), .I1(n830), 
            .I2(VCC_net), .I3(n25159), .O(n883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_566_9_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n25158), .O(n884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_CARRY encoder0_position_23__I_0_add_566_9 (.CI(n25158), .I0(n831), 
            .I1(VCC_net), .CO(n25159));
    SB_LUT4 encoder0_position_23__I_0_add_566_8_lut (.I0(GND_net), .I1(n832), 
            .I2(VCC_net), .I3(n25157), .O(n885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_8 (.CI(n25157), .I0(n832), 
            .I1(VCC_net), .CO(n25158));
    SB_LUT4 encoder0_position_23__I_0_add_566_7_lut (.I0(GND_net), .I1(n833), 
            .I2(GND_net), .I3(n25156), .O(n886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_7 (.CI(n25156), .I0(n833), 
            .I1(GND_net), .CO(n25157));
    SB_LUT4 encoder0_position_23__I_0_add_566_6_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(n25155), .O(n887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28281_3_lut (.I0(n33956), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n33957));   // verilog/pwm.v(21[8:24])
    defparam i28281_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i12789_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4216), .I3(GND_net), .O(n16898));   // verilog/coms.v(127[12] 300[6])
    defparam i12789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4605));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.data_o({quadA_debounced_adj_4504, 
            quadB_debounced_adj_4505}), .GND_net(GND_net), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n32056(n32056), .reg_B({reg_B_adj_4715}), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .VCC_net(VCC_net), .n16872(n16872), 
            .ENCODER1_B_c_0(ENCODER1_B_c_0), .n17382(n17382)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(194[15] 199[4])
    SB_LUT4 i28180_3_lut (.I0(n33957), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n33856));   // verilog/pwm.v(21[8:24])
    defparam i28180_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4604));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4603));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_558_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4571));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4573));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4577));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4576));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4575));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4569));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4579));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4580));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4578));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_558_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4582));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_558_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4584));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4585));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4581));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_558_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_41_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[0]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4602));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4539));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_41_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[1]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12819_3_lut (.I0(\data_in_frame[18] [7]), .I1(rx_data[7]), 
            .I2(n29535), .I3(GND_net), .O(n16928));   // verilog/coms.v(127[12] 300[6])
    defparam i12819_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12820_3_lut (.I0(\data_in_frame[18] [6]), .I1(rx_data[6]), 
            .I2(n29535), .I3(GND_net), .O(n16929));   // verilog/coms.v(127[12] 300[6])
    defparam i12820_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12821_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n29535), .I3(GND_net), .O(n16930));   // verilog/coms.v(127[12] 300[6])
    defparam i12821_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12822_3_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n29535), .I3(GND_net), .O(n16931));   // verilog/coms.v(127[12] 300[6])
    defparam i12822_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12823_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n29535), .I3(GND_net), .O(n16932));   // verilog/coms.v(127[12] 300[6])
    defparam i12823_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12824_3_lut (.I0(\data_in_frame[18] [2]), .I1(rx_data[2]), 
            .I2(n29535), .I3(GND_net), .O(n16933));   // verilog/coms.v(127[12] 300[6])
    defparam i12824_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12825_3_lut (.I0(\data_in_frame[18] [1]), .I1(rx_data[1]), 
            .I2(n29535), .I3(GND_net), .O(n16934));   // verilog/coms.v(127[12] 300[6])
    defparam i12825_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12826_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n29535), .I3(GND_net), .O(n16935));   // verilog/coms.v(127[12] 300[6])
    defparam i12826_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_41_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[2]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4601));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4600));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4599));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4598));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_41_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[3]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4597));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4538));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4537));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4596));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_41_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[4]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4595));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_41_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[5]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4594));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4593));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_41_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4529), .I3(n15_adj_4531), .O(motor_state_23__N_74[6]));   // verilog/TinyFPGA_B.v(167[5] 169[10])
    defparam mux_41_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4592));   // verilog/TinyFPGA_B.v(202[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4536));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    motorControl control (.\Kp[2] (Kp[2]), .GND_net(GND_net), .\Kp[0] (Kp[0]), 
            .\Kp[1] (Kp[1]), .\Kp[3] (Kp[3]), .\Kp[6] (Kp[6]), .\Kp[4] (Kp[4]), 
            .\Ki[8] (Ki[8]), .\Kp[5] (Kp[5]), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), 
            .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
            .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
            .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), 
            .\Ki[15] (Ki[15]), .PWMLimit({PWMLimit}), .IntegralLimit({IntegralLimit}), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), 
            .\Kp[15] (Kp[15]), .n29(n29), .\duty_23__N_3516[14] (duty_23__N_3516[14]), 
            .duty({duty}), .clk32MHz(clk32MHz), .setpoint({setpoint}), 
            .motor_state({motor_state}), .n34501(n34501), .VCC_net(VCC_net), 
            .n18701(n18701)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(171[16] 183[4])
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4528));   // verilog/TinyFPGA_B.v(203[21:65])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12843_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n29538), .I3(GND_net), .O(n16952));   // verilog/coms.v(127[12] 300[6])
    defparam i12843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12844_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n29538), .I3(GND_net), .O(n16953));   // verilog/coms.v(127[12] 300[6])
    defparam i12844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12845_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n29538), .I3(GND_net), .O(n16954));   // verilog/coms.v(127[12] 300[6])
    defparam i12845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12846_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n29538), .I3(GND_net), .O(n16955));   // verilog/coms.v(127[12] 300[6])
    defparam i12846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12847_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n29538), .I3(GND_net), .O(n16956));   // verilog/coms.v(127[12] 300[6])
    defparam i12847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12848_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n29538), .I3(GND_net), .O(n16957));   // verilog/coms.v(127[12] 300[6])
    defparam i12848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12849_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n29538), .I3(GND_net), .O(n16958));   // verilog/coms.v(127[12] 300[6])
    defparam i12849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12850_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n29538), .I3(GND_net), .O(n16959));   // verilog/coms.v(127[12] 300[6])
    defparam i12850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_4652), .I3(control_mode[2]), .O(n15450));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12851_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n29541), .I3(GND_net), .O(n16960));   // verilog/coms.v(127[12] 300[6])
    defparam i12851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12852_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n29541), .I3(GND_net), .O(n16961));   // verilog/coms.v(127[12] 300[6])
    defparam i12852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12853_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n29541), .I3(GND_net), .O(n16962));   // verilog/coms.v(127[12] 300[6])
    defparam i12853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12854_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n29541), .I3(GND_net), .O(n16963));   // verilog/coms.v(127[12] 300[6])
    defparam i12854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12855_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n29541), .I3(GND_net), .O(n16964));   // verilog/coms.v(127[12] 300[6])
    defparam i12855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12856_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n29541), .I3(GND_net), .O(n16965));   // verilog/coms.v(127[12] 300[6])
    defparam i12856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12857_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n29541), .I3(GND_net), .O(n16966));   // verilog/coms.v(127[12] 300[6])
    defparam i12857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12858_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n29541), .I3(GND_net), .O(n16967));   // verilog/coms.v(127[12] 300[6])
    defparam i12858_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .GND_net(GND_net), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .setpoint({setpoint}), 
         .clk32MHz(clk32MHz), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n63(n63_adj_4566), .n771(n771), .n63_adj_3(n63), .\FRAME_MATCHER.i_31__N_2364 (\FRAME_MATCHER.i_31__N_2364 ), 
         .n29497(n29497), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .n12869(n12869), .n2329(n2329), .n4452(n4452), .\data_in[0] ({\data_in[0] }), 
         .\data_in[2] ({\data_in[2] }), .\data_in[3] ({\data_in[3] }), .\data_in[1] ({\data_in[1] }), 
         .\FRAME_MATCHER.i_31__N_2370 (\FRAME_MATCHER.i_31__N_2370 ), .PWMLimit({PWMLimit}), 
         .\duty_23__N_3516[14] (duty_23__N_3516[14]), .n29(n29), .rx_data({rx_data}), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_in_frame[18] ({\data_in_frame[18] }), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .tx_active(tx_active), 
         .\FRAME_MATCHER.state[2] (\FRAME_MATCHER.state [2]), .rx_data_ready(rx_data_ready), 
         .n16911(n16911), .\data_in_frame[21] ({\data_in_frame[21] }), .n16910(n16910), 
         .n16909(n16909), .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n4218(n4218), .n16908(n16908), .n16907(n16907), .\data_in_frame[9] ({\data_in_frame[9] [7], 
         Open_0, Open_1, Open_2, Open_3, Open_4, Open_5, Open_6}), 
         .\data_in_frame[9][5] (\data_in_frame[9] [5]), .\data_in_frame[9][4] (\data_in_frame[9] [4]), 
         .\data_in_frame[9][3] (\data_in_frame[9] [3]), .\data_in_frame[9][2] (\data_in_frame[9] [2]), 
         .\data_in_frame[9][1] (\data_in_frame[9] [1]), .\data_in_frame[9][0] (\data_in_frame[9] [0]), 
         .n16906(n16906), .n78(n78), .n16905(n16905), .n16904(n16904), 
         .n16903(n16903), .control_mode({control_mode}), .n16902(n16902), 
         .\data_in_frame[10] ({\data_in_frame[10] [7:3], Open_7, Open_8, 
         Open_9}), .\data_in_frame[5] ({\data_in_frame[5] }), .n16901(n16901), 
         .\data_in_frame[15] ({\data_in_frame[15] }), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[14] ({\data_in_frame[14] }), 
         .n16900(n16900), .n16899(n16899), .n12944(n12944), .\data_in_frame[10][1] (\data_in_frame[10] [1]), 
         .n2(n2_adj_4638), .DE_c(DE_c), .n8868(n8868), .n16898(n16898), 
         .n16897(n16897), .n16896(n16896), .n16894(n16894), .n16893(n16893), 
         .n16892(n16892), .n16891(n16891), .n16890(n16890), .n16889(n16889), 
         .n16888(n16888), .n16887(n16887), .n16886(n16886), .n16885(n16885), 
         .n16884(n16884), .n16882(n16882), .n16881(n16881), .n16880(n16880), 
         .n16879(n16879), .n16878(n16878), .n16877(n16877), .n16876(n16876), 
         .n16875(n16875), .n16874(n16874), .n35073(n35073), .n28937(n28937), 
         .n16867(n16867), .VCC_net(VCC_net), .n17373(n17373), .IntegralLimit({IntegralLimit}), 
         .n17372(n17372), .n17371(n17371), .n17370(n17370), .n17369(n17369), 
         .n17368(n17368), .n17367(n17367), .n17335(n17335), .n17334(n17334), 
         .n17333(n17333), .n17332(n17332), .n17331(n17331), .n17330(n17330), 
         .n17329(n17329), .n17328(n17328), .n17327(n17327), .n17326(n17326), 
         .n17325(n17325), .n17324(n17324), .n17323(n17323), .n17322(n17322), 
         .n17321(n17321), .n17320(n17320), .n17314(n17314), .n17313(n17313), 
         .n17312(n17312), .n17311(n17311), .n17310(n17310), .n17309(n17309), 
         .n17308(n17308), .n17307(n17307), .n17306(n17306), .n17305(n17305), 
         .n17304(n17304), .n17303(n17303), .n17302(n17302), .n17301(n17301), 
         .n17300(n17300), .n17299(n17299), .n17298(n17298), .n17297(n17297), 
         .n17296(n17296), .n17295(n17295), .n17294(n17294), .n17293(n17293), 
         .n17292(n17292), .n17291(n17291), .n17290(n17290), .n17289(n17289), 
         .n17288(n17288), .n17287(n17287), .n17286(n17286), .n17285(n17285), 
         .n17284(n17284), .n17283(n17283), .\Kp[1] (Kp[1]), .n17282(n17282), 
         .\Kp[2] (Kp[2]), .n17281(n17281), .\Kp[3] (Kp[3]), .n17280(n17280), 
         .\Kp[4] (Kp[4]), .n17279(n17279), .\Kp[5] (Kp[5]), .n17278(n17278), 
         .\Kp[6] (Kp[6]), .n17277(n17277), .\Kp[7] (Kp[7]), .n17276(n17276), 
         .\Kp[8] (Kp[8]), .n17275(n17275), .\Kp[9] (Kp[9]), .n17274(n17274), 
         .\Kp[10] (Kp[10]), .n17273(n17273), .\Kp[11] (Kp[11]), .n17272(n17272), 
         .\Kp[12] (Kp[12]), .n17271(n17271), .\Kp[13] (Kp[13]), .n17270(n17270), 
         .\Kp[14] (Kp[14]), .n17269(n17269), .\Kp[15] (Kp[15]), .n17268(n17268), 
         .\Ki[1] (Ki[1]), .n17267(n17267), .\Ki[2] (Ki[2]), .n17266(n17266), 
         .\Ki[3] (Ki[3]), .n17265(n17265), .\Ki[4] (Ki[4]), .n17264(n17264), 
         .\Ki[5] (Ki[5]), .n17263(n17263), .\Ki[6] (Ki[6]), .n17262(n17262), 
         .\Ki[7] (Ki[7]), .n17261(n17261), .\Ki[8] (Ki[8]), .n17260(n17260), 
         .\Ki[9] (Ki[9]), .n17259(n17259), .\Ki[10] (Ki[10]), .n17258(n17258), 
         .\Ki[11] (Ki[11]), .n17257(n17257), .\Ki[12] (Ki[12]), .n17256(n17256), 
         .\Ki[13] (Ki[13]), .n17255(n17255), .\Ki[14] (Ki[14]), .n17254(n17254), 
         .\Ki[15] (Ki[15]), .n17253(n17253), .n17252(n17252), .n17251(n17251), 
         .n17250(n17250), .n17249(n17249), .n17248(n17248), .n17247(n17247), 
         .n17246(n17246), .n17245(n17245), .n17244(n17244), .n17243(n17243), 
         .n17242(n17242), .n17241(n17241), .n17240(n17240), .n17239(n17239), 
         .n17238(n17238), .n17237(n17237), .n17236(n17236), .n17235(n17235), 
         .n17234(n17234), .n17233(n17233), .n17232(n17232), .n4216(n4216), 
         .n122(n122), .n5(n5_adj_4590), .n35368(n35368), .n17231(n17231), 
         .n17230(n17230), .n17229(n17229), .n17228(n17228), .n17227(n17227), 
         .n17226(n17226), .n17225(n17225), .n17224(n17224), .n17223(n17223), 
         .n17222(n17222), .n17221(n17221), .n17220(n17220), .n17219(n17219), 
         .n17218(n17218), .n17217(n17217), .n17216(n17216), .n17215(n17215), 
         .n17214(n17214), .n17213(n17213), .n17212(n17212), .n17211(n17211), 
         .n17210(n17210), .n17209(n17209), .n17208(n17208), .n17207(n17207), 
         .n17206(n17206), .n17205(n17205), .n17204(n17204), .n17203(n17203), 
         .n17202(n17202), .n17201(n17201), .n17200(n17200), .n17199(n17199), 
         .n17198(n17198), .n17197(n17197), .n17196(n17196), .n17195(n17195), 
         .n17194(n17194), .n17193(n17193), .n17192(n17192), .n17191(n17191), 
         .n17190(n17190), .n17189(n17189), .n17188(n17188), .n17187(n17187), 
         .n17186(n17186), .n17185(n17185), .n17184(n17184), .n17183(n17183), 
         .n17182(n17182), .n17181(n17181), .n17180(n17180), .n17179(n17179), 
         .n17178(n17178), .n17177(n17177), .n17176(n17176), .n17175(n17175), 
         .n17174(n17174), .n17173(n17173), .n17172(n17172), .n17171(n17171), 
         .n17170(n17170), .n17169(n17169), .n17168(n17168), .n17167(n17167), 
         .n17166(n17166), .n17165(n17165), .n17164(n17164), .n17163(n17163), 
         .n17162(n17162), .n17161(n17161), .n17160(n17160), .n17159(n17159), 
         .n17158(n17158), .n17157(n17157), .n17156(n17156), .n17155(n17155), 
         .n17154(n17154), .n17153(n17153), .n17152(n17152), .n17151(n17151), 
         .n17150(n17150), .n17149(n17149), .n17148(n17148), .n17147(n17147), 
         .n17146(n17146), .n17145(n17145), .n17144(n17144), .n17143(n17143), 
         .n17142(n17142), .n17141(n17141), .n17140(n17140), .n17139(n17139), 
         .n17138(n17138), .n17137(n17137), .n17136(n17136), .n17135(n17135), 
         .n17134(n17134), .n17133(n17133), .n17132(n17132), .n17131(n17131), 
         .n17130(n17130), .n17129(n17129), .n17128(n17128), .n17127(n17127), 
         .n17126(n17126), .n17125(n17125), .n17124(n17124), .n17123(n17123), 
         .n17122(n17122), .n17121(n17121), .n17120(n17120), .n17119(n17119), 
         .n17118(n17118), .n17117(n17117), .n17116(n17116), .n29535(n29535), 
         .n17115(n17115), .n17114(n17114), .n17113(n17113), .n17112(n17112), 
         .n17111(n17111), .LED_c(LED_c), .n17110(n17110), .n29532(n29532), 
         .n17109(n17109), .n17108(n17108), .n17107(n17107), .n17106(n17106), 
         .n17105(n17105), .n17104(n17104), .n17103(n17103), .n17102(n17102), 
         .n17101(n17101), .neopxl_color({neopxl_color}), .n17100(n17100), 
         .n17099(n17099), .n17098(n17098), .n17097(n17097), .n17096(n17096), 
         .n17095(n17095), .n17094(n17094), .n17093(n17093), .n17092(n17092), 
         .n17091(n17091), .n17090(n17090), .n17089(n17089), .n17088(n17088), 
         .n17087(n17087), .n17086(n17086), .n17085(n17085), .n17084(n17084), 
         .n17083(n17083), .n17082(n17082), .n17081(n17081), .n17080(n17080), 
         .n17079(n17079), .n16865(n16865), .n16864(n16864), .\Ki[0] (Ki[0]), 
         .n16863(n16863), .\Kp[0] (Kp[0]), .n16862(n16862), .n16853(n16853), 
         .n17031(n17031), .n17030(n17030), .n17029(n17029), .n17028(n17028), 
         .n17027(n17027), .n17026(n17026), .n17025(n17025), .n17024(n17024), 
         .n17023(n17023), .n17022(n17022), .n17021(n17021), .n17020(n17020), 
         .n17019(n17019), .n17018(n17018), .n17017(n17017), .n17016(n17016), 
         .n16967(n16967), .n16966(n16966), .n16965(n16965), .n16964(n16964), 
         .n16963(n16963), .n16962(n16962), .n16961(n16961), .n16960(n16960), 
         .n16959(n16959), .n16958(n16958), .n16957(n16957), .n16956(n16956), 
         .n16955(n16955), .n16954(n16954), .n16953(n16953), .n16952(n16952), 
         .n16935(n16935), .n16934(n16934), .n16933(n16933), .n16932(n16932), 
         .n16931(n16931), .n16930(n16930), .n16929(n16929), .n16928(n16928), 
         .n18701(n18701), .n29541(n29541), .n29542(n29542), .n29538(n29538), 
         .n29539(n29539), .n6(n6_adj_4624), .\r_SM_Main[1] (r_SM_Main_adj_4704[1]), 
         .tx_o(tx_o), .n4(n4_adj_4494), .n16871(n16871), .n8947(n8947), 
         .tx_enable(tx_enable), .n16710(n16710), .n16802(n16802), .n21215(n21215), 
         .n4_adj_4(n4), .r_Rx_Data(r_Rx_Data), .n4_adj_5(n4_adj_4535), 
         .\r_Bit_Index[0] (r_Bit_Index[0]), .n15595(n15595), .RX_N_2(RX_N_2), 
         .n15590(n15590), .n4_adj_6(n4_adj_4530), .n17376(n17376), .n17380(n17380), 
         .n16861(n16861), .n16860(n16860), .n16859(n16859), .n16858(n16858), 
         .n16857(n16857), .n16856(n16856), .n16855(n16855)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(138[8] 161[4])
    pwm PWM (.n33856(n33856), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n15455(n15455), .pwm_counter({pwm_counter}), .GND_net(GND_net), 
        .n15453(n15453)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(90[6] 95[3])
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, GND_net, data_o, 
            clk32MHz, n31883, reg_B, VCC_net, n16870, ENCODER0_B_c_0, 
            n17381, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input GND_net;
    output [1:0]data_o;
    input clk32MHz;
    output n31883;
    output [1:0]reg_B;
    input VCC_net;
    input n16870;
    input ENCODER0_B_c_0;
    input n17381;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2549;
    
    wire n2545, n24956, n24957, n24955, A_delayed, B_delayed, count_enable, 
        n24954, n24953, count_direction, n24952, n24975, n24974, 
        n24973, n24972, n24971, n24970, n24969, n24968, n24967, 
        n24966, n24965, n24964, n24963, n24962, n24961, n24960, 
        n24959, n24958;
    
    SB_LUT4 add_555_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2545), 
            .I3(n24956), .O(n2549[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_6 (.CI(n24956), .I0(encoder0_position[4]), .I1(n2545), 
            .CO(n24957));
    SB_LUT4 add_555_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2545), 
            .I3(n24955), .O(n2549[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_5 (.CI(n24955), .I0(encoder0_position[3]), .I1(n2545), 
            .CO(n24956));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_555_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2545), 
            .I3(n24954), .O(n2549[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_4 (.CI(n24954), .I0(encoder0_position[2]), .I1(n2545), 
            .CO(n24955));
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2549[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_555_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2545), 
            .I3(n24953), .O(n2549[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_3 (.CI(n24953), .I0(encoder0_position[1]), .I1(n2545), 
            .CO(n24954));
    SB_LUT4 add_555_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n24952), .O(n2549[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_2 (.CI(n24952), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n24953));
    SB_CARRY add_555_1 (.CI(GND_net), .I0(n2545), .I1(n2545), .CO(n24952));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_555_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2545), 
            .I3(n24975), .O(n2549[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2545), 
            .I3(n24974), .O(n2549[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_24 (.CI(n24974), .I0(encoder0_position[22]), .I1(n2545), 
            .CO(n24975));
    SB_LUT4 add_555_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2545), 
            .I3(n24973), .O(n2549[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_23 (.CI(n24973), .I0(encoder0_position[21]), .I1(n2545), 
            .CO(n24974));
    SB_LUT4 add_555_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2545), 
            .I3(n24972), .O(n2549[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_22 (.CI(n24972), .I0(encoder0_position[20]), .I1(n2545), 
            .CO(n24973));
    SB_LUT4 add_555_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2545), 
            .I3(n24971), .O(n2549[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_21 (.CI(n24971), .I0(encoder0_position[19]), .I1(n2545), 
            .CO(n24972));
    SB_LUT4 add_555_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2545), 
            .I3(n24970), .O(n2549[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_20 (.CI(n24970), .I0(encoder0_position[18]), .I1(n2545), 
            .CO(n24971));
    SB_LUT4 add_555_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2545), 
            .I3(n24969), .O(n2549[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_19 (.CI(n24969), .I0(encoder0_position[17]), .I1(n2545), 
            .CO(n24970));
    SB_LUT4 add_555_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2545), 
            .I3(n24968), .O(n2549[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_18 (.CI(n24968), .I0(encoder0_position[16]), .I1(n2545), 
            .CO(n24969));
    SB_LUT4 add_555_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2545), 
            .I3(n24967), .O(n2549[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_17 (.CI(n24967), .I0(encoder0_position[15]), .I1(n2545), 
            .CO(n24968));
    SB_LUT4 add_555_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2545), 
            .I3(n24966), .O(n2549[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_16 (.CI(n24966), .I0(encoder0_position[14]), .I1(n2545), 
            .CO(n24967));
    SB_LUT4 add_555_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2545), 
            .I3(n24965), .O(n2549[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_15 (.CI(n24965), .I0(encoder0_position[13]), .I1(n2545), 
            .CO(n24966));
    SB_LUT4 add_555_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2545), 
            .I3(n24964), .O(n2549[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_14 (.CI(n24964), .I0(encoder0_position[12]), .I1(n2545), 
            .CO(n24965));
    SB_LUT4 add_555_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2545), 
            .I3(n24963), .O(n2549[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_13 (.CI(n24963), .I0(encoder0_position[11]), .I1(n2545), 
            .CO(n24964));
    SB_LUT4 add_555_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2545), 
            .I3(n24962), .O(n2549[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_12 (.CI(n24962), .I0(encoder0_position[10]), .I1(n2545), 
            .CO(n24963));
    SB_LUT4 add_555_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2545), 
            .I3(n24961), .O(n2549[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_11 (.CI(n24961), .I0(encoder0_position[9]), .I1(n2545), 
            .CO(n24962));
    SB_LUT4 add_555_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2545), 
            .I3(n24960), .O(n2549[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_10 (.CI(n24960), .I0(encoder0_position[8]), .I1(n2545), 
            .CO(n24961));
    SB_LUT4 add_555_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2545), 
            .I3(n24959), .O(n2549[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_9 (.CI(n24959), .I0(encoder0_position[7]), .I1(n2545), 
            .CO(n24960));
    SB_LUT4 add_555_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2545), 
            .I3(n24958), .O(n2549[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_8 (.CI(n24958), .I0(encoder0_position[6]), .I1(n2545), 
            .CO(n24959));
    SB_LUT4 add_555_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2545), 
            .I3(n24957), .O(n2549[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_7 (.CI(n24957), .I0(encoder0_position[5]), .I1(n2545), 
            .CO(n24958));
    SB_LUT4 i846_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2545));   // quad.v(37[5] 40[8])
    defparam i846_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,100)_U0  debounce (.n31883(n31883), .reg_B({reg_B}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .n16870(n16870), .data_o({data_o}), .ENCODER0_B_c_0(ENCODER0_B_c_0), 
            .n17381(n17381), .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (n31883, reg_B, GND_net, clk32MHz, 
            VCC_net, n16870, data_o, ENCODER0_B_c_0, n17381, ENCODER0_A_c_1);
    output n31883;
    output [1:0]reg_B;
    input GND_net;
    input clk32MHz;
    input VCC_net;
    input n16870;
    output [1:0]data_o;
    input ENCODER0_B_c_0;
    input n17381;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3600;
    wire [6:0]n33;
    
    wire n25582, n25581, n25580, n25579, n25578, n25577;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[3]), .I1(cnt_reg[5]), .I2(cnt_reg[1]), 
            .I3(cnt_reg[0]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[6]), .I1(n12), .I2(cnt_reg[2]), .I3(cnt_reg[4]), 
            .O(n31883));
    defparam i6_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n31883), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1131_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n25582), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1131_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1131_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n25581), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1131_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1131_add_4_7 (.CI(n25581), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n25582));
    SB_LUT4 cnt_reg_1131_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n25580), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1131_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1131_add_4_6 (.CI(n25580), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n25581));
    SB_LUT4 cnt_reg_1131_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n25579), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1131_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1131_add_4_5 (.CI(n25579), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n25580));
    SB_LUT4 cnt_reg_1131_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n25578), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1131_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1131_add_4_4 (.CI(n25578), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n25579));
    SB_LUT4 cnt_reg_1131_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n25577), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1131_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1131_add_4_3 (.CI(n25577), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n25578));
    SB_LUT4 cnt_reg_1131_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1131_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1131_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n25577));
    SB_DFFSR cnt_reg_1131__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n16870));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n17381));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1131__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1131__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1131__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1131__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1131__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1131__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (\neo_pixel_transmitter.done , clk32MHz, GND_net, VCC_net, 
            timer, \neo_pixel_transmitter.t0 , \state_3__N_272[1] , start, 
            LED_c, \state[0] , n21971, \state[1] , n22115, neopxl_color, 
            n16698, n30267, n28583, n28495, n17366, n17365, n17364, 
            n17363, n17362, n17361, n17360, n17359, n17358, n17357, 
            n17356, n17355, n17354, n17353, n17352, n17351, n17350, 
            n17349, n17348, n17347, n17346, n17345, n17344, n17343, 
            n17342, n17341, n17340, n17339, n17338, n17337, n17336, 
            n17316, NEOPXL_c, n16852) /* synthesis syn_module_defined=1 */ ;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    input GND_net;
    input VCC_net;
    output [31:0]timer;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output \state_3__N_272[1] ;
    output start;
    input LED_c;
    output \state[0] ;
    output n21971;
    output \state[1] ;
    output n22115;
    input [23:0]neopxl_color;
    output n16698;
    output n30267;
    output n28583;
    input n28495;
    input n17366;
    input n17365;
    input n17364;
    input n17363;
    input n17362;
    input n17361;
    input n17360;
    input n17359;
    input n17358;
    input n17357;
    input n17356;
    input n17355;
    input n17354;
    input n17353;
    input n17352;
    input n17351;
    input n17350;
    input n17349;
    input n17348;
    input n17347;
    input n17346;
    input n17345;
    input n17344;
    input n17343;
    input n17342;
    input n17341;
    input n17340;
    input n17339;
    input n17338;
    input n17337;
    input n17336;
    input n17316;
    output NEOPXL_c;
    input n16852;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n44, \neo_pixel_transmitter.done_N_480 , n34806, n2498, n2399, 
        n2423, n25696, n25697, n2499, n2400, n25695, n2500, n2401, 
        n25694, n2501, n2402, n25693, n2502, n2403, n25692, n2503, 
        n2404, n25691, n2504, n2405, n25690, n2505, n2406, n25689;
    wire [31:0]n255;
    
    wire n16688, n16807, n1409, n21925, n1405, n1403, n1406, n16, 
        n1402, n1404, n1400, n1407, n17, n1408, n1401, n1433, 
        n1037, n34504, n2;
    wire [31:0]n971;
    
    wire n1007, n1006, n906, n1005, n905, n30427, n32222, n1304, 
        n1305, n10, n1303, n1309, n12, n1306, n1308, n1302, 
        n16_adj_4339, n1307, n1301, n1334, n16727, n14162, n1009, 
        n1008, n32274, n6, n4, n2506, n2407, n25688, n2507, 
        n2408, n25687, n2508, n2409, n34489, n25686, n2194, n2095, 
        n2126, n25781, n25782, n2324, n34500, n2509, n2588, n2489, 
        n2522, n25685, n2589, n2490, n25684, n1235, n34497, n30, 
        n43, n2195, n2096, n25780, n3116, n34503, n2590, n2491, 
        n25683;
    wire [31:0]one_wire_N_423;
    wire [31:0]n1;
    
    wire n25004, n2196, n2097, n25779, n25005, n2197, n2098, n25778, 
        n2591, n2492, n25682, n2592, n2493, n25681, n2593, n2494, 
        n25680, n2594, n2495, n25679, n2198, n2099, n25777, n2595, 
        n2496, n25678, n2596, n2497, n25677, n2597, n25676, n24812, 
        n2199, n2100, n25776, n2598, n25675, n2599, n25674, n2600, 
        n25673, n2601, n25672, n3102, n3090, n3103, n3085, n42, 
        n3089, n3094, n3101, n3098, n46, n3099, n3091, n3106, 
        n3100, n44_adj_4340, n3097, n3088, n3104, n3092, n45, 
        n3105, n3083, n3093, n3096, n43_adj_4341, n3108, n3109, 
        n40, n2602, n25671, n2603, n25670, n3107, n3087, n3086, 
        n48, n2604, n25669, n52, n3095, n3084, n39, n1205, n1206, 
        n1204, n1207, n14, n1203, n1209, n9, n1202, n1208, n1136, 
        n34495, n2605, n25668, n3017, n34502, n45_adj_4342, n47, 
        n46_adj_4343, n48_adj_4344, n54, n1109, n21895, n1105, n1103, 
        n1108, n12_adj_4345, n1107, n1106, n1104, n2206, n2204, 
        n28_adj_4346, n2209, n21889, n2193, n32_adj_4347, n2208, 
        n2192, n2205, n2201, n30_adj_4348, n2207, n31_adj_4349, 
        n2202, n2200, n2203, n29, n2225, n2819, n34494, n2606, 
        n25667, n34490, n2798, n2804, n2791, n2795, n40_adj_4350, 
        n2796, n2793, n2788, n2808, n38, n2789, n2800, n2803, 
        n2805, n39_adj_4351, n2792, n2787, n2801, n2799, n37, 
        n2786, n2797, n34, n2794, n2806, n2807, n2790, n42_adj_4352, 
        n46_adj_4353, n2802, n2809, n33_adj_4354, n2720, n34493, 
        n2607, n25666, n2608, n34491, n25665, n2609, n2687, n2621, 
        n25664, n2688, n25663, n2101, n25775, n2689, n25662, n2690, 
        n25661, n2691, n25660, n2692, n25659, n2693, n25658, n2694, 
        n25657, n49, n2695, n25656, n2696, n25655, n2697, n25654, 
        n2704, n28_adj_4357, n2699, n2706, n38_adj_4358, n2709, 
        n21903, n2701, n36, n2700, n2705, n42_adj_4359, n2702, 
        n2708, n40_adj_4360, n2703, n41, n2698, n2707, n39_adj_4361, 
        n34492, n36_adj_4362, n25, n34_adj_4363, n40_adj_4364, n38_adj_4365, 
        n39_adj_4366, n37_adj_4367, n2102, n25774, n25653, n2103, 
        n25773, n25652, n25651, n25650, n25649, n25648, n25647, 
        n25646, n25645, n25644, n25643, n25642, n25641, n25640, 
        n25639, n26419, n25638, n25637, n25636, n2104, n25772, 
        n25635, n25003, n25634, n25633, n25632, n25631, n25630, 
        n25629, n2105, n25771, n25628, n25627, n25002, n25626, 
        n25625, n24820, n2106, n25770, n25624, n25623, n15574, 
        n26673, n30348, n15581, n14_adj_4368, n9_adj_4369, n15471, 
        n2107, n25769, n25622, n25621, n25620, n2108, n25768, 
        n831, n2885, n25619, n2886, n25618, n2887, n25617, n2888, 
        n25616, n2889, n25615, n2890, n25614, n2109, n25767, n2891, 
        n25613, n2892, n25612, n2893, n25611, n2894, n25610, n2895, 
        n25609, n2896, n25608, n2897, n25607, n2898, n25606, n2899, 
        n25605, n2900, n25604, n2901, n25603, n2902, n25602, n33493, 
        n33192, n30455, n33494, n30475, \neo_pixel_transmitter.done_N_486 , 
        n2903, n25601, n2904, n25600, n2905, n25599, n2906, n25598, 
        n2907, n25597, n2908, n25596, n2909, n2291, n25766, n25595, 
        n25594, n25593, n2292, n25765, n25592, n25591, n24, n34_adj_4373, 
        n22, n38_adj_4374, n36_adj_4375, n37_adj_4376, n35, n25590, 
        n22039, n25001, n25589, n25144, n25143, n2293, n25764, 
        n25142, n25141, n25000, n4_adj_4377, n3209, n21917, n35_adj_4378, 
        n11, n29_adj_4379, n51, n48_adj_4380, n37_adj_4381, n23, 
        n53, n39_adj_4382, n46_adj_4383, n27, n57, n63, n43_adj_4384, 
        n47_adj_4385, n25_adj_4386, n33_adj_4387, n47_adj_4388, n61, 
        n45_adj_4389, n59, n17_adj_4390, n15_adj_4391, n55, n44_adj_4392, 
        n31_adj_4393, n41_adj_4394, n49_adj_4395, n43_adj_4396, n54_adj_4397, 
        n45_adj_4398, n13_adj_4399, n19_adj_4400, n21_adj_4401, n49_adj_4402, 
        n26709, n35413, n25140;
    wire [4:0]color_bit_N_466;
    
    wire n34714, n34612, n33147, n2294, n25763, n25139, n34528;
    wire [3:0]state_3__N_272;
    
    wire n2295, n25762, n25138, n25137, n4081, n2296, n25761, 
        n18_adj_4404, n21887, n2093, n30_adj_4405, n2094, n28_adj_4406, 
        n29_adj_4407, n27_adj_4408, n2297, n25760, n25136, n2298, 
        n25759, n2299, n25758, n2300, n25757, n25135, n33174, 
        n2301, n25756, n25134, n25133, n25132;
    wire [31:0]n133;
    
    wire n25530, n25529, n25528, n25527, n25131, n2302, n25755, 
        n25526, n25525, n25524, n2303, n25754, n25523, n25522, 
        n25521, n25520, n25519, n25518, n25130, n3004, n2989, 
        n2990, n3007, n40_adj_4409, n3006, n2984, n2988, n2986, 
        n44_adj_4410, n3008, n3003, n2994, n3002, n42_adj_4411, 
        n2999, n3000, n2992, n2997, n43_adj_4412, n2996, n2985, 
        n2995, n2987, n41_adj_4413, n3001, n2993, n38_adj_4414, 
        n2998, n2991, n46_adj_4415, n50, n3005, n3009, n37_adj_4416, 
        n2918, n34499, n25517, n25516, n25515, n24813, n25129, 
        n25514, n2304, n25753, n25513, n25512, n25511, n25510, 
        n25509, n25508, n25507, n34498, n25128, n25506, n25505, 
        n25504, n2305, n25752, n25503, n25502, n25501, n25500, 
        n25499, n25498, n24821, n25497, n25496, n25495, n25494, 
        n25493, n25492, n25491, n24840, n25127, n25490, n24839, 
        n25489, n25126, n25488, n24838, n2306, n25751, n25125, 
        n25487, n25124, n2307, n25750, n25486, n25123, n25485, 
        n25484, n2308, n34496, n25749, n2309, n22_adj_4417, n2390, 
        n25748, n30_adj_4418, n2391, n25747, n34_adj_4419, n2392, 
        n25746, n2393, n25745, n25483, n32_adj_4420, n33_adj_4421, 
        n25482, n25481, n25480, n25479, n25478, n2394, n25744, 
        n25477, n24837, n2395, n25743, n2396, n25742, n2397, n25741, 
        n25476, n31_adj_4422, n24836, n25475, n24835, n2398, n25740, 
        n25474, n25473, n25739, n838, n25472, n807, n60, n25738, 
        n25471, n608, n708, n21867, n6706, n30429, n14164, n33_adj_4423, 
        n41_adj_4424, n38_adj_4425, n43_adj_4426, n40_adj_4427, n46_adj_4428, 
        n25470, n39_adj_4429, n47_adj_4430, n25469, n25468, n25467, 
        n25466, n25465, n25737, n25464, n25463, n25462, n25461, 
        n25460, n25459, n25458, n24834, n25457, n25456, n25455, 
        n25454, n25453, n25452, n25451, n25736, n25450, n25449, 
        n25735, n25448, n25734, n25447, n25733, n25732, n25446, 
        n25445, n25444, n25443, n25442, n25441, n25440, n25439, 
        n25438, n25437, n25436, n25435, n25434, n25433, n25432, 
        n25431, n25430, n25429, n25731, n25428, n25427, n25426, 
        n25425, n25424, n25423, n25422, n24819, n25730, n30302, 
        n33100, n30261, n27_adj_4431, n33_adj_4432, n34711, n32_adj_4433, 
        n31_adj_4434, n845, n35_adj_4435, n37_adj_4436, n21_adj_4437, 
        n23_adj_4438, n22_adj_4439, n24_adj_4440, n36_adj_4441, n25_adj_4442, 
        n27_adj_4443, n26, n28_adj_4444, n37_adj_4445, n29_adj_4446, 
        n30_adj_4447, n34675, n32383, n30350, n29563, n111, n34663, 
        n32389, n34609, n34597, n33801, n24833, n24832, n25030, 
        n25029, n25028, n24811, n25027, n25026, n24818, n25025, 
        n116, n16_adj_4451, n24831, n25024, n24817, n25023, n24810, 
        n24830, n24816, n24829, n24828, n25022, n30370, n7_adj_4454, 
        n22071, n25021, n18_adj_4456, n25705, n25704, n25020, n25703, 
        n24827, n25702, n25701, n25700, n25699, n25698, n25019, 
        n25018, n25017, n25016, n32089, n25015, n24826, n25014, 
        n25013, n25012, n25011, n25880, n25879, n25878, n25877, 
        n25876, n25875, n1499, n25874, n1500, n25873, n1501, n25872, 
        n1502, n25871, n1503, n25870, n1504, n25869, n1505, n25868, 
        n1506, n25867, n1507, n25866, n1508, n34505, n25865, n1509, 
        n1598, n1532, n25864, n1599, n25863, n1600, n25862, n1601, 
        n25861, n1602, n25860, n24825, n1603, n25859, n1604, n25858, 
        n25010, n1605, n25857, n1606, n25856, n1607, n25855, n1608, 
        n34506, n25854, n1609, n1697, n1631, n25853, n1698, n25852, 
        n1699, n25851, n1700, n25850, n1701, n25849, n1702, n25848, 
        n25009, n1703, n25847, n1704, n25846, n1705, n25845, n1706, 
        n25844, n1707, n25843, n1708, n34507, n25842, n24824, 
        n1709, n1796, n1730, n25841, n1797, n25840, n1798, n25839, 
        n24815, n1799, n25838, n1800, n25837, n1801, n25836, n1802, 
        n25835, n1803, n25834, n1804, n25833, n25008, n1805, n25832, 
        n1806, n25831, n1807, n25830, n1808, n34508, n25829, n25007, 
        n1809, n1895, n1829, n25828, n1896, n25827, n1897, n25826, 
        n25006, n1898, n25825, n24823, n1899, n25824, n1900, n25823, 
        n1901, n25822, n1902, n25821, n1903, n25820, n1904, n25819, 
        n1905, n25818, n1906, n25817, n1907, n25816, n24814, n1908, 
        n34509, n25815, n1909, n1994, n1928, n25814, n1995, n25813, 
        n1996, n25812, n24822, n1997, n25811, n1998, n25810, n1999, 
        n25809, n2000, n25808, n2001, n25807, n2002, n25806, n2003, 
        n25805, n2004, n25804, n2005, n25803, n2006, n25802, n2007, 
        n25801, n2008, n34510, n25800, n2009, n2027, n25799, n25798, 
        n25797, n25796, n25795, n25794, n25793, n25792, n25791, 
        n25790, n25789, n25788, n25787, n25786, n25785, n34511, 
        n25784, n25783, n34516, n34525, n34513, n18_adj_4463, n28_adj_4464, 
        n26_adj_4465, n27_adj_4466, n25_adj_4467, n26_adj_4468, n19_adj_4469, 
        n16_adj_4470, n24_adj_4471, n28_adj_4472, n24_adj_4473, n22_adj_4474, 
        n23_adj_4475, n21_adj_4476, n17_adj_4477, n21_adj_4478, n20_adj_4479, 
        n24_adj_4480, n20_adj_4481, n13_adj_4482, n18_adj_4483, n22_adj_4484, 
        n18_adj_4485, n20_adj_4486, n15_adj_4487;
    
    SB_LUT4 i16_4_lut (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n34806), .D(\neo_pixel_transmitter.done_N_480 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n25696), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n25696), .I0(n2399), .I1(n2423), .CO(n25697));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n25695), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n25695), .I0(n2400), .I1(n2423), .CO(n25696));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n25694), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n25694), .I0(n2401), .I1(n2423), .CO(n25695));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n25693), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n25693), .I0(n2402), .I1(n2423), .CO(n25694));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n25692), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n25692), .I0(n2403), .I1(n2423), .CO(n25693));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n25691), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n25691), .I0(n2404), .I1(n2423), .CO(n25692));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n25690), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n25690), .I0(n2405), .I1(n2423), .CO(n25691));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n25689), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n16688), 
            .D(n255[5]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i17824_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n21925));
    defparam i17824_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut (.I0(n1405), .I1(n21925), .I2(n1403), .I3(n1406), 
            .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(n1408), .I2(n16), .I3(n1401), .O(n1433));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28830_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34504));
    defparam i28830_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28376_2_lut (.I0(n2), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i28376_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY mod_5_add_1674_6 (.CI(n25689), .I0(n2406), .I1(n2423), .CO(n25690));
    SB_LUT4 i28374_2_lut (.I0(n2), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i28374_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26549_3_lut (.I0(n906), .I1(n905), .I2(n30427), .I3(GND_net), 
            .O(n32222));
    defparam i26549_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1487 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10), 
            .O(n16_adj_4339));
    defparam i7_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1307), .I1(n16_adj_4339), .I2(n12), .I3(n1301), 
            .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(n16727), .I1(n32222), .I2(bit_ctr[26]), .I3(n14162), 
            .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h0111;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n14162), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26600_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n32274));
    defparam i26600_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut (.I0(n2), .I1(n6), .I2(n1005), .I3(n32274), .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i28380_2_lut (.I0(n2), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4));   // verilog/neopixel.v(22[26:36])
    defparam i28380_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n25688), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n25688), .I0(n2407), .I1(n2423), .CO(n25689));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n25687), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n25687), .I0(n2408), .I1(n2423), .CO(n25688));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n34489), 
            .I3(n25686), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n25781), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n25781), .I0(n2095), .I1(n2126), .CO(n25782));
    SB_LUT4 i28826_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34500));
    defparam i28826_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1674_3 (.CI(n25686), .I0(n2409), .I1(n34489), .CO(n25687));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n34489), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n34489), 
            .CO(n25686));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n25685), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n16688), 
            .D(n255[4]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n16688), 
            .D(n255[3]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n16688), 
            .D(n255[2]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n16688), 
            .D(n255[1]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n25684), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28823_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34497));
    defparam i28823_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut (.I0(bit_ctr[3]), .I1(n30), .I2(bit_ctr[13]), .I3(bit_ctr[4]), 
            .O(n43));
    defparam i15_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n25780), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n25684), .I0(n2490), .I1(n2522), .CO(n25685));
    SB_LUT4 i28829_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34503));
    defparam i28829_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1473_16 (.CI(n25780), .I0(n2096), .I1(n2126), .CO(n25781));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n25683), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n25683), .I0(n2491), .I1(n2522), .CO(n25684));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n25004), .O(one_wire_N_423[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n25779), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n25779), .I0(n2097), .I1(n2126), .CO(n25780));
    SB_CARRY sub_14_add_2_7 (.CI(n25004), .I0(timer[5]), .I1(n1[5]), .CO(n25005));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n25778), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n25682), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_20 (.CI(n25682), .I0(n2492), .I1(n2522), .CO(n25683));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n25681), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n25681), .I0(n2493), .I1(n2522), .CO(n25682));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n25680), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n25680), .I0(n2494), .I1(n2522), .CO(n25681));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n25679), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n25679), .I0(n2495), .I1(n2522), .CO(n25680));
    SB_CARRY mod_5_add_1473_14 (.CI(n25778), .I0(n2098), .I1(n2126), .CO(n25779));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n25777), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n25678), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n25678), .I0(n2496), .I1(n2522), .CO(n25679));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n25677), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n25677), .I0(n2497), .I1(n2522), .CO(n25678));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n25676), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n24812), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_13 (.CI(n25777), .I0(n2099), .I1(n2126), .CO(n25778));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n25776), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n25676), .I0(n2498), .I1(n2522), .CO(n25677));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n25675), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n25675), .I0(n2499), .I1(n2522), .CO(n25676));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n25674), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n25674), .I0(n2500), .I1(n2522), .CO(n25675));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n25673), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n25673), .I0(n2501), .I1(n2522), .CO(n25674));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n25672), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n25776), .I0(n2100), .I1(n2126), .CO(n25777));
    SB_CARRY mod_5_add_1741_10 (.CI(n25672), .I0(n2502), .I1(n2522), .CO(n25673));
    SB_LUT4 i15_4_lut_adj_1488 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42));
    defparam i15_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44_adj_4340));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1489 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43_adj_4341));
    defparam i16_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), .I3(GND_net), 
            .O(n40));
    defparam i13_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n25671), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n25671), .I0(n2503), .I1(n2522), .CO(n25672));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n25670), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n25670), .I0(n2504), .I1(n2522), .CO(n25671));
    SB_LUT4 i21_4_lut (.I0(n3107), .I1(n42), .I2(n3087), .I3(n3086), 
            .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n25669), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25_4_lut (.I0(n43_adj_4341), .I1(n45), .I2(n44_adj_4340), 
            .I3(n46), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_2_lut (.I0(n3095), .I1(n3084), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1741_7 (.CI(n25669), .I0(n2505), .I1(n2522), .CO(n25670));
    SB_LUT4 i6_4_lut_adj_1490 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14));
    defparam i6_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n39), .I1(n52), .I2(n48), .I3(n40), .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), .I3(GND_net), 
            .O(n9));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1491 (.I0(n9), .I1(n14), .I2(n1202), .I3(n1208), 
            .O(n1235));
    defparam i7_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_LUT4 i28821_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34495));
    defparam i28821_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n25668), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28828_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34502));
    defparam i28828_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26_4_lut_adj_1492 (.I0(n45_adj_4342), .I1(n47), .I2(n46_adj_4343), 
            .I3(n48_adj_4344), .O(n54));
    defparam i26_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 i17794_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n21895));
    defparam i17794_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n21895), .I3(n1108), 
            .O(n12_adj_4345));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1493 (.I0(n1107), .I1(n12_adj_4345), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n2206), .I1(n2204), .I2(n2194), .I3(n2196), 
            .O(n28_adj_4346));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17788_2_lut (.I0(bit_ctr[13]), .I1(n2209), .I2(GND_net), 
            .I3(GND_net), .O(n21889));
    defparam i17788_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14_3_lut (.I0(n2193), .I1(n28_adj_4346), .I2(n2198), .I3(GND_net), 
            .O(n32_adj_4347));
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut (.I0(n2208), .I1(n2192), .I2(n2205), .I3(n2201), 
            .O(n30_adj_4348));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2195), .I1(n2207), .I2(n21889), .I3(n2197), 
            .O(n31_adj_4349));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2202), .I1(n2200), .I2(n2199), .I3(n2203), 
            .O(n29));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1494 (.I0(n29), .I1(n31_adj_4349), .I2(n30_adj_4348), 
            .I3(n32_adj_4347), .O(n2225));
    defparam i17_4_lut_adj_1494.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_6 (.CI(n25668), .I0(n2506), .I1(n2522), .CO(n25669));
    SB_LUT4 i28820_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34494));
    defparam i28820_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n25667), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28816_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34490));
    defparam i28816_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1495 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4350));
    defparam i16_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1496 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4351));
    defparam i15_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1497 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37));
    defparam i13_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1498 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4352));
    defparam i18_4_lut_adj_1498.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n37), .I1(n39_adj_4351), .I2(n38), .I3(n40_adj_4350), 
            .O(n46_adj_4353));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4354));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut (.I0(n33_adj_4354), .I1(n46_adj_4353), .I2(n42_adj_4352), 
            .I3(n34), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28819_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34493));
    defparam i28819_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_5 (.CI(n25667), .I0(n2507), .I1(n2522), .CO(n25668));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n25666), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n25666), .I0(n2508), .I1(n2522), .CO(n25667));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n34491), 
            .I3(n25665), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_3 (.CI(n25665), .I0(n2509), .I1(n34491), .CO(n25666));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n34491), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n34491), 
            .CO(n25665));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n25664), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n25663), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n25663), .I0(n2589), .I1(n2621), .CO(n25664));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n25775), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n25662), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n25662), .I0(n2590), .I1(n2621), .CO(n25663));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n25661), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_21 (.CI(n25661), .I0(n2591), .I1(n2621), .CO(n25662));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n25660), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n25660), .I0(n2592), .I1(n2621), .CO(n25661));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n25659), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n25659), .I0(n2593), .I1(n2621), .CO(n25660));
    SB_CARRY mod_5_add_1473_11 (.CI(n25775), .I0(n2101), .I1(n2126), .CO(n25776));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n25658), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n25658), .I0(n2594), .I1(n2621), .CO(n25659));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n25657), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n16688), 
            .D(n255[31]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i21_4_lut_adj_1499 (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1808_17 (.CI(n25657), .I0(n2595), .I1(n2621), .CO(n25658));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n25656), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n25656), .I0(n2596), .I1(n2621), .CO(n25657));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n25655), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n25655), .I0(n2597), .I1(n2621), .CO(n25656));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n25654), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4357));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1500 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4358));
    defparam i15_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 i17802_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n21903));
    defparam i17802_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1501 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n21903), 
            .O(n36));
    defparam i13_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1502 (.I0(n2700), .I1(n38_adj_4358), .I2(n28_adj_4357), 
            .I3(n2705), .O(n42_adj_4359));
    defparam i19_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1503 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4360));
    defparam i17_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1504 (.I0(n2687), .I1(n36), .I2(n2703), .I3(n2695), 
            .O(n41));
    defparam i18_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1505 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4361));
    defparam i16_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1506 (.I0(n39_adj_4361), .I1(n41), .I2(n40_adj_4360), 
            .I3(n42_adj_4359), .O(n2720));
    defparam i22_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i28818_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34492));
    defparam i28818_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_14 (.CI(n25654), .I0(n2598), .I1(n2621), .CO(n25655));
    SB_LUT4 i14_4_lut_adj_1507 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4362));
    defparam i14_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1508 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25));
    defparam i3_3_lut_adj_1508.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1509 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4363));
    defparam i12_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1510 (.I0(n25), .I1(n36_adj_4362), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4364));
    defparam i18_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1511 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4365));
    defparam i16_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4363), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4366));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1512 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4367));
    defparam i15_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1513 (.I0(n37_adj_4367), .I1(n39_adj_4366), .I2(n38_adj_4365), 
            .I3(n40_adj_4364), .O(n2621));
    defparam i21_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n25774), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28817_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34491));
    defparam i28817_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1473_10 (.CI(n25774), .I0(n2102), .I1(n2126), .CO(n25775));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n25653), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n25653), .I0(n2599), .I1(n2621), .CO(n25654));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n25773), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n25652), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n25652), .I0(n2600), .I1(n2621), .CO(n25653));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n25651), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n25651), .I0(n2601), .I1(n2621), .CO(n25652));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n25650), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n25650), .I0(n2602), .I1(n2621), .CO(n25651));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n25649), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n25649), .I0(n2603), .I1(n2621), .CO(n25650));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n25648), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n25648), .I0(n2604), .I1(n2621), .CO(n25649));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n25647), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n25647), .I0(n2605), .I1(n2621), .CO(n25648));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n25646), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n25646), .I0(n2606), .I1(n2621), .CO(n25647));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n25645), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n25645), .I0(n2607), .I1(n2621), .CO(n25646));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n25644), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n25644), .I0(n2608), .I1(n2621), .CO(n25645));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n34492), 
            .I3(n25643), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n25643), .I0(n2609), .I1(n34492), .CO(n25644));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n34492), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n34492), 
            .CO(n25643));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n25642), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n25641), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n25641), .I0(n2688), .I1(n2720), .CO(n25642));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n25640), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n25640), .I0(n2689), .I1(n2720), .CO(n25641));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n25639), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n25773), .I0(n2103), .I1(n2126), .CO(n25774));
    SB_CARRY mod_5_add_1875_22 (.CI(n25639), .I0(n2690), .I1(n2720), .CO(n25640));
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_272[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1514 (.I0(one_wire_N_423[3]), .I1(one_wire_N_423[4]), 
            .I2(one_wire_N_423[2]), .I3(GND_net), .O(n26419));
    defparam i2_3_lut_adj_1514.LUT_INIT = 16'h8080;
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n25638), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n25638), .I0(n2691), .I1(n2720), .CO(n25639));
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n16688), 
            .D(n255[15]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n25637), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n25637), .I0(n2692), .I1(n2720), .CO(n25638));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n25636), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n25636), .I0(n2693), .I1(n2720), .CO(n25637));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n25772), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n25635), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n16688), 
            .D(n255[14]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n25003), .O(one_wire_N_423[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_8 (.CI(n25772), .I0(n2104), .I1(n2126), .CO(n25773));
    SB_CARRY mod_5_add_1875_18 (.CI(n25635), .I0(n2694), .I1(n2720), .CO(n25636));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n25634), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n25634), .I0(n2695), .I1(n2720), .CO(n25635));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n25633), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n25633), .I0(n2696), .I1(n2720), .CO(n25634));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n25632), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n25632), .I0(n2697), .I1(n2720), .CO(n25633));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n25631), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n25631), .I0(n2698), .I1(n2720), .CO(n25632));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n25630), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n25630), .I0(n2699), .I1(n2720), .CO(n25631));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n25629), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n25629), .I0(n2700), .I1(n2720), .CO(n25630));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n25771), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_6 (.CI(n25003), .I0(timer[4]), .I1(n1[4]), .CO(n25004));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n25628), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n25628), .I0(n2701), .I1(n2720), .CO(n25629));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n25627), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n25627), .I0(n2702), .I1(n2720), .CO(n25628));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n25002), .O(one_wire_N_423[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n25626), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n25626), .I0(n2703), .I1(n2720), .CO(n25627));
    SB_CARRY mod_5_add_1473_7 (.CI(n25771), .I0(n2105), .I1(n2126), .CO(n25772));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n25625), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n24820), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_8 (.CI(n25625), .I0(n2704), .I1(n2720), .CO(n25626));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n25770), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n25624), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n25624), .I0(n2705), .I1(n2720), .CO(n25625));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n25623), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n25770), .I0(n2106), .I1(n2126), .CO(n25771));
    SB_CARRY mod_5_add_1875_6 (.CI(n25623), .I0(n2706), .I1(n2720), .CO(n25624));
    SB_LUT4 i1_2_lut_adj_1515 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n15574));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut_adj_1515.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_3_lut_adj_1516 (.I0(n26673), .I1(one_wire_N_423[4]), .I2(one_wire_N_423[3]), 
            .I3(GND_net), .O(n30348));
    defparam i1_3_lut_adj_1516.LUT_INIT = 16'hecec;
    SB_LUT4 i6_4_lut_adj_1517 (.I0(one_wire_N_423[5]), .I1(one_wire_N_423[11]), 
            .I2(one_wire_N_423[7]), .I3(n15581), .O(n14_adj_4368));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n16688), 
            .D(n255[8]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i7_4_lut_adj_1518 (.I0(n9_adj_4369), .I1(n14_adj_4368), .I2(one_wire_N_423[10]), 
            .I3(one_wire_N_423[8]), .O(n15471));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n25769), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n25622), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n25769), .I0(n2107), .I1(n2126), .CO(n25770));
    SB_CARRY mod_5_add_1875_5 (.CI(n25622), .I0(n2707), .I1(n2720), .CO(n25623));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n25621), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n25621), .I0(n2708), .I1(n2720), .CO(n25622));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n34493), 
            .I3(n25620), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n25620), .I0(n2709), .I1(n34493), .CO(n25621));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n25768), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n25768), .I0(n2108), .I1(n2126), .CO(n25769));
    SB_LUT4 i181_2_lut (.I0(LED_c), .I1(\state_3__N_272[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/neopixel.v(40[18] 45[12])
    defparam i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n34493), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n34493), 
            .CO(n25620));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n25619), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n25618), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n25618), .I0(n2787), .I1(n2819), .CO(n25619));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n25617), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n25617), .I0(n2788), .I1(n2819), .CO(n25618));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n25616), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n25616), .I0(n2789), .I1(n2819), .CO(n25617));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n25615), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n25615), .I0(n2790), .I1(n2819), .CO(n25616));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n25614), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n16688), 
            .D(n255[7]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1942_21 (.CI(n25614), .I0(n2791), .I1(n2819), .CO(n25615));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n34490), 
            .I3(n25767), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n25613), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n25613), .I0(n2792), .I1(n2819), .CO(n25614));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n25612), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n25612), .I0(n2793), .I1(n2819), .CO(n25613));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n25611), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n25611), .I0(n2794), .I1(n2819), .CO(n25612));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n25610), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n25610), .I0(n2795), .I1(n2819), .CO(n25611));
    SB_CARRY mod_5_add_1473_3 (.CI(n25767), .I0(n2109), .I1(n34490), .CO(n25768));
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n25609), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n25609), .I0(n2796), .I1(n2819), .CO(n25610));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n25608), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n25608), .I0(n2797), .I1(n2819), .CO(n25609));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n25607), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n25607), .I0(n2798), .I1(n2819), .CO(n25608));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n34490), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n25606), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n25606), .I0(n2799), .I1(n2819), .CO(n25607));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n25605), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n25605), .I0(n2800), .I1(n2819), .CO(n25606));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n25604), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n25604), .I0(n2801), .I1(n2819), .CO(n25605));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n25603), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n25603), .I0(n2802), .I1(n2819), .CO(n25604));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n25602), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n25602), .I0(n2803), .I1(n2819), .CO(n25603));
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n34490), 
            .CO(n25767));
    SB_CARRY sub_14_add_2_5 (.CI(n25002), .I0(timer[3]), .I1(n1[3]), .CO(n25003));
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28024_4_lut (.I0(n26419), .I1(n30348), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n33493));
    defparam i28024_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i27822_2_lut (.I0(n30348), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n33192));
    defparam i27822_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53_4_lut (.I0(n33192), .I1(n21971), .I2(\state[1] ), .I3(n15471), 
            .O(n30455));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n30455), .I1(n33494), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n30475));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i80_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_486 ));
    defparam i80_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n25601), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n25601), .I0(n2804), .I1(n2819), .CO(n25602));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n25600), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n25600), .I0(n2805), .I1(n2819), .CO(n25601));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n25599), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n25599), .I0(n2806), .I1(n2819), .CO(n25600));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n25598), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n25598), .I0(n2807), .I1(n2819), .CO(n25599));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n25597), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n25597), .I0(n2808), .I1(n2819), .CO(n25598));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n34494), 
            .I3(n25596), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n25596), .I0(n2809), .I1(n34494), .CO(n25597));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n34494), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n34494), 
            .CO(n25596));
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n25766), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n25595), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n25594), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n25594), .I0(n1104), .I1(n1136), .CO(n25595));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n25593), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n25593), .I0(n1105), .I1(n1136), .CO(n25594));
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n25765), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n25592), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n25592), .I0(n1106), .I1(n1136), .CO(n25593));
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n25591), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1519 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4373));
    defparam i13_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1520 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22));
    defparam i1_3_lut_adj_1520.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1521 (.I0(n2490), .I1(n34_adj_4373), .I2(n24), 
            .I3(n2494), .O(n38_adj_4374));
    defparam i17_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1522 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4375));
    defparam i15_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1523 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22), 
            .O(n37_adj_4376));
    defparam i16_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1524 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35));
    defparam i14_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37_adj_4376), .I2(n36_adj_4375), 
            .I3(n38_adj_4374), .O(n2522));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_803_5 (.CI(n25591), .I0(n1107), .I1(n1136), .CO(n25592));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n25590), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(n15471), .I1(n30348), .I2(GND_net), .I3(GND_net), 
            .O(n22039));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n25001), .O(one_wire_N_423[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_4 (.CI(n25590), .I0(n1108), .I1(n1136), .CO(n25591));
    SB_CARRY sub_14_add_2_4 (.CI(n25001), .I0(timer[2]), .I1(n1[2]), .CO(n25002));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n34495), 
            .I3(n25589), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n25589), .I0(n1109), .I1(n34495), .CO(n25590));
    SB_CARRY mod_5_add_1540_19 (.CI(n25765), .I0(n2193), .I1(n2225), .CO(n25766));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n34495), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n34495), 
            .CO(n25589));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n25144), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n25143), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n25764), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n25143), .I0(n1203), .I1(n1235), .CO(n25144));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n25142), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n25142), .I0(n1204), .I1(n1235), .CO(n25143));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n25141), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4377), .I1(timer[1]), .I2(n1[1]), 
            .I3(n25000), .O(n26673)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_3 (.CI(n25000), .I0(timer[1]), .I1(n1[1]), .CO(n25001));
    SB_LUT4 i17816_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n21917));
    defparam i17816_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1525 (.I0(n35_adj_4378), .I1(n11), .I2(n29_adj_4379), 
            .I3(n51), .O(n48_adj_4380));
    defparam i20_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1526 (.I0(n37_adj_4381), .I1(n23), .I2(n53), 
            .I3(n39_adj_4382), .O(n46_adj_4383));
    defparam i18_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_870_7 (.CI(n25141), .I0(n1205), .I1(n1235), .CO(n25142));
    SB_LUT4 i19_4_lut_adj_1527 (.I0(n27), .I1(n57), .I2(n63), .I3(n43_adj_4384), 
            .O(n47_adj_4385));
    defparam i19_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1528 (.I0(n25_adj_4386), .I1(n33_adj_4387), .I2(n47_adj_4388), 
            .I3(n61), .O(n45_adj_4389));
    defparam i17_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1529 (.I0(n59), .I1(n17_adj_4390), .I2(n15_adj_4391), 
            .I3(n55), .O(n44_adj_4392));
    defparam i16_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1530 (.I0(n31_adj_4393), .I1(n41_adj_4394), .I2(n49_adj_4395), 
            .I3(n21917), .O(n43_adj_4396));
    defparam i15_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1531 (.I0(n45_adj_4389), .I1(n47_adj_4385), .I2(n46_adj_4383), 
            .I3(n48_adj_4380), .O(n54_adj_4397));
    defparam i26_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1532 (.I0(n45_adj_4398), .I1(n13_adj_4399), .I2(n19_adj_4400), 
            .I3(n21_adj_4401), .O(n49_adj_4402));
    defparam i21_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut_adj_1533 (.I0(n49_adj_4402), .I1(n54_adj_4397), .I2(n43_adj_4396), 
            .I3(n44_adj_4392), .O(n26709));
    defparam i27_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_rep_240_2_lut (.I0(bit_ctr[3]), .I1(n26709), .I2(GND_net), 
            .I3(GND_net), .O(n35413));
    defparam i1_rep_240_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n25140), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i27912_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n26709), .I3(GND_net), 
            .O(color_bit_N_466[4]));
    defparam i27912_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i27992_4_lut (.I0(n34714), .I1(n35413), .I2(n34612), .I3(bit_ctr[2]), 
            .O(n33147));
    defparam i27992_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY mod_5_add_1540_18 (.CI(n25764), .I0(n2194), .I1(n2225), .CO(n25765));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n25763), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n25140), .I0(n1206), .I1(n1235), .CO(n25141));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n25139), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n25139), .I0(n1207), .I1(n1235), .CO(n25140));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_423[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_adj_4377)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i17070_4_lut (.I0(n34528), .I1(\state_3__N_272[1] ), .I2(n33147), 
            .I3(color_bit_N_466[4]), .O(state_3__N_272[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i17070_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n25000));
    SB_CARRY mod_5_add_1540_17 (.CI(n25763), .I0(n2195), .I1(n2225), .CO(n25764));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n25762), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n25138), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n25138), .I0(n1208), .I1(n1235), .CO(n25139));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n34497), 
            .I3(n25137), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i2846_4_lut (.I0(n22039), .I1(n831), .I2(\state[1] ), .I3(n15574), 
            .O(n4081));
    defparam i2846_4_lut.LUT_INIT = 16'h3f35;
    SB_CARRY mod_5_add_870_3 (.CI(n25137), .I0(n1209), .I1(n34497), .CO(n25138));
    SB_CARRY mod_5_add_1540_16 (.CI(n25762), .I0(n2196), .I1(n2225), .CO(n25763));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n25761), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n25761), .I0(n2197), .I1(n2225), .CO(n25762));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n34497), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_1534 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4404));
    defparam i1_2_lut_adj_1534.LUT_INIT = 16'heeee;
    SB_LUT4 i17786_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n21887));
    defparam i17786_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1535 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_4404), 
            .O(n30_adj_4405));
    defparam i13_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1536 (.I0(n2098), .I1(n21887), .I2(n2094), .I3(n2099), 
            .O(n28_adj_4406));
    defparam i11_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1537 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4407));
    defparam i12_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1538 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4408));
    defparam i10_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n25760), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n34497), 
            .CO(n25137));
    SB_CARRY mod_5_add_1540_14 (.CI(n25760), .I0(n2198), .I1(n2225), .CO(n25761));
    SB_LUT4 i16_4_lut_adj_1539 (.I0(n27_adj_4408), .I1(n29_adj_4407), .I2(n28_adj_4406), 
            .I3(n30_adj_4405), .O(n2126));
    defparam i16_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n25136), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n25759), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n25759), .I0(n2199), .I1(n2225), .CO(n25760));
    SB_LUT4 i28815_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34489));
    defparam i28815_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n25758), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n25758), .I0(n2200), .I1(n2225), .CO(n25759));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n25757), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n25757), .I0(n2201), .I1(n2225), .CO(n25758));
    SB_LUT4 i2_2_lut_adj_1540 (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30));
    defparam i2_2_lut_adj_1540.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_1541 (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48_adj_4344));
    defparam i20_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n25135), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18_4_lut_adj_1542 (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46_adj_4343));
    defparam i18_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1543 (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1544 (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45_adj_4342));
    defparam i17_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i28367_4_lut (.I0(\state[1] ), .I1(n33174), .I2(\state[0] ), 
            .I3(n4081), .O(n16688));
    defparam i28367_4_lut.LUT_INIT = 16'h01f1;
    SB_CARRY mod_5_add_937_10 (.CI(n25135), .I0(n1302), .I1(n1334), .CO(n25136));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n25756), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n25134), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n25134), .I0(n1303), .I1(n1334), .CO(n25135));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n25133), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n25133), .I0(n1304), .I1(n1334), .CO(n25134));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n25132), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1125_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n25530), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1125_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n25529), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_32 (.CI(n25529), .I0(GND_net), .I1(timer[30]), 
            .CO(n25530));
    SB_CARRY mod_5_add_1540_10 (.CI(n25756), .I0(n2202), .I1(n2225), .CO(n25757));
    SB_LUT4 timer_1125_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n25528), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_7 (.CI(n25132), .I0(n1305), .I1(n1334), .CO(n25133));
    SB_CARRY timer_1125_add_4_31 (.CI(n25528), .I0(GND_net), .I1(timer[29]), 
            .CO(n25529));
    SB_LUT4 timer_1125_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n25527), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n25131), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n25755), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1125_add_4_30 (.CI(n25527), .I0(GND_net), .I1(timer[28]), 
            .CO(n25528));
    SB_CARRY mod_5_add_1540_9 (.CI(n25755), .I0(n2203), .I1(n2225), .CO(n25756));
    SB_LUT4 timer_1125_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n25526), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_29 (.CI(n25526), .I0(GND_net), .I1(timer[27]), 
            .CO(n25527));
    SB_LUT4 timer_1125_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n25525), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_28 (.CI(n25525), .I0(GND_net), .I1(timer[26]), 
            .CO(n25526));
    SB_LUT4 timer_1125_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n25524), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_27 (.CI(n25524), .I0(GND_net), .I1(timer[25]), 
            .CO(n25525));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n25754), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1125_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n25523), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_26 (.CI(n25523), .I0(GND_net), .I1(timer[24]), 
            .CO(n25524));
    SB_LUT4 timer_1125_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n25522), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_25 (.CI(n25522), .I0(GND_net), .I1(timer[23]), 
            .CO(n25523));
    SB_LUT4 timer_1125_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n25521), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_24 (.CI(n25521), .I0(GND_net), .I1(timer[22]), 
            .CO(n25522));
    SB_CARRY mod_5_add_937_6 (.CI(n25131), .I0(n1306), .I1(n1334), .CO(n25132));
    SB_CARRY mod_5_add_1540_8 (.CI(n25754), .I0(n2204), .I1(n2225), .CO(n25755));
    SB_LUT4 timer_1125_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n25520), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_23 (.CI(n25520), .I0(GND_net), .I1(timer[21]), 
            .CO(n25521));
    SB_LUT4 timer_1125_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n25519), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_22 (.CI(n25519), .I0(GND_net), .I1(timer[20]), 
            .CO(n25520));
    SB_LUT4 timer_1125_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n25518), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n25130), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n25130), .I0(n1307), .I1(n1334), .CO(n25131));
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n16688), 
            .D(n255[0]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i14_4_lut_adj_1545 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4409));
    defparam i14_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1546 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4410));
    defparam i18_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1547 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_4411));
    defparam i16_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1548 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4412));
    defparam i17_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1549 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4413));
    defparam i15_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut_adj_1550 (.I0(n3001), .I1(n2993), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4414));
    defparam i12_2_lut_adj_1550.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4409), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4415));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n41_adj_4413), .I1(n43_adj_4412), .I2(n42_adj_4411), 
            .I3(n44_adj_4410), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4416));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut_adj_1551 (.I0(n37_adj_4416), .I1(n50), .I2(n46_adj_4415), 
            .I3(n38_adj_4414), .O(n3017));
    defparam i25_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i28825_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34499));
    defparam i28825_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1125_add_4_21 (.CI(n25518), .I0(GND_net), .I1(timer[19]), 
            .CO(n25519));
    SB_LUT4 timer_1125_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n25517), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_20 (.CI(n25517), .I0(GND_net), .I1(timer[18]), 
            .CO(n25518));
    SB_LUT4 timer_1125_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n25516), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_19 (.CI(n25516), .I0(GND_net), .I1(timer[17]), 
            .CO(n25517));
    SB_LUT4 timer_1125_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n25515), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_18 (.CI(n25515), .I0(GND_net), .I1(timer[16]), 
            .CO(n25516));
    SB_CARRY add_21_5 (.CI(n24812), .I0(bit_ctr[3]), .I1(GND_net), .CO(n24813));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n25129), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1125_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n25514), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_17 (.CI(n25514), .I0(GND_net), .I1(timer[15]), 
            .CO(n25515));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n25753), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1125_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n25513), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_16 (.CI(n25513), .I0(GND_net), .I1(timer[14]), 
            .CO(n25514));
    SB_LUT4 timer_1125_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n25512), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_15 (.CI(n25512), .I0(GND_net), .I1(timer[13]), 
            .CO(n25513));
    SB_LUT4 timer_1125_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n25511), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_14 (.CI(n25511), .I0(GND_net), .I1(timer[12]), 
            .CO(n25512));
    SB_LUT4 timer_1125_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n25510), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_13 (.CI(n25510), .I0(GND_net), .I1(timer[11]), 
            .CO(n25511));
    SB_LUT4 timer_1125_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n25509), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_12 (.CI(n25509), .I0(GND_net), .I1(timer[10]), 
            .CO(n25510));
    SB_LUT4 timer_1125_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n25508), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_11 (.CI(n25508), .I0(GND_net), .I1(timer[9]), 
            .CO(n25509));
    SB_CARRY mod_5_add_1540_7 (.CI(n25753), .I0(n2205), .I1(n2225), .CO(n25754));
    SB_CARRY mod_5_add_937_4 (.CI(n25129), .I0(n1308), .I1(n1334), .CO(n25130));
    SB_LUT4 timer_1125_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n25507), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n34498), 
            .I3(n25128), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1125_add_4_10 (.CI(n25507), .I0(GND_net), .I1(timer[8]), 
            .CO(n25508));
    SB_LUT4 timer_1125_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n25506), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_9 (.CI(n25506), .I0(GND_net), .I1(timer[7]), 
            .CO(n25507));
    SB_LUT4 timer_1125_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n25505), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_8 (.CI(n25505), .I0(GND_net), .I1(timer[6]), 
            .CO(n25506));
    SB_LUT4 timer_1125_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n25504), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_3 (.CI(n25128), .I0(n1309), .I1(n34498), .CO(n25129));
    SB_CARRY timer_1125_add_4_7 (.CI(n25504), .I0(GND_net), .I1(timer[5]), 
            .CO(n25505));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n25752), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n16688), 
            .D(n255[30]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_1125_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n25503), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_6 (.CI(n25503), .I0(GND_net), .I1(timer[4]), 
            .CO(n25504));
    SB_LUT4 timer_1125_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n25502), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_5 (.CI(n25502), .I0(GND_net), .I1(timer[3]), 
            .CO(n25503));
    SB_LUT4 timer_1125_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n25501), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_4 (.CI(n25501), .I0(GND_net), .I1(timer[2]), 
            .CO(n25502));
    SB_LUT4 timer_1125_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n25500), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1125_add_4_3 (.CI(n25500), .I0(GND_net), .I1(timer[1]), 
            .CO(n25501));
    SB_LUT4 timer_1125_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1125_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n34498), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1125_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n25500));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n25499), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n25498), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n34498), 
            .CO(n25128));
    SB_CARRY mod_5_add_1540_6 (.CI(n25752), .I0(n2206), .I1(n2225), .CO(n25753));
    SB_CARRY mod_5_add_2009_26 (.CI(n25498), .I0(n2886), .I1(n2918), .CO(n25499));
    SB_CARRY add_21_13 (.CI(n24820), .I0(bit_ctr[11]), .I1(GND_net), .CO(n24821));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n25497), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n25497), .I0(n2887), .I1(n2918), .CO(n25498));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n25496), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n25496), .I0(n2888), .I1(n2918), .CO(n25497));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n25495), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n25495), .I0(n2889), .I1(n2918), .CO(n25496));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n25494), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n25494), .I0(n2890), .I1(n2918), .CO(n25495));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n25493), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n25493), .I0(n2891), .I1(n2918), .CO(n25494));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n25492), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n25492), .I0(n2892), .I1(n2918), .CO(n25493));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n25491), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n24840), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n25127), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_19 (.CI(n25491), .I0(n2893), .I1(n2918), .CO(n25492));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n25490), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n24839), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_18 (.CI(n25490), .I0(n2894), .I1(n2918), .CO(n25491));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n25489), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n25126), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_17 (.CI(n25489), .I0(n2895), .I1(n2918), .CO(n25490));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n25488), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_32 (.CI(n24839), .I0(bit_ctr[30]), .I1(GND_net), .CO(n24840));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n24838), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n25751), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n25488), .I0(n2896), .I1(n2918), .CO(n25489));
    SB_CARRY mod_5_add_669_6 (.CI(n25126), .I0(n906), .I1(VCC_net), .CO(n25127));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n30427), .I2(VCC_net), 
            .I3(n25125), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n25487), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_5 (.CI(n25125), .I0(n30427), .I1(VCC_net), 
            .CO(n25126));
    SB_CARRY mod_5_add_1540_5 (.CI(n25751), .I0(n2207), .I1(n2225), .CO(n25752));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n16727), .I2(VCC_net), 
            .I3(n25124), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n25124), .I0(n16727), .I1(VCC_net), 
            .CO(n25125));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n25750), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n25487), .I0(n2897), .I1(n2918), .CO(n25488));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n25486), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n25486), .I0(n2898), .I1(n2918), .CO(n25487));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n14162), .I2(GND_net), 
            .I3(n25123), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n25485), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_3 (.CI(n25123), .I0(n14162), .I1(GND_net), 
            .CO(n25124));
    SB_CARRY mod_5_add_2009_13 (.CI(n25485), .I0(n2899), .I1(n2918), .CO(n25486));
    SB_CARRY add_21_31 (.CI(n24838), .I0(bit_ctr[29]), .I1(GND_net), .CO(n24839));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n25484), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n25484), .I0(n2900), .I1(n2918), .CO(n25485));
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n25123));
    SB_CARRY mod_5_add_1540_4 (.CI(n25750), .I0(n2208), .I1(n2225), .CO(n25751));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n34496), 
            .I3(n25749), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n25749), .I0(n2209), .I1(n34496), .CO(n25750));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n34496), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_2_lut_adj_1552 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4417));
    defparam i3_2_lut_adj_1552.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n34496), 
            .CO(n25749));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n25748), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_1553 (.I0(bit_ctr[12]), .I1(n22_adj_4417), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4418));
    defparam i11_4_lut_adj_1553.LUT_INIT = 16'hfefc;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n25747), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n25747), .I0(n2292), .I1(n2324), .CO(n25748));
    SB_LUT4 i15_4_lut_adj_1554 (.I0(n2294), .I1(n30_adj_4418), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4419));
    defparam i15_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n25746), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n25746), .I0(n2293), .I1(n2324), .CO(n25747));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n25745), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n25483), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n25483), .I0(n2901), .I1(n2918), .CO(n25484));
    SB_CARRY mod_5_add_1607_18 (.CI(n25745), .I0(n2294), .I1(n2324), .CO(n25746));
    SB_LUT4 i13_4_lut_adj_1555 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4420));
    defparam i13_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1556 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4421));
    defparam i14_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n25482), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n25482), .I0(n2902), .I1(n2918), .CO(n25483));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n25481), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n25481), .I0(n2903), .I1(n2918), .CO(n25482));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n25480), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n25480), .I0(n2904), .I1(n2918), .CO(n25481));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n25479), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n25479), .I0(n2905), .I1(n2918), .CO(n25480));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n25478), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n25478), .I0(n2906), .I1(n2918), .CO(n25479));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n25744), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n25477), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n24837), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_17 (.CI(n25744), .I0(n2295), .I1(n2324), .CO(n25745));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n25743), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_30 (.CI(n24837), .I0(bit_ctr[28]), .I1(GND_net), .CO(n24838));
    SB_CARRY mod_5_add_1607_16 (.CI(n25743), .I0(n2296), .I1(n2324), .CO(n25744));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n25742), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n25477), .I0(n2907), .I1(n2918), .CO(n25478));
    SB_CARRY mod_5_add_1607_15 (.CI(n25742), .I0(n2297), .I1(n2324), .CO(n25743));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n25741), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n25741), .I0(n2298), .I1(n2324), .CO(n25742));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n25476), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_4_lut_adj_1557 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4422));
    defparam i12_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1558 (.I0(n31_adj_4422), .I1(n33_adj_4421), .I2(n32_adj_4420), 
            .I3(n34_adj_4419), .O(n2324));
    defparam i18_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i28822_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34496));
    defparam i28822_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n24836), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n24836), .I0(bit_ctr[27]), .I1(GND_net), .CO(n24837));
    SB_CARRY mod_5_add_2009_4 (.CI(n25476), .I0(n2908), .I1(n2918), .CO(n25477));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n34499), 
            .I3(n25475), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n24835), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n25740), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_28 (.CI(n24835), .I0(bit_ctr[26]), .I1(GND_net), .CO(n24836));
    SB_CARRY mod_5_add_2009_3 (.CI(n25475), .I0(n2909), .I1(n34499), .CO(n25476));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n34499), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_13 (.CI(n25740), .I0(n2299), .I1(n2324), .CO(n25741));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n34499), 
            .CO(n25475));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n25474), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n25473), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n25739), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1559 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n14162));
    defparam i1_2_lut_adj_1559.LUT_INIT = 16'h9999;
    SB_CARRY mod_5_add_2076_27 (.CI(n25473), .I0(n2985), .I1(n3017), .CO(n25474));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n25472), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_CARRY mod_5_add_2076_26 (.CI(n25472), .I0(n2986), .I1(n3017), .CO(n25473));
    SB_CARRY mod_5_add_1607_12 (.CI(n25739), .I0(n2300), .I1(n2324), .CO(n25740));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n25738), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n25471), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17702_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i17702_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n21867), .I2(n6706), .I3(n608), 
            .O(n30429));
    defparam i2_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_adj_1560 (.I0(bit_ctr[28]), .I1(n30429), .I2(GND_net), 
            .I3(GND_net), .O(n14164));
    defparam i1_2_lut_adj_1560.LUT_INIT = 16'h9999;
    SB_LUT4 i26525_3_lut (.I0(n30429), .I1(n708), .I2(n6706), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam i26525_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_DFF timer_1125__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4423));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n16688), 
            .D(n255[29]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i16_4_lut_adj_1561 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_4424));
    defparam i16_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut_adj_1562 (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_4425));
    defparam i13_3_lut_adj_1562.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1563 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43_adj_4426));
    defparam i18_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1564 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_4427));
    defparam i15_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1565 (.I0(n41_adj_4424), .I1(n33_adj_4423), .I2(n2889), 
            .I3(n2901), .O(n46_adj_4428));
    defparam i21_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_25 (.CI(n25471), .I0(n2987), .I1(n3017), .CO(n25472));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n25470), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n25470), .I0(n2988), .I1(n3017), .CO(n25471));
    SB_LUT4 i14_4_lut_adj_1566 (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39_adj_4429));
    defparam i14_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1567 (.I0(n43_adj_4426), .I1(n2904), .I2(n38_adj_4425), 
            .I3(n2893), .O(n47_adj_4430));
    defparam i22_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n25469), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n25469), .I0(n2989), .I1(n3017), .CO(n25470));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n25468), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i24_4_lut_adj_1568 (.I0(n47_adj_4430), .I1(n39_adj_4429), .I2(n46_adj_4428), 
            .I3(n40_adj_4427), .O(n2918));
    defparam i24_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_22 (.CI(n25468), .I0(n2990), .I1(n3017), .CO(n25469));
    SB_CARRY mod_5_add_1607_11 (.CI(n25738), .I0(n2301), .I1(n2324), .CO(n25739));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n25467), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n25467), .I0(n2991), .I1(n3017), .CO(n25468));
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n16688), 
            .D(n255[28]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n25466), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n25466), .I0(n2992), .I1(n3017), .CO(n25467));
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n16688), 
            .D(n255[13]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n16688), 
            .D(n255[27]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n25465), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n25737), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n25465), .I0(n2993), .I1(n3017), .CO(n25466));
    SB_CARRY mod_5_add_1607_10 (.CI(n25737), .I0(n2302), .I1(n2324), .CO(n25738));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n25464), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28824_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34498));
    defparam i28824_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_18 (.CI(n25464), .I0(n2994), .I1(n3017), .CO(n25465));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n25463), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n25463), .I0(n2995), .I1(n3017), .CO(n25464));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n25462), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n25462), .I0(n2996), .I1(n3017), .CO(n25463));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n25461), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n25461), .I0(n2997), .I1(n3017), .CO(n25462));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n25460), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n25460), .I0(n2998), .I1(n3017), .CO(n25461));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n25459), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n25459), .I0(n2999), .I1(n3017), .CO(n25460));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n25458), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n24834), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_12 (.CI(n25458), .I0(n3000), .I1(n3017), .CO(n25459));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n25457), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n25457), .I0(n3001), .I1(n3017), .CO(n25458));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n25456), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n25456), .I0(n3002), .I1(n3017), .CO(n25457));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n25455), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n25455), .I0(n3003), .I1(n3017), .CO(n25456));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n25454), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n25454), .I0(n3004), .I1(n3017), .CO(n25455));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n25453), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n25453), .I0(n3005), .I1(n3017), .CO(n25454));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n25452), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n25452), .I0(n3006), .I1(n3017), .CO(n25453));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n25451), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n25736), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n25451), .I0(n3007), .I1(n3017), .CO(n25452));
    SB_CARRY mod_5_add_1607_9 (.CI(n25736), .I0(n2303), .I1(n2324), .CO(n25737));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n25450), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n25450), .I0(n3008), .I1(n3017), .CO(n25451));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n34502), 
            .I3(n25449), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n25449), .I0(n3009), .I1(n34502), .CO(n25450));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n34502), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n34502), 
            .CO(n25449));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n25735), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n25735), .I0(n2304), .I1(n2324), .CO(n25736));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n25448), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n25734), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n25734), .I0(n2305), .I1(n2324), .CO(n25735));
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n25447), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n25733), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n25733), .I0(n2306), .I1(n2324), .CO(n25734));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n25732), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n25447), .I0(n3084), .I1(n3116), .CO(n25448));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n25446), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n25446), .I0(n3085), .I1(n3116), .CO(n25447));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n25445), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n25445), .I0(n3086), .I1(n3116), .CO(n25446));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n25444), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n25444), .I0(n3087), .I1(n3116), .CO(n25445));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n25443), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n25443), .I0(n3088), .I1(n3116), .CO(n25444));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n25442), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n25442), .I0(n3089), .I1(n3116), .CO(n25443));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n25441), .O(n49_adj_4395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n25441), .I0(n3090), .I1(n3116), .CO(n25442));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n25440), .O(n47_adj_4388)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n25440), .I0(n3091), .I1(n3116), .CO(n25441));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n25439), .O(n45_adj_4398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n25439), .I0(n3092), .I1(n3116), .CO(n25440));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n25438), .O(n43_adj_4384)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n25438), .I0(n3093), .I1(n3116), .CO(n25439));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n25437), .O(n41_adj_4394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n25437), .I0(n3094), .I1(n3116), .CO(n25438));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n25436), .O(n39_adj_4382)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n25436), .I0(n3095), .I1(n3116), .CO(n25437));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n25435), .O(n37_adj_4381)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n25435), .I0(n3096), .I1(n3116), .CO(n25436));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n25434), .O(n35_adj_4378)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n25434), .I0(n3097), .I1(n3116), .CO(n25435));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n25433), .O(n33_adj_4387)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n25433), .I0(n3098), .I1(n3116), .CO(n25434));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n25432), .O(n31_adj_4393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n25732), .I0(n2307), .I1(n2324), .CO(n25733));
    SB_CARRY mod_5_add_2143_13 (.CI(n25432), .I0(n3099), .I1(n3116), .CO(n25433));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n25431), .O(n29_adj_4379)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n25431), .I0(n3100), .I1(n3116), .CO(n25432));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n25430), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n25430), .I0(n3101), .I1(n3116), .CO(n25431));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n25429), .O(n25_adj_4386)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n25731), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n25429), .I0(n3102), .I1(n3116), .CO(n25430));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n25428), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n25428), .I0(n3103), .I1(n3116), .CO(n25429));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n25427), .O(n21_adj_4401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n25427), .I0(n3104), .I1(n3116), .CO(n25428));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n25426), .O(n19_adj_4400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n25426), .I0(n3105), .I1(n3116), .CO(n25427));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n25425), .O(n17_adj_4390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n25425), .I0(n3106), .I1(n3116), .CO(n25426));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n25424), .O(n15_adj_4391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n25424), .I0(n3107), .I1(n3116), .CO(n25425));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n25423), .O(n13_adj_4399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n25423), .I0(n3108), .I1(n3116), .CO(n25424));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n34503), 
            .I3(n25422), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n25422), .I0(n3109), .I1(n34503), .CO(n25423));
    SB_CARRY mod_5_add_1607_4 (.CI(n25731), .I0(n2308), .I1(n2324), .CO(n25732));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n34503), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n34503), 
            .CO(n25422));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n24819), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n34500), 
            .I3(n25730), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i4550_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n30429), .I2(bit_ctr[27]), 
            .I3(n30302), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i4550_2_lut_3_lut_4_lut.LUT_INIT = 16'hff60;
    SB_CARRY mod_5_add_1607_3 (.CI(n25730), .I0(n2309), .I1(n34500), .CO(n25731));
    SB_CARRY add_21_27 (.CI(n24834), .I0(bit_ctr[25]), .I1(GND_net), .CO(n24835));
    SB_LUT4 i27529_2_lut_3_lut (.I0(n21971), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[0] ), .I3(GND_net), .O(n33100));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27529_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut (.I0(n22115), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n30261));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), .I3(GND_net), 
            .O(n27_adj_4431));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1569 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4432));
    defparam i13_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n34711));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n34711_bdd_4_lut (.I0(n34711), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n34714));
    defparam n34711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1570 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4433));
    defparam i12_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1571 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4434));
    defparam i11_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i195_2_lut (.I0(n21971), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n845));   // verilog/neopixel.v(103[9] 111[12])
    defparam i195_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1572 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4435));
    defparam i15_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(\state[0] ), .I1(n30261), .I2(n845), .I3(\state[1] ), 
            .O(n16698));
    defparam i1_4_lut.LUT_INIT = 16'hafcc;
    SB_LUT4 i17_4_lut_adj_1573 (.I0(n33_adj_4432), .I1(n27_adj_4431), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4436));
    defparam i17_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1574 (.I0(n22115), .I1(n33100), .I2(\state[1] ), 
            .I3(n15574), .O(n30267));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1574.LUT_INIT = 16'h303a;
    SB_LUT4 i19_4_lut_adj_1575 (.I0(n37_adj_4436), .I1(n35_adj_4435), .I2(n31_adj_4434), 
            .I3(n32_adj_4433), .O(n2423));
    defparam i19_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1576 (.I0(n21_adj_4437), .I1(n23_adj_4438), .I2(n22_adj_4439), 
            .I3(n24_adj_4440), .O(n36_adj_4441));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1577 (.I0(n25_adj_4442), .I1(n27_adj_4443), .I2(n26), 
            .I3(n28_adj_4444), .O(n37_adj_4445));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1578 (.I0(n37_adj_4445), .I1(n29_adj_4446), .I2(n36_adj_4441), 
            .I3(n30_adj_4447), .O(n15581));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_29001 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n34675));
    defparam bit_ctr_0__bdd_4_lut_29001.LUT_INIT = 16'he4aa;
    SB_LUT4 n34675_bdd_4_lut (.I0(n34675), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n32383));
    defparam n34675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i24686_2_lut (.I0(\state[1] ), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n30350));
    defparam i24686_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28355_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n29563));
    defparam i28355_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(one_wire_N_423[4]), .I1(one_wire_N_423[3]), 
            .I2(n29563), .I3(n26673), .O(n111));
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'h5155;
    SB_LUT4 bit_ctr_0__bdd_4_lut_28971 (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n34663));
    defparam bit_ctr_0__bdd_4_lut_28971.LUT_INIT = 16'he4aa;
    SB_LUT4 n34663_bdd_4_lut (.I0(n34663), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n32389));
    defparam n34663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n34500), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n34500), 
            .CO(n25730));
    SB_LUT4 bit_ctr_0__bdd_4_lut_28961 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n34609));
    defparam bit_ctr_0__bdd_4_lut_28961.LUT_INIT = 16'he4aa;
    SB_LUT4 n34609_bdd_4_lut (.I0(n34609), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n34612));
    defparam n34609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_28917 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n34597));
    defparam bit_ctr_0__bdd_4_lut_28917.LUT_INIT = 16'he4aa;
    SB_LUT4 n34597_bdd_4_lut (.I0(n34597), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n33801));
    defparam n34597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n16688), 
            .D(n255[6]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n24833), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n16688), 
            .D(n255[26]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_26 (.CI(n24833), .I0(bit_ctr[24]), .I1(GND_net), .CO(n24834));
    SB_CARRY add_21_12 (.CI(n24819), .I0(bit_ctr[10]), .I1(GND_net), .CO(n24820));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n24832), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_423[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n25030), .O(n22_adj_4439)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_423[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n25029), .O(n23_adj_4438)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n25029), .I0(timer[30]), .I1(n1[30]), 
            .CO(n25030));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_423[19]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n25028), .O(n28_adj_4444)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n16688), 
            .D(n255[25]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n24811), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_31 (.CI(n25028), .I0(timer[29]), .I1(n1[29]), 
            .CO(n25029));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_423[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n25027), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n25027), .I0(timer[28]), .I1(n1[28]), 
            .CO(n25028));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_423[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n25026), .O(n21_adj_4437)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n25026), .I0(timer[27]), .I1(n1[27]), 
            .CO(n25027));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n24818), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n25025), .O(one_wire_N_423[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_25 (.CI(n24832), .I0(bit_ctr[23]), .I1(GND_net), .CO(n24833));
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n16688), 
            .D(n255[12]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n16688), 
            .D(n255[11]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n16688), 
            .D(n255[24]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n16688), 
            .D(n255[23]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n16688), 
            .D(n255[10]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i1_4_lut_adj_1580 (.I0(n111), .I1(n29563), .I2(one_wire_N_423[2]), 
            .I3(one_wire_N_423[3]), .O(n116));
    defparam i1_4_lut_adj_1580.LUT_INIT = 16'haeee;
    SB_LUT4 i6_4_lut_adj_1581 (.I0(one_wire_N_423[8]), .I1(one_wire_N_423[10]), 
            .I2(n30350), .I3(n116), .O(n16_adj_4451));
    defparam i6_4_lut_adj_1581.LUT_INIT = 16'h0100;
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n16688), 
            .D(n255[9]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n16688), 
            .D(n255[22]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_28 (.CI(n25025), .I0(timer[26]), .I1(n1[26]), 
            .CO(n25026));
    SB_CARRY add_21_11 (.CI(n24818), .I0(bit_ctr[9]), .I1(GND_net), .CO(n24819));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n24831), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n25024), .O(one_wire_N_423[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_4 (.CI(n24811), .I0(bit_ctr[2]), .I1(GND_net), .CO(n24812));
    SB_CARRY add_21_24 (.CI(n24831), .I0(bit_ctr[22]), .I1(GND_net), .CO(n24832));
    SB_CARRY sub_14_add_2_27 (.CI(n25024), .I0(timer[25]), .I1(n1[25]), 
            .CO(n25025));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n24817), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n25023), .O(one_wire_N_423[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n24810), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_26 (.CI(n25023), .I0(timer[24]), .I1(n1[24]), 
            .CO(n25024));
    SB_CARRY add_21_10 (.CI(n24817), .I0(bit_ctr[8]), .I1(GND_net), .CO(n24818));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n24830), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n24816), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n24830), .I0(bit_ctr[21]), .I1(GND_net), .CO(n24831));
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n24829), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_22 (.CI(n24829), .I0(bit_ctr[20]), .I1(GND_net), .CO(n24830));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n24828), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_423[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n25022), .O(n30_adj_4447)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i24704_4_lut (.I0(n15471), .I1(n30348), .I2(n26419), .I3(\state[0] ), 
            .O(n30370));
    defparam i24704_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut_adj_1582 (.I0(n30370), .I1(\state[1] ), .I2(start), 
            .I3(\neo_pixel_transmitter.done ), .O(n7_adj_4454));
    defparam i20_4_lut_adj_1582.LUT_INIT = 16'hcfcd;
    SB_LUT4 i1_4_lut_adj_1583 (.I0(n22115), .I1(n7_adj_4454), .I2(n15574), 
            .I3(\state[1] ), .O(n28583));
    defparam i1_4_lut_adj_1583.LUT_INIT = 16'hccc4;
    SB_LUT4 i3_4_lut_4_lut (.I0(n30302), .I1(n14164), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n14164), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n30302), .O(n30427));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i3338_2_lut_3_lut (.I0(bit_ctr[29]), .I1(n22071), .I2(bit_ctr[28]), 
            .I3(GND_net), .O(n6706));
    defparam i3338_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i27732_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n22071), .I2(n30429), 
            .I3(bit_ctr[28]), .O(n30302));
    defparam i27732_3_lut_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 i17767_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n21867));   // verilog/neopixel.v(22[26:36])
    defparam i17767_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(n22071), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut.LUT_INIT = 16'hd222;
    SB_CARRY sub_14_add_2_25 (.CI(n25022), .I0(timer[23]), .I1(n1[23]), 
            .CO(n25023));
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n28495));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_24_lut (.I0(one_wire_N_423[13]), .I1(timer[22]), 
            .I2(n1[22]), .I3(n25021), .O(n24_adj_4440)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i8_3_lut_adj_1584 (.I0(one_wire_N_423[5]), .I1(n16_adj_4451), 
            .I2(n15581), .I3(GND_net), .O(n18_adj_4456));
    defparam i8_3_lut_adj_1584.LUT_INIT = 16'h0404;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n17366));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n17365));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n17364));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n17363));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n17362));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n17361));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n17360));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n17359));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n17358));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n17357));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n17356));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n17355));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n17354));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n17353));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n17352));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n17351));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n17350));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n17349));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n17348));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n17347));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n17346));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n17345));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_21 (.CI(n24828), .I0(bit_ctr[19]), .I1(GND_net), .CO(n24829));
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n17344));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n17343));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n17342));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n17341));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n17340));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n17339));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n17338));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n17337));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n17336));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n17316));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i24779_4_lut (.I0(n15471), .I1(n26419), .I2(n30348), .I3(\state[0] ), 
            .O(n22115));
    defparam i24779_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i17869_4_lut (.I0(one_wire_N_423[9]), .I1(n15581), .I2(one_wire_N_423[11]), 
            .I3(one_wire_N_423[10]), .O(n21971));
    defparam i17869_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF timer_1125__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n16688), 
            .D(n255[21]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n16688), 
            .D(n255[20]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i3_4_lut_adj_1585 (.I0(n9_adj_4369), .I1(one_wire_N_423[11]), 
            .I2(n18_adj_4456), .I3(one_wire_N_423[7]), .O(n34806));
    defparam i3_4_lut_adj_1585.LUT_INIT = 16'hffef;
    SB_LUT4 mux_589_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_480 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_589_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_CARRY sub_14_add_2_24 (.CI(n25021), .I0(timer[22]), .I1(n1[22]), 
            .CO(n25022));
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n16688), 
            .D(n255[19]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n16688), 
            .D(n255[18]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n16688), 
            .D(n255[17]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n25705), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n25704), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n16688), 
            .D(n255[16]), .R(n16807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_423[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n25020), .O(n25_adj_4442)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n16698), .D(state_3__N_272[0]), 
            .S(n30267));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_21 (.CI(n25704), .I0(n2391), .I1(n2423), .CO(n25705));
    SB_CARRY sub_14_add_2_23 (.CI(n25020), .I0(timer[21]), .I1(n1[21]), 
            .CO(n25021));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n25703), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n24827), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_20 (.CI(n25703), .I0(n2392), .I1(n2423), .CO(n25704));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n25702), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n25702), .I0(n2393), .I1(n2423), .CO(n25703));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n25701), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n25701), .I0(n2394), .I1(n2423), .CO(n25702));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n25700), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n25700), .I0(n2395), .I1(n2423), .CO(n25701));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n25699), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n25699), .I0(n2396), .I1(n2423), .CO(n25700));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n25698), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n25698), .I0(n2397), .I1(n2423), .CO(n25699));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n25697), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_423[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n25019), .O(n29_adj_4446)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1674_14 (.CI(n25697), .I0(n2398), .I1(n2423), .CO(n25698));
    SB_CARRY sub_14_add_2_22 (.CI(n25019), .I0(timer[20]), .I1(n1[20]), 
            .CO(n25020));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n25018), .O(one_wire_N_423[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_21 (.CI(n25018), .I0(timer[19]), .I1(n1[19]), 
            .CO(n25019));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n25017), .O(one_wire_N_423[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n25017), .I0(timer[18]), .I1(n1[18]), 
            .CO(n25018));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_423[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n25016), .O(n27_adj_4443)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_20 (.CI(n24827), .I0(bit_ctr[18]), .I1(GND_net), .CO(n24828));
    SB_CARRY sub_14_add_2_19 (.CI(n25016), .I0(timer[17]), .I1(n1[17]), 
            .CO(n25017));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n30475), .D(\neo_pixel_transmitter.done_N_486 ), 
            .R(n32089));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_DFF timer_1125__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n25015), .O(one_wire_N_423[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF timer_1125__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1125__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY sub_14_add_2_18 (.CI(n25015), .I0(timer[16]), .I1(n1[16]), 
            .CO(n25016));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n24826), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n25014), .O(one_wire_N_423[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_17 (.CI(n25014), .I0(timer[15]), .I1(n1[15]), 
            .CO(n25015));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n25013), .O(one_wire_N_423[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_19 (.CI(n24826), .I0(bit_ctr[17]), .I1(GND_net), .CO(n24827));
    SB_CARRY sub_14_add_2_16 (.CI(n25013), .I0(timer[14]), .I1(n1[14]), 
            .CO(n25014));
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n16852));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n25012), .O(one_wire_N_423[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_15 (.CI(n25012), .I0(timer[13]), .I1(n1[13]), 
            .CO(n25013));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n25011), .O(one_wire_N_423[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_14 (.CI(n25011), .I0(timer[12]), .I1(n1[12]), 
            .CO(n25012));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4), .I1(n4), .I2(n1037), .I3(n25880), 
            .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n25879), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n25879), .I0(n1005), .I1(n1037), .CO(n25880));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n25878), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17969_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n22071));   // verilog/neopixel.v(22[26:36])
    defparam i17969_2_lut_3_lut.LUT_INIT = 16'h6464;
    SB_CARRY mod_5_add_736_6 (.CI(n25878), .I0(n1006), .I1(n1037), .CO(n25879));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n25877), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n25877), .I0(n1007), .I1(n1037), .CO(n25878));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n25876), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n25876), .I0(n1008), .I1(n1037), .CO(n25877));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n34504), 
            .I3(n25875), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n25875), .I0(n1009), .I1(n34504), .CO(n25876));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n34504), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n34504), 
            .CO(n25875));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n25874), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n25873), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n25873), .I0(n1401), .I1(n1433), .CO(n25874));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n25872), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n25872), .I0(n1402), .I1(n1433), .CO(n25873));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n25871), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n25871), .I0(n1403), .I1(n1433), .CO(n25872));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n25870), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n25870), .I0(n1404), .I1(n1433), .CO(n25871));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n25869), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n25869), .I0(n1405), .I1(n1433), .CO(n25870));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n25868), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n25868), .I0(n1406), .I1(n1433), .CO(n25869));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n25867), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n25867), .I0(n1407), .I1(n1433), .CO(n25868));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n25866), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n25866), .I0(n1408), .I1(n1433), .CO(n25867));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n34505), 
            .I3(n25865), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n25865), .I0(n1409), .I1(n34505), .CO(n25866));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n34505), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n34505), 
            .CO(n25865));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n25864), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n25863), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n25863), .I0(n1500), .I1(n1532), .CO(n25864));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n25862), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n25862), .I0(n1501), .I1(n1532), .CO(n25863));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n25861), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n25861), .I0(n1502), .I1(n1532), .CO(n25862));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n25860), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n24825), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_9 (.CI(n25860), .I0(n1503), .I1(n1532), .CO(n25861));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n25859), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n25859), .I0(n1504), .I1(n1532), .CO(n25860));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n25858), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n25858), .I0(n1505), .I1(n1532), .CO(n25859));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n25010), .O(one_wire_N_423[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n25857), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_18 (.CI(n24825), .I0(bit_ctr[16]), .I1(GND_net), .CO(n24826));
    SB_CARRY mod_5_add_1071_6 (.CI(n25857), .I0(n1506), .I1(n1532), .CO(n25858));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n25856), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n25856), .I0(n1507), .I1(n1532), .CO(n25857));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n25855), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n25855), .I0(n1508), .I1(n1532), .CO(n25856));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n34506), 
            .I3(n25854), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_3 (.CI(n25854), .I0(n1509), .I1(n34506), .CO(n25855));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n34506), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n34506), 
            .CO(n25854));
    SB_CARRY sub_14_add_2_13 (.CI(n25010), .I0(timer[11]), .I1(n1[11]), 
            .CO(n25011));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n25853), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n25852), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n25852), .I0(n1599), .I1(n1631), .CO(n25853));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n25851), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n25851), .I0(n1600), .I1(n1631), .CO(n25852));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n25850), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n25850), .I0(n1601), .I1(n1631), .CO(n25851));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n25849), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n25849), .I0(n1602), .I1(n1631), .CO(n25850));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n25848), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n25009), .O(one_wire_N_423[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_9 (.CI(n25848), .I0(n1603), .I1(n1631), .CO(n25849));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n25847), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n25847), .I0(n1604), .I1(n1631), .CO(n25848));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n25846), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n25846), .I0(n1605), .I1(n1631), .CO(n25847));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n25845), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n25845), .I0(n1606), .I1(n1631), .CO(n25846));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n25844), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n25844), .I0(n1607), .I1(n1631), .CO(n25845));
    SB_CARRY sub_14_add_2_12 (.CI(n25009), .I0(timer[10]), .I1(n1[10]), 
            .CO(n25010));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n25843), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n25843), .I0(n1608), .I1(n1631), .CO(n25844));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n34507), 
            .I3(n25842), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n24824), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_3 (.CI(n25842), .I0(n1609), .I1(n34507), .CO(n25843));
    SB_CARRY add_21_9 (.CI(n24816), .I0(bit_ctr[7]), .I1(GND_net), .CO(n24817));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n34507), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n34507), 
            .CO(n25842));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n25841), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n25840), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n25840), .I0(n1698), .I1(n1730), .CO(n25841));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n25839), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n24815), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_13 (.CI(n25839), .I0(n1699), .I1(n1730), .CO(n25840));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n25838), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n25838), .I0(n1700), .I1(n1730), .CO(n25839));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n25837), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n25837), .I0(n1701), .I1(n1730), .CO(n25838));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n25836), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n25836), .I0(n1702), .I1(n1730), .CO(n25837));
    SB_CARRY add_21_17 (.CI(n24824), .I0(bit_ctr[15]), .I1(GND_net), .CO(n24825));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n25835), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n25835), .I0(n1703), .I1(n1730), .CO(n25836));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n25834), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n25834), .I0(n1704), .I1(n1730), .CO(n25835));
    SB_CARRY add_21_3 (.CI(n24810), .I0(bit_ctr[1]), .I1(GND_net), .CO(n24811));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n25833), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n25833), .I0(n1705), .I1(n1730), .CO(n25834));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n25008), .O(one_wire_N_423[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n25832), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n25832), .I0(n1706), .I1(n1730), .CO(n25833));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n25831), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n25831), .I0(n1707), .I1(n1730), .CO(n25832));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n25830), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n25830), .I0(n1708), .I1(n1730), .CO(n25831));
    SB_CARRY sub_14_add_2_11 (.CI(n25008), .I0(timer[9]), .I1(n1[9]), 
            .CO(n25009));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n34508), 
            .I3(n25829), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n25007), .O(one_wire_N_423[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_3 (.CI(n25829), .I0(n1709), .I1(n34508), .CO(n25830));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n34508), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_10 (.CI(n25007), .I0(timer[8]), .I1(n1[8]), 
            .CO(n25008));
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n34508), 
            .CO(n25829));
    SB_LUT4 i27737_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n30429), .I2(bit_ctr[27]), 
            .I3(n838), .O(n16727));
    defparam i27737_3_lut_4_lut.LUT_INIT = 16'h6696;
    SB_CARRY add_21_8 (.CI(n24815), .I0(bit_ctr[6]), .I1(GND_net), .CO(n24816));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n25828), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n25827), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n25827), .I0(n1797), .I1(n1829), .CO(n25828));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n25826), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n25826), .I0(n1798), .I1(n1829), .CO(n25827));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n25006), .O(one_wire_N_423[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n25825), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n25825), .I0(n1799), .I1(n1829), .CO(n25826));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n24823), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n25824), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_16 (.CI(n24823), .I0(bit_ctr[14]), .I1(GND_net), .CO(n24824));
    SB_CARRY mod_5_add_1272_12 (.CI(n25824), .I0(n1800), .I1(n1829), .CO(n25825));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n25823), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n25823), .I0(n1801), .I1(n1829), .CO(n25824));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n25822), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n25822), .I0(n1802), .I1(n1829), .CO(n25823));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n25821), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n25821), .I0(n1803), .I1(n1829), .CO(n25822));
    SB_CARRY sub_14_add_2_9 (.CI(n25006), .I0(timer[7]), .I1(n1[7]), .CO(n25007));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n25820), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_423[9]), .I1(timer[6]), .I2(n1[6]), 
            .I3(n25005), .O(n9_adj_4369)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1272_8 (.CI(n25820), .I0(n1804), .I1(n1829), .CO(n25821));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n25819), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n25819), .I0(n1805), .I1(n1829), .CO(n25820));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n25818), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n25818), .I0(n1806), .I1(n1829), .CO(n25819));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n25817), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_5 (.CI(n25817), .I0(n1807), .I1(n1829), .CO(n25818));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n25816), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n25816), .I0(n1808), .I1(n1829), .CO(n25817));
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n24814), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n34509), 
            .I3(n25815), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n25815), .I0(n1809), .I1(n34509), .CO(n25816));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n34509), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n34509), 
            .CO(n25815));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n25814), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n25813), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n25813), .I0(n1896), .I1(n1928), .CO(n25814));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n25812), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n25812), .I0(n1897), .I1(n1928), .CO(n25813));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n24822), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n25811), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n25811), .I0(n1898), .I1(n1928), .CO(n25812));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n25810), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n25810), .I0(n1899), .I1(n1928), .CO(n25811));
    SB_CARRY sub_14_add_2_8 (.CI(n25005), .I0(timer[6]), .I1(n1[6]), .CO(n25006));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n25809), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n25809), .I0(n1900), .I1(n1928), .CO(n25810));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n25808), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n25808), .I0(n1901), .I1(n1928), .CO(n25809));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n25807), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n25807), .I0(n1902), .I1(n1928), .CO(n25808));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n25806), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n25806), .I0(n1903), .I1(n1928), .CO(n25807));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n25805), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_15 (.CI(n24822), .I0(bit_ctr[13]), .I1(GND_net), .CO(n24823));
    SB_CARRY mod_5_add_1339_8 (.CI(n25805), .I0(n1904), .I1(n1928), .CO(n25806));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n25804), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n25804), .I0(n1905), .I1(n1928), .CO(n25805));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n25803), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n25803), .I0(n1906), .I1(n1928), .CO(n25804));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n25802), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n25802), .I0(n1907), .I1(n1928), .CO(n25803));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n25801), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n24810));
    SB_CARRY mod_5_add_1339_4 (.CI(n25801), .I0(n1908), .I1(n1928), .CO(n25802));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n34510), 
            .I3(n25800), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_3 (.CI(n25800), .I0(n1909), .I1(n34510), .CO(n25801));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n34510), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n34510), 
            .CO(n25800));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n25799), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n25798), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n25798), .I0(n1995), .I1(n2027), .CO(n25799));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n25797), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_7 (.CI(n24814), .I0(bit_ctr[5]), .I1(GND_net), .CO(n24815));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n24813), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n24821), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_16 (.CI(n25797), .I0(n1996), .I1(n2027), .CO(n25798));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n25796), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n25796), .I0(n1997), .I1(n2027), .CO(n25797));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n25795), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n25795), .I0(n1998), .I1(n2027), .CO(n25796));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n25794), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n25794), .I0(n1999), .I1(n2027), .CO(n25795));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n25793), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n25793), .I0(n2000), .I1(n2027), .CO(n25794));
    SB_CARRY add_21_14 (.CI(n24821), .I0(bit_ctr[12]), .I1(GND_net), .CO(n24822));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n25792), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n25792), .I0(n2001), .I1(n2027), .CO(n25793));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n25791), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n25791), .I0(n2002), .I1(n2027), .CO(n25792));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n25790), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_6 (.CI(n24813), .I0(bit_ctr[4]), .I1(GND_net), .CO(n24814));
    SB_CARRY mod_5_add_1406_9 (.CI(n25790), .I0(n2003), .I1(n2027), .CO(n25791));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n25789), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n25789), .I0(n2004), .I1(n2027), .CO(n25790));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n25788), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n25788), .I0(n2005), .I1(n2027), .CO(n25789));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n25787), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n25787), .I0(n2006), .I1(n2027), .CO(n25788));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n25786), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_5 (.CI(n25786), .I0(n2007), .I1(n2027), .CO(n25787));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n25785), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n25785), .I0(n2008), .I1(n2027), .CO(n25786));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n34511), 
            .I3(n25784), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_3 (.CI(n25784), .I0(n2009), .I1(n34511), .CO(n25785));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n34511), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n34511), 
            .CO(n25784));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n25783), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n25782), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n25782), .I0(n2094), .I1(n2126), .CO(n25783));
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n34516), .I2(n32383), 
            .I3(n35413), .O(n34525));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n34525_bdd_4_lut (.I0(n34525), .I1(n33801), .I2(n32389), .I3(n35413), 
            .O(n34528));
    defparam n34525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_28908 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n34513));
    defparam bit_ctr_0__bdd_4_lut_28908.LUT_INIT = 16'he4aa;
    SB_LUT4 n34513_bdd_4_lut (.I0(n34513), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n34516));
    defparam n34513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i28837_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34511));
    defparam i28837_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i27780_3_lut_4_lut (.I0(n26419), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n15471), .O(n33174));
    defparam i27780_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_272[1] ), .O(n16807));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i27818_3_lut_4_lut (.I0(n15471), .I1(n33493), .I2(\state[1] ), 
            .I3(start), .O(n33494));
    defparam i27818_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1586 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4463));
    defparam i2_2_lut_adj_1586.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1587 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4464));
    defparam i12_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1588 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4465));
    defparam i10_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1589 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4466));
    defparam i11_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1590 (.I0(bit_ctr[15]), .I1(n18_adj_4463), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4467));
    defparam i9_4_lut_adj_1590.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1591 (.I0(n25_adj_4467), .I1(n27_adj_4466), .I2(n26_adj_4465), 
            .I3(n28_adj_4464), .O(n2027));
    defparam i15_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i28836_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34510));
    defparam i28836_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut_adj_1592 (.I0(n21971), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n32089));
    defparam i3_4_lut_4_lut_adj_1592.LUT_INIT = 16'h0004;
    SB_LUT4 i11_4_lut_adj_1593 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4468));
    defparam i11_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), .I3(GND_net), 
            .O(n19_adj_4469));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1594 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4470));
    defparam i1_2_lut_adj_1594.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1595 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4471));
    defparam i9_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1596 (.I0(n19_adj_4469), .I1(n26_adj_4468), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4472));
    defparam i13_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1597 (.I0(n1896), .I1(n28_adj_4472), .I2(n24_adj_4471), 
            .I3(n16_adj_4470), .O(n1928));
    defparam i14_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i28835_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34509));
    defparam i28835_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1598 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_4473));
    defparam i10_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1599 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_4474));
    defparam i8_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1600 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_4475));
    defparam i9_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1601 (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_4476));
    defparam i7_3_lut_adj_1601.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1602 (.I0(n21_adj_4476), .I1(n23_adj_4475), .I2(n22_adj_4474), 
            .I3(n24_adj_4473), .O(n1829));
    defparam i13_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28834_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34508));
    defparam i28834_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1603 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_4477));
    defparam i4_3_lut_adj_1603.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1604 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4478));
    defparam i8_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1605 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4479));
    defparam i7_3_lut_adj_1605.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1606 (.I0(n21_adj_4478), .I1(n17_adj_4477), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4480));
    defparam i11_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1607 (.I0(n1700), .I1(n24_adj_4480), .I2(n20_adj_4479), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i28833_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34507));
    defparam i28833_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1608 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4481));
    defparam i8_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1609 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4482));
    defparam i1_3_lut_adj_1609.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4483));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1610 (.I0(n13_adj_4482), .I1(n20_adj_4481), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4484));
    defparam i10_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1611 (.I0(n1601), .I1(n22_adj_4484), .I2(n18_adj_4483), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i28832_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34506));
    defparam i28832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1612 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4485));
    defparam i7_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1613 (.I0(n1504), .I1(n18_adj_4485), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4486));
    defparam i9_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1614 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4487));
    defparam i4_3_lut_adj_1614.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1615 (.I0(n15_adj_4487), .I1(n20_adj_4486), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i28831_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34505));
    defparam i28831_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (data_o, GND_net, encoder1_position, 
            clk32MHz, n32056, reg_B, ENCODER1_A_c_1, VCC_net, n16872, 
            ENCODER1_B_c_0, n17382) /* synthesis syn_module_defined=1 */ ;
    output [1:0]data_o;
    input GND_net;
    output [23:0]encoder1_position;
    input clk32MHz;
    output n32056;
    output [1:0]reg_B;
    input ENCODER1_A_c_1;
    input VCC_net;
    input n16872;
    input ENCODER1_B_c_0;
    input n17382;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire B_delayed, count_direction, A_delayed, count_enable;
    wire [23:0]n2499;
    
    wire n2476, n24999, n24998, n24997, n24996, n24995, n24994, 
        n24993, n24992, n24991, n24990, n24989, n24988, n24987, 
        n24986, n24985, n24984, n24983, n24982, n24981, n24980, 
        n24979, n24978, n24977, n24976;
    
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2499[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_529_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2476), 
            .I3(n24999), .O(n2499[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_529_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2476), 
            .I3(n24998), .O(n2499[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_24 (.CI(n24998), .I0(encoder1_position[22]), .I1(n2476), 
            .CO(n24999));
    SB_LUT4 add_529_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2476), 
            .I3(n24997), .O(n2499[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_23 (.CI(n24997), .I0(encoder1_position[21]), .I1(n2476), 
            .CO(n24998));
    SB_LUT4 add_529_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2476), 
            .I3(n24996), .O(n2499[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_22 (.CI(n24996), .I0(encoder1_position[20]), .I1(n2476), 
            .CO(n24997));
    SB_LUT4 add_529_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2476), 
            .I3(n24995), .O(n2499[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_21 (.CI(n24995), .I0(encoder1_position[19]), .I1(n2476), 
            .CO(n24996));
    SB_LUT4 add_529_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2476), 
            .I3(n24994), .O(n2499[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_20 (.CI(n24994), .I0(encoder1_position[18]), .I1(n2476), 
            .CO(n24995));
    SB_LUT4 add_529_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2476), 
            .I3(n24993), .O(n2499[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_19 (.CI(n24993), .I0(encoder1_position[17]), .I1(n2476), 
            .CO(n24994));
    SB_LUT4 add_529_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2476), 
            .I3(n24992), .O(n2499[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_18 (.CI(n24992), .I0(encoder1_position[16]), .I1(n2476), 
            .CO(n24993));
    SB_LUT4 add_529_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2476), 
            .I3(n24991), .O(n2499[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_17 (.CI(n24991), .I0(encoder1_position[15]), .I1(n2476), 
            .CO(n24992));
    SB_LUT4 add_529_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2476), 
            .I3(n24990), .O(n2499[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_16 (.CI(n24990), .I0(encoder1_position[14]), .I1(n2476), 
            .CO(n24991));
    SB_LUT4 add_529_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2476), 
            .I3(n24989), .O(n2499[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_15 (.CI(n24989), .I0(encoder1_position[13]), .I1(n2476), 
            .CO(n24990));
    SB_LUT4 add_529_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2476), 
            .I3(n24988), .O(n2499[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_14 (.CI(n24988), .I0(encoder1_position[12]), .I1(n2476), 
            .CO(n24989));
    SB_LUT4 add_529_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2476), 
            .I3(n24987), .O(n2499[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_13 (.CI(n24987), .I0(encoder1_position[11]), .I1(n2476), 
            .CO(n24988));
    SB_LUT4 add_529_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2476), 
            .I3(n24986), .O(n2499[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_12 (.CI(n24986), .I0(encoder1_position[10]), .I1(n2476), 
            .CO(n24987));
    SB_LUT4 add_529_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2476), 
            .I3(n24985), .O(n2499[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_11 (.CI(n24985), .I0(encoder1_position[9]), .I1(n2476), 
            .CO(n24986));
    SB_LUT4 add_529_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2476), 
            .I3(n24984), .O(n2499[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_10 (.CI(n24984), .I0(encoder1_position[8]), .I1(n2476), 
            .CO(n24985));
    SB_LUT4 add_529_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2476), 
            .I3(n24983), .O(n2499[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_9 (.CI(n24983), .I0(encoder1_position[7]), .I1(n2476), 
            .CO(n24984));
    SB_LUT4 add_529_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2476), 
            .I3(n24982), .O(n2499[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_8 (.CI(n24982), .I0(encoder1_position[6]), .I1(n2476), 
            .CO(n24983));
    SB_LUT4 add_529_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2476), 
            .I3(n24981), .O(n2499[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_7 (.CI(n24981), .I0(encoder1_position[5]), .I1(n2476), 
            .CO(n24982));
    SB_LUT4 add_529_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2476), 
            .I3(n24980), .O(n2499[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_6 (.CI(n24980), .I0(encoder1_position[4]), .I1(n2476), 
            .CO(n24981));
    SB_LUT4 add_529_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2476), 
            .I3(n24979), .O(n2499[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_5 (.CI(n24979), .I0(encoder1_position[3]), .I1(n2476), 
            .CO(n24980));
    SB_LUT4 add_529_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2476), 
            .I3(n24978), .O(n2499[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_4 (.CI(n24978), .I0(encoder1_position[2]), .I1(n2476), 
            .CO(n24979));
    SB_LUT4 add_529_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2476), 
            .I3(n24977), .O(n2499[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_3 (.CI(n24977), .I0(encoder1_position[1]), .I1(n2476), 
            .CO(n24978));
    SB_LUT4 add_529_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n24976), .O(n2499[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_529_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_529_2 (.CI(n24976), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n24977));
    SB_CARRY add_529_1 (.CI(GND_net), .I0(n2476), .I1(n2476), .CO(n24976));
    SB_LUT4 i863_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2476));   // quad.v(37[5] 40[8])
    defparam i863_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,100)  debounce (.n32056(n32056), .reg_B({reg_B}), .GND_net(GND_net), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .n16872(n16872), .data_o({data_o}), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n17382(n17382));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (n32056, reg_B, GND_net, ENCODER1_A_c_1, 
            clk32MHz, VCC_net, n16872, data_o, ENCODER1_B_c_0, n17382);
    output n32056;
    output [1:0]reg_B;
    input GND_net;
    input ENCODER1_A_c_1;
    input clk32MHz;
    input VCC_net;
    input n16872;
    output [1:0]data_o;
    input ENCODER1_B_c_0;
    input n17382;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3600;
    wire [6:0]n33;
    
    wire n25588, n25587, n25586, n25585, n25584, n25583;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n32056));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n32056), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1132_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n25588), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1132_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1132_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n25587), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1132_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1132_add_4_7 (.CI(n25587), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n25588));
    SB_LUT4 cnt_reg_1132_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n25586), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1132_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1132_add_4_6 (.CI(n25586), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n25587));
    SB_LUT4 cnt_reg_1132_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n25585), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1132_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1132_add_4_5 (.CI(n25585), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n25586));
    SB_LUT4 cnt_reg_1132_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n25584), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1132_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1132_add_4_4 (.CI(n25584), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n25585));
    SB_LUT4 cnt_reg_1132_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n25583), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1132_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1132_add_4_3 (.CI(n25583), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n25584));
    SB_LUT4 cnt_reg_1132_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1132_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1132_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n25583));
    SB_DFFSR cnt_reg_1132__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n16872));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n17382));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1132__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1132__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1132__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1132__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1132__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1132__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3600));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[2] , GND_net, \Kp[0] , \Kp[1] , \Kp[3] , 
            \Kp[6] , \Kp[4] , \Ki[8] , \Kp[5] , \Ki[1] , \Ki[0] , 
            \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , \Ki[6] , \Ki[7] , 
            \Ki[9] , \Ki[10] , \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , 
            \Ki[15] , PWMLimit, IntegralLimit, \Kp[7] , \Kp[8] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[15] , 
            n29, \duty_23__N_3516[14] , duty, clk32MHz, setpoint, 
            motor_state, n34501, VCC_net, n18701) /* synthesis syn_module_defined=1 */ ;
    input \Kp[2] ;
    input GND_net;
    input \Kp[0] ;
    input \Kp[1] ;
    input \Kp[3] ;
    input \Kp[6] ;
    input \Kp[4] ;
    input \Ki[8] ;
    input \Kp[5] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input [23:0]PWMLimit;
    input [23:0]IntegralLimit;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input n29;
    output \duty_23__N_3516[14] ;
    output [23:0]duty;
    input clk32MHz;
    input [23:0]setpoint;
    input [23:0]motor_state;
    output n34501;
    input VCC_net;
    input n18701;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    
    wire n204, n24918;
    wire [47:0]n106;
    wire [47:0]n155;
    
    wire n24919;
    wire [1:0]n8422;
    
    wire n24855;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    wire [23:0]n2629;
    
    wire n24856, n24846, n24847, n4_adj_3913;
    wire [2:0]n8417;
    wire [3:0]n8411;
    
    wire n490, n12, n6_adj_3914, n8_adj_3915, n11, n6_adj_3916;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3416 ;
    
    wire n621, n24650, n18, n13, n4_adj_3917, n30955, n77, n8_adj_3918, 
        n150, n223, n296, n369, n442, n515, n588, n661, n734, 
        n807, n880, n953, n1026, n1099, n530, n603, \PID_CONTROLLER.integral_23__N_3464 , 
        n676, n749, n822, n895, n968, n1041, n1114, n95, n26, 
        n168, n241, n314, n387, n460, n533, n606, n679, n752, 
        n825, n898;
    wire [23:0]n1_adj_4337;
    
    wire n77_adj_3921, n8_adj_3922, n150_adj_3924, n223_adj_3925, n74, 
        n5_adj_3927, n147, n220, n293, n296_adj_3928, n366, n439, 
        n512, n585, n658, n731, n369_adj_3929, n804, n877, n950, 
        n1023;
    wire [5:0]n8693;
    
    wire n31043, n490_adj_3930, n26372;
    wire [4:0]n8701;
    
    wire n417, n26371, n344, n26370, n271, n26369, n198, n26368, 
        n56, n125;
    wire [6:0]n8684;
    
    wire n560, n26367, n487, n26366, n414, n26365, n341, n26364, 
        n268, n26363, n195, n26362, n53, n122;
    wire [7:0]n8674;
    
    wire n630, n26361, n557, n26360, n484, n26359, n411, n26358, 
        n338, n26357, n265, n26356, n192, n26355, n50, n119;
    wire [8:0]n8663;
    
    wire n700, n26354, n627, n26353, n554, n26352, n481, n26351, 
        n408, n26350, n335, n26349, n262, n26348, n189, n26347, 
        n47, n116;
    wire [9:0]n8651;
    
    wire n770, n26346, n697, n26345, n1096, n971, n624, n26344, 
        n1044, n442_adj_3932, n551, n26343, n35222, n33677, n33675, 
        n478, n26342, n1117, n405, n26341, n332, n26340, n98, 
        n29_c, n171, n244, n317, n390, n463, n80, n11_adj_3934;
    wire [23:0]duty_23__N_3516;
    
    wire n24917, n536, n609, n153, n226, n299, n372, n682, n445, 
        n259, n26339, n518;
    wire [23:0]n257;
    
    wire n256;
    wire [23:0]duty_23__N_3491;
    
    wire duty_23__N_3515;
    wire [23:0]duty_23__N_3392;
    
    wire n515_adj_3935, n755, n591, n588_adj_3936, n186_adj_3937, 
        n26338, n664, n661_adj_3938, n737, n810, n883, n956, n24845, 
        n1029, n1102, n83, n14_adj_3939, n734_adj_3940, n156, n229, 
        n807_adj_3941, n302, n375, n448, n521, n594, n667, n740, 
        n35216, n880_adj_3942, n813, n886, n959, n1032, n953_adj_3943, 
        n1026_adj_3944, n44, n113, n828, n901, n974, n1099_adj_3945, 
        n1047;
    wire [10:0]n8638;
    
    wire n840, n26337, n1105, n1120, n767, n26336, n86, n17_adj_3946, 
        n101, n694, n26335, n32, n174, n247, n320, n393, n466, 
        n539, n612, n685, n758, n831, n904, n977, n1050, n104, 
        n35, n177, n250, n27, n15_adj_3948, n13_adj_3949, n11_adj_3950, 
        n33357, n323, n396, n469, n542, n615, n688, n761, n834, 
        n41, n39, n45, n26334, n37, n31, n43, n548, n26333, 
        n475, n26332, n23_adj_3951, n402, n26331, n329, n26330, 
        n25_adj_3952, n256_adj_3953, n26329, n183, n26328, n41_adj_3954, 
        n110;
    wire [11:0]n8624;
    
    wire n910, n26327, n35_adj_3955, n837, n26326, n11_adj_3956, 
        n13_adj_3957, n15_adj_3958, n27_adj_3959, n764, n26325, n33, 
        n691, n26324, n9_adj_3960, n17_adj_3961, n618, n26323, n19, 
        n21, n545, n26322, n33321, n33315, n12_adj_3962, n472, 
        n26321, n399, n26320, n10, n30, n326, n26319, n33331, 
        n33603, n33599, n33909, n33751, n33962, n16_adj_3964, n6_adj_3965, 
        n33895, n33896, n8_adj_3966, n24_adj_3967, n33301, n33299, 
        n33769, n24854, n33836, n4_adj_3968, n33885, n33886, n33311, 
        n33309, n33972, n33838, n34021, n34022, n34003, n33303, 
        n33925, n40, n33927, n24916;
    wire [23:0]n1_adj_4338;
    
    wire n24844, n39_adj_3971, n41_adj_3972, n45_adj_3974, n43_adj_3975, 
        n37_adj_3976, n29_adj_3977, n31_adj_3978, n23_adj_3979, n25_adj_3980, 
        n35_adj_3981, n33_adj_3983, n253, n26318, n11_adj_3984, n13_adj_3985, 
        n15_adj_3986, n27_adj_3988, n9_adj_3989, n17_adj_3990, n19_adj_3991, 
        n21_adj_3993, n33285, n33278, n12_adj_3994, n10_adj_3995, 
        n30_adj_3996, n33296, n33570, n33566, n33901, n33735, n33960, 
        n16_adj_3997, n6_adj_3998, n33881, n33882, n8_adj_3999, n24_adj_4000, 
        n33263, n33261, n33771, n33842, n4_adj_4001, n33879, n33880, 
        n33274, n33272, n33974, n33844, n34023, n34024, n34001, 
        n33265, n33931, n40_adj_4002, n33933, n907, n980, n107, 
        n38, n180, n26317;
    wire [12:0]n8609;
    
    wire n26316, n26315, n26314, n26313, n26312, n26311, n26310, 
        n26309, n26308, n26307, n21_adj_4005, n19_adj_4006, n17_adj_4007, 
        n9_adj_4008, n33366, n26306, n26305;
    wire [13:0]n8593;
    
    wire n26304, n26303, n26302, n43_adj_4009, n16_adj_4010, n33333, 
        n26301, n26300, n26299, n26298, n26297, n24843, n8_adj_4011, 
        n26296, n26295, n24853, n26294, n26293, n74_adj_4014, n5_adj_4015, 
        n147_adj_4016, n220_adj_4017, n293_adj_4018, n366_adj_4019, 
        n439_adj_4020, n512_adj_4022, n585_adj_4024, n658_adj_4025, 
        n731_adj_4027, n804_adj_4028, n26292, n877_adj_4031;
    wire [14:0]n8576;
    
    wire n26291, n950_adj_4032, n1023_adj_4033, n1096_adj_4034, n45_adj_4035, 
        n24_adj_4036, n26290, n80_adj_4037, n26289, n11_adj_4038, 
        n153_adj_4039, n226_adj_4040, n299_adj_4041, n372_adj_4042, 
        n445_adj_4043, n518_adj_4044, n26288, n591_adj_4045, n24915, 
        n664_adj_4047, n737_adj_4048, n810_adj_4049, n6_adj_4050;
    wire [3:0]n8708;
    
    wire n204_adj_4051;
    wire [1:0]n8719;
    
    wire n26287, n131, n62, n7_adj_4052, n5_adj_4053, n33398, n33650, 
        n33646, n25_adj_4054, n23_adj_4055, n33937, n31_adj_4056, 
        n29_adj_4057, n33777, n37_adj_4058, n35_adj_4059, n33_adj_4060, 
        n33964, n35239, n11_adj_4061, n33681, n35209, n33669, n26286, 
        n4_adj_4062;
    wire [2:0]n8714;
    
    wire n26285, n12_adj_4063, n8_adj_4064, n26284, n26283, n26282, 
        n26281, n11_adj_4065, n26280, n26279, n26278, n6_adj_4066;
    wire [15:0]n8558;
    
    wire n26277, n26276, n26275, n24914, n24782, n26274, n24852, 
        n18_adj_4067, n13_adj_4068, n4_adj_4069, n26273, n26272, n26271, 
        n26270, n26269, n26268, n26267, n26266, n26265, n26264, 
        n24913, n26263;
    wire [16:0]n8539;
    
    wire n26262, n25053, n26261, n24851, n24842, n25052, n24850, 
        n24841, n24912, n26260, n26259, n26258, n26257, n26256, 
        n26255, n26254, n24849, n26253, n26252, n457, n26251, 
        n25051, n883_adj_4072, n956_adj_4073, n35204, n12_adj_4074, 
        n1029_adj_4075, n33414, n35227, n10_adj_4076, n30_adj_4077, 
        n33679, n33865, n1102_adj_4078, n384, n26250, n33422, n83_adj_4079, 
        n311, n26249, n24848, n238, n26248, n165, n26247, n23_adj_4080, 
        n92, n14_adj_4081, n156_adj_4082, n229_adj_4083, n302_adj_4084, 
        n159, n375_adj_4085, n448_adj_4086, n232, n521_adj_4087, n305, 
        n378, n451, n524, n594_adj_4089, n667_adj_4090, n597, n740_adj_4091, 
        n813_adj_4093, n886_adj_4094, n959_adj_4095, n1032_adj_4096, 
        n1105_adj_4097, n670, n743, n816, n889;
    wire [17:0]n8519;
    
    wire n26246, n24911, n25050, n25049, n26245, n25048, n26244, 
        n962, n1035, n1108, n35207, n24910, n89, n20_adj_4104, 
        n24909, n33793, n1111, n26243, n35233, n162, n25047, n235, 
        n308, n1038, n26242, n965, n26241, n892, n26240, n819, 
        n26239, n746, n26238, n673, n26237, n600, n26236, n24908, 
        n33942, n381, n527, n26235, n454, n26234, n25122, n25121, 
        n26233, n25120, n26232, n26231, n26230, n25046;
    wire [18:0]n8498;
    
    wire n26229, n26228, n26227, n26226, n26225, n26224, n26223, 
        n25119, n25118, n25117, n25116, n25045, n25115, n35198, 
        n33996, n35195, n16_adj_4111, n33400, n24_adj_4112, n6_adj_4113, 
        n33813, n33814, n33402, n8_adj_4114, n35193, n33765, n33620;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3467 ;
    
    wire n3_adj_4115, n4_adj_4116, n33805, n33806, n12_adj_4117, n33345, 
        n10_adj_4118, n30_adj_4119, n26222, n25114, n26221, n26220, 
        n26219, n25113, n26218, n26217, n25112, n24907, n26216, 
        n26215, n26214, n26213, n26212, n24625, n33351, n33970, 
        n33633, n34019, n34020, n39_adj_4121, n34005, n6_adj_4122, 
        n33831, n33832, n33335, n33767;
    wire [19:0]n8476;
    
    wire n26211, n26210, n26209, n26208, n26207, n25044, n26206, 
        n33440, n33631, n41_adj_4124, n33337, n33919, n26205, n26204, 
        n40_adj_4125, n33921, n4_adj_4126, n33811, n26203, n33812, 
        n33416, n33954, n33622, n34006, n26202, n34007, n33981, 
        n33407, n33915, n33628, \PID_CONTROLLER.integral_23__N_3466 , 
        n33966, n25043, n26201, n25042, n26200, n26199, n26198, 
        n26197, n26196, n26195, n26194, n26193;
    wire [20:0]n8453;
    
    wire n26192, n26191, n26190, n26189, n26188, n26187, n26186, 
        n26185, n26184, n26183, n26182, n26181, n26180, n26179, 
        n26178, n26177, n24548;
    wire [4:0]n8404;
    
    wire n4_adj_4128, n26176, n26175, n26174, n24906, n26173;
    wire [0:0]n6842;
    wire [21:0]n8429;
    
    wire n26172, n26171, n25041, n26170, n26169, n26168, n25111, 
        n24905, n26167, n26166, n26165, n26164, n25040, n25110, 
        n26163, n26162, n26161, n26160, n26159, n9_adj_4132, n33437, 
        n25039, n26158, n26157, n62_adj_4133, n131_adj_4134, n26156, 
        n26155, n26154, n26153, n26152, n26151, n26150, n25109, 
        n26149, n25108, n24904, n25038, n25107, n25106, n24903, 
        n26148, n25037, n26147, n26146, n26145, n26144, n26143, 
        n26142, n26141, n26140, n26139, n26138, n26137, n26136, 
        n26135, n26134, n26133, n26132, n26131, n26130;
    wire [5:0]n8396;
    
    wire n26129, n417_adj_4136, n26128, n344_adj_4137, n26127, n271_adj_4138, 
        n26126, n198_adj_4139, n26125, n56_adj_4140, n125_adj_4141;
    wire [6:0]n8387;
    
    wire n560_adj_4142, n26124, n487_adj_4143, n26123, n414_adj_4144, 
        n26122, n341_adj_4145, n26121, n268_adj_4146, n26120, n195_adj_4147, 
        n26119, n53_adj_4148, n122_adj_4149, n25036;
    wire [7:0]n8377;
    
    wire n630_adj_4150, n26118, n557_adj_4151, n26117, n25105, n24902, 
        n484_adj_4154, n26116, n86_adj_4155, n17_adj_4156, n25104, 
        n159_adj_4158, n25035, n25034, n411_adj_4159, n26115, n338_adj_4160, 
        n26114, n25103, n25033, n265_adj_4162, n26113, n25102, n25101, 
        n192_adj_4165, n26112, n50_adj_4166, n119_adj_4167;
    wire [8:0]n8366;
    
    wire n700_adj_4168, n26111, n627_adj_4169, n26110, n25032, n554_adj_4170, 
        n26109, n481_adj_4171, n26108, n408_adj_4172, n26107, n335_adj_4173, 
        n26106, n262_adj_4174, n26105, n25100, n25031, n189_adj_4176, 
        n26104, n47_adj_4177, n116_adj_4178;
    wire [9:0]n8354;
    
    wire n770_adj_4179, n26103, n25099, n697_adj_4181, n26102, n624_adj_4182, 
        n26101, n551_adj_4183, n26100, n478_adj_4184, n26099, n405_adj_4185, 
        n26098, n332_adj_4186, n26097, n259_adj_4187, n26096, n33799, 
        n186_adj_4188, n26095, n25098, n25097, n44_adj_4191, n113_adj_4192;
    wire [10:0]n8341;
    
    wire n840_adj_4193, n26094, n767_adj_4194, n26093, n232_adj_4195, 
        n694_adj_4196, n26092, n17_adj_4197, n621_adj_4198, n26091, 
        n548_adj_4199, n26090, n475_adj_4200, n26089, n402_adj_4201, 
        n26088, n329_adj_4202, n26087, n305_adj_4203, n256_adj_4204, 
        n26086, n183_adj_4205, n26085, n41_adj_4206, n110_adj_4207;
    wire [11:0]n8327;
    
    wire n910_adj_4208, n26084, n837_adj_4209, n26083, n764_adj_4210, 
        n26082, n691_adj_4211, n26081, n618_adj_4212, n26080, n545_adj_4213, 
        n26079, n378_adj_4214, n472_adj_4215, n26078, n399_adj_4216, 
        n26077, n326_adj_4217, n26076, n253_adj_4218, n26075, n180_adj_4219, 
        n26074, n38_adj_4220, n107_adj_4221;
    wire [12:0]n8312;
    
    wire n980_adj_4222, n26073, n907_adj_4223, n26072, n834_adj_4224, 
        n26071, n761_adj_4225, n26070, n688_adj_4226, n26069, n615_adj_4227, 
        n26068, n542_adj_4228, n26067, n469_adj_4229, n26066, n396_adj_4230, 
        n26065, n323_adj_4231, n26064, n250_adj_4232, n26063, n177_adj_4233, 
        n26062, n25096, n35_adj_4235, n104_adj_4236;
    wire [13:0]n8296;
    
    wire n1050_adj_4237, n26061, n977_adj_4238, n26060, n904_adj_4239, 
        n26059, n831_adj_4240, n26058, n758_adj_4241, n26057, n25095, 
        n685_adj_4243, n26056, n612_adj_4244, n26055, n539_adj_4245, 
        n26054, n466_adj_4246, n26053, n393_adj_4247, n26052, n320_adj_4248, 
        n26051, n247_adj_4249, n26050, n174_adj_4250, n26049, n32_adj_4251, 
        n101_adj_4252, n451_adj_4253, n25094;
    wire [14:0]n8279;
    
    wire n1120_adj_4255, n26048, n1047_adj_4256, n26047, n974_adj_4257, 
        n26046, n24863, n524_adj_4258, n901_adj_4259, n26045, n25093, 
        n828_adj_4261, n26044, n755_adj_4262, n26043, n597_adj_4263, 
        n682_adj_4264, n26042, n24862, n670_adj_4265, n609_adj_4266, 
        n26041, n743_adj_4267, n816_adj_4268, n536_adj_4269, n26040, 
        n889_adj_4270, n463_adj_4271, n26039, n390_adj_4272, n26038, 
        n317_adj_4273, n26037, n244_adj_4274, n26036, n171_adj_4275, 
        n26035, n29_adj_4276, n98_adj_4277;
    wire [15:0]n8261;
    
    wire n26034, n1117_adj_4278, n26033, n1044_adj_4279, n26032, n971_adj_4280, 
        n26031, n898_adj_4281, n26030, n825_adj_4282, n26029, n752_adj_4283, 
        n26028, n679_adj_4284, n26027, n606_adj_4285, n26026, n533_adj_4286, 
        n26025, n460_adj_4287, n26024, n387_adj_4288, n26023, n314_adj_4289, 
        n26022, n241_adj_4290, n26021, n168_adj_4291, n26020, n25092, 
        n26_adj_4293, n95_adj_4294;
    wire [16:0]n8242;
    
    wire n26019, n26018, n24861, n1114_adj_4295, n26017, n25091, 
        n1041_adj_4297, n26016, n968_adj_4298, n26015, n895_adj_4299, 
        n26014, n822_adj_4300, n26013, n749_adj_4301, n26012, n676_adj_4302, 
        n26011, n25090, n603_adj_4304, n26010, n530_adj_4305, n26009, 
        n457_adj_4306, n26008, n384_adj_4307, n26007, n25089, n311_adj_4309, 
        n26006, n238_adj_4310, n26005, n165_adj_4311, n26004, n23_adj_4312, 
        n92_adj_4313;
    wire [17:0]n8222;
    
    wire n26003, n26002, n26001, n1111_adj_4314, n26000, n1038_adj_4315, 
        n25999, n965_adj_4316, n25998, n892_adj_4317, n25997, n819_adj_4318, 
        n25996, n746_adj_4319, n25995, n25088, n673_adj_4321, n25994, 
        n24860, n600_adj_4322, n25993, n527_adj_4323, n25992, n454_adj_4324, 
        n25991, n381_adj_4325, n25990, n308_adj_4326, n25989, n25087, 
        n235_adj_4329, n25988, n162_adj_4330, n25987, n20_adj_4331, 
        n89_adj_4332;
    wire [18:0]n8201;
    
    wire n25986, n25985, n25984, n25983, n1108_adj_4333, n25982, 
        n1035_adj_4334, n25981, n24859, n962_adj_4335, n25980, n25086, 
        n25979, n25978, n25977, n25976, n25975, n25974, n25973, 
        n25972, n25971, n25970, n25969;
    wire [19:0]n8179;
    
    wire n25968, n25085, n25967, n25966, n25965, n25964, n25963, 
        n25962, n25961, n25960, n25959, n25958, n25957, n25956, 
        n25955, n25954, n25953, n25952, n25951, n25950;
    wire [20:0]n8156;
    
    wire n25949, n25948, n25947, n25946, n25945, n25944, n25943, 
        n25942, n25941, n25940, n25084, n25939, n25938, n25937, 
        n25936, n25935, n25934, n25933, n25932, n25931, n25930;
    wire [0:0]n6838;
    wire [21:0]n8132;
    
    wire n25929, n25928, n25927, n25926, n25925, n25924, n25923, 
        n25922, n25921, n25920, n25919, n25918, n25083, n24858, 
        n25082, n24924, n25917, n24857, n25081, n25916, n25080, 
        n25915, n25914, n24923, n25079, n25913, n25078, n4_adj_4336, 
        n25912, n25911, n25910, n25909, n24680, n25908, n25077, 
        n25901, n25900, n25899, n25898, n25897, n25896, n25895, 
        n25894, n25893, n25892, n25891, n25890, n25889, n25888, 
        n25887, n25886, n25885, n25884, n25883, n25882, n25881, 
        n24757, n24922, n24921, n24920;
    
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_19 (.CI(n24918), .I0(n106[17]), .I1(n155[17]), .CO(n24919));
    SB_LUT4 i20563_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n8422[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20563_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_563_17 (.CI(n24855), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n2629[15]), .CO(n24856));
    SB_CARRY add_563_8 (.CI(n24846), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n2629[6]), .CO(n24847));
    SB_LUT4 i2_4_lut (.I0(n4_adj_3913), .I1(\Kp[3] ), .I2(n8417[1]), .I3(n1[19]), 
            .O(n8411[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1471 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1471.LUT_INIT = 16'h9c50;
    SB_LUT4 i20499_4_lut (.I0(n8411[2]), .I1(\Kp[4] ), .I2(n6_adj_3914), 
            .I3(n1[18]), .O(n8_adj_3915));   // verilog/motorControl.v(34[16:22])
    defparam i20499_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), .I3(n1[21]), 
            .O(n11));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i20530_4_lut (.I0(n8417[1]), .I1(\Kp[3] ), .I2(n4_adj_3913), 
            .I3(n1[19]), .O(n6_adj_3916));   // verilog/motorControl.v(34[16:22])
    defparam i20530_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20565_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n24650));   // verilog/motorControl.v(34[16:22])
    defparam i20565_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_3916), .I1(n11), .I2(n8_adj_3915), .I3(n12), 
            .O(n18));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), .I3(n1[22]), 
            .O(n13));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13), .I1(n18), .I2(n24650), .I3(n4_adj_3917), 
            .O(n30955));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3918));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17462_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17462_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17454_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17454_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17463_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17455_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17464_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_3921));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3922));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_3924));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_3925));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3927));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_3928));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_3929));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4693_7_lut (.I0(GND_net), .I1(n31043), .I2(n490_adj_3930), 
            .I3(n26372), .O(n8693[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4693_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4693_6_lut (.I0(GND_net), .I1(n8701[3]), .I2(n417), .I3(n26371), 
            .O(n8693[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4693_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4693_6 (.CI(n26371), .I0(n8701[3]), .I1(n417), .CO(n26372));
    SB_LUT4 add_4693_5_lut (.I0(GND_net), .I1(n8701[2]), .I2(n344), .I3(n26370), 
            .O(n8693[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4693_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4693_5 (.CI(n26370), .I0(n8701[2]), .I1(n344), .CO(n26371));
    SB_LUT4 add_4693_4_lut (.I0(GND_net), .I1(n8701[1]), .I2(n271), .I3(n26369), 
            .O(n8693[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4693_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4693_4 (.CI(n26369), .I0(n8701[1]), .I1(n271), .CO(n26370));
    SB_LUT4 add_4693_3_lut (.I0(GND_net), .I1(n8701[0]), .I2(n198), .I3(n26368), 
            .O(n8693[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4693_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4693_3 (.CI(n26368), .I0(n8701[0]), .I1(n198), .CO(n26369));
    SB_LUT4 add_4693_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n8693[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4693_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4693_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n26368));
    SB_LUT4 add_4692_8_lut (.I0(GND_net), .I1(n8693[5]), .I2(n560), .I3(n26367), 
            .O(n8684[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4692_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4692_7_lut (.I0(GND_net), .I1(n8693[4]), .I2(n487), .I3(n26366), 
            .O(n8684[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4692_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4692_7 (.CI(n26366), .I0(n8693[4]), .I1(n487), .CO(n26367));
    SB_LUT4 add_4692_6_lut (.I0(GND_net), .I1(n8693[3]), .I2(n414), .I3(n26365), 
            .O(n8684[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4692_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4692_6 (.CI(n26365), .I0(n8693[3]), .I1(n414), .CO(n26366));
    SB_LUT4 add_4692_5_lut (.I0(GND_net), .I1(n8693[2]), .I2(n341), .I3(n26364), 
            .O(n8684[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4692_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4692_5 (.CI(n26364), .I0(n8693[2]), .I1(n341), .CO(n26365));
    SB_LUT4 add_4692_4_lut (.I0(GND_net), .I1(n8693[1]), .I2(n268), .I3(n26363), 
            .O(n8684[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4692_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4692_4 (.CI(n26363), .I0(n8693[1]), .I1(n268), .CO(n26364));
    SB_LUT4 add_4692_3_lut (.I0(GND_net), .I1(n8693[0]), .I2(n195), .I3(n26362), 
            .O(n8684[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4692_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4692_3 (.CI(n26362), .I0(n8693[0]), .I1(n195), .CO(n26363));
    SB_LUT4 add_4692_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n8684[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4692_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4692_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n26362));
    SB_LUT4 add_4691_9_lut (.I0(GND_net), .I1(n8684[6]), .I2(n630), .I3(n26361), 
            .O(n8674[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4691_8_lut (.I0(GND_net), .I1(n8684[5]), .I2(n557), .I3(n26360), 
            .O(n8674[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4691_8 (.CI(n26360), .I0(n8684[5]), .I1(n557), .CO(n26361));
    SB_LUT4 add_4691_7_lut (.I0(GND_net), .I1(n8684[4]), .I2(n484), .I3(n26359), 
            .O(n8674[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4691_7 (.CI(n26359), .I0(n8684[4]), .I1(n484), .CO(n26360));
    SB_LUT4 add_4691_6_lut (.I0(GND_net), .I1(n8684[3]), .I2(n411), .I3(n26358), 
            .O(n8674[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4691_6 (.CI(n26358), .I0(n8684[3]), .I1(n411), .CO(n26359));
    SB_LUT4 add_4691_5_lut (.I0(GND_net), .I1(n8684[2]), .I2(n338), .I3(n26357), 
            .O(n8674[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4691_5 (.CI(n26357), .I0(n8684[2]), .I1(n338), .CO(n26358));
    SB_LUT4 add_4691_4_lut (.I0(GND_net), .I1(n8684[1]), .I2(n265), .I3(n26356), 
            .O(n8674[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4691_4 (.CI(n26356), .I0(n8684[1]), .I1(n265), .CO(n26357));
    SB_LUT4 add_4691_3_lut (.I0(GND_net), .I1(n8684[0]), .I2(n192), .I3(n26355), 
            .O(n8674[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4691_3 (.CI(n26355), .I0(n8684[0]), .I1(n192), .CO(n26356));
    SB_LUT4 add_4691_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n8674[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4691_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4691_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n26355));
    SB_LUT4 add_4690_10_lut (.I0(GND_net), .I1(n8674[7]), .I2(n700), .I3(n26354), 
            .O(n8663[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4690_9_lut (.I0(GND_net), .I1(n8674[6]), .I2(n627), .I3(n26353), 
            .O(n8663[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_9 (.CI(n26353), .I0(n8674[6]), .I1(n627), .CO(n26354));
    SB_LUT4 add_4690_8_lut (.I0(GND_net), .I1(n8674[5]), .I2(n554), .I3(n26352), 
            .O(n8663[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_8 (.CI(n26352), .I0(n8674[5]), .I1(n554), .CO(n26353));
    SB_LUT4 add_4690_7_lut (.I0(GND_net), .I1(n8674[4]), .I2(n481), .I3(n26351), 
            .O(n8663[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_7 (.CI(n26351), .I0(n8674[4]), .I1(n481), .CO(n26352));
    SB_LUT4 add_4690_6_lut (.I0(GND_net), .I1(n8674[3]), .I2(n408), .I3(n26350), 
            .O(n8663[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_6 (.CI(n26350), .I0(n8674[3]), .I1(n408), .CO(n26351));
    SB_LUT4 add_4690_5_lut (.I0(GND_net), .I1(n8674[2]), .I2(n335), .I3(n26349), 
            .O(n8663[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_5 (.CI(n26349), .I0(n8674[2]), .I1(n335), .CO(n26350));
    SB_LUT4 add_4690_4_lut (.I0(GND_net), .I1(n8674[1]), .I2(n262), .I3(n26348), 
            .O(n8663[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_4 (.CI(n26348), .I0(n8674[1]), .I1(n262), .CO(n26349));
    SB_LUT4 add_4690_3_lut (.I0(GND_net), .I1(n8674[0]), .I2(n189), .I3(n26347), 
            .O(n8663[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_3 (.CI(n26347), .I0(n8674[0]), .I1(n189), .CO(n26348));
    SB_LUT4 add_4690_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n8663[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n26347));
    SB_LUT4 add_4689_11_lut (.I0(GND_net), .I1(n8663[8]), .I2(n770), .I3(n26346), 
            .O(n8651[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4689_10_lut (.I0(GND_net), .I1(n8663[7]), .I2(n697), .I3(n26345), 
            .O(n8651[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17465_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4689_10 (.CI(n26345), .I0(n8663[7]), .I1(n697), .CO(n26346));
    SB_LUT4 add_4689_9_lut (.I0(GND_net), .I1(n8663[6]), .I2(n624), .I3(n26344), 
            .O(n8651[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4689_9 (.CI(n26344), .I0(n8663[6]), .I1(n624), .CO(n26345));
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_3932));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4689_8_lut (.I0(GND_net), .I1(n8663[5]), .I2(n551), .I3(n26343), 
            .O(n8651[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4689_8 (.CI(n26343), .I0(n8663[5]), .I1(n551), .CO(n26344));
    SB_LUT4 i27999_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n35222), 
            .I2(IntegralLimit[11]), .I3(n33677), .O(n33675));
    defparam i27999_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_4689_7_lut (.I0(GND_net), .I1(n8663[4]), .I2(n478), .I3(n26342), 
            .O(n8651[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4689_7 (.CI(n26342), .I0(n8663[4]), .I1(n478), .CO(n26343));
    SB_LUT4 add_4689_6_lut (.I0(GND_net), .I1(n8663[3]), .I2(n405), .I3(n26341), 
            .O(n8651[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4689_6 (.CI(n26341), .I0(n8663[3]), .I1(n405), .CO(n26342));
    SB_LUT4 add_4689_5_lut (.I0(GND_net), .I1(n8663[2]), .I2(n332), .I3(n26340), 
            .O(n8651[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4689_5 (.CI(n26340), .I0(n8663[2]), .I1(n332), .CO(n26341));
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3934));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n24917), .O(duty_23__N_3516[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4689_4_lut (.I0(GND_net), .I1(n8663[1]), .I2(n259), .I3(n26339), 
            .O(n8651[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3516[1]), .I1(n257[1]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3491[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_3935));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4689_4 (.CI(n26339), .I0(n8663[1]), .I1(n259), .CO(n26340));
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_3936));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4689_3_lut (.I0(GND_net), .I1(n8663[0]), .I2(n186_adj_3937), 
            .I3(n26338), .O(n8651[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4689_3 (.CI(n26338), .I0(n8663[0]), .I1(n186_adj_3937), 
            .CO(n26339));
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_3938));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_563_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n2629[5]), .I3(n24845), .O(\PID_CONTROLLER.integral_23__N_3416 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_7 (.CI(n24845), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n2629[5]), .CO(n24846));
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3939));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_3940));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_3941));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_43_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n35216));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_3942));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_3943));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_3944));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4689_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n8651[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4689_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_3945));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4689_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n26338));
    SB_LUT4 add_4688_12_lut (.I0(GND_net), .I1(n8651[9]), .I2(n840), .I3(n26337), 
            .O(n8638[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4688_11_lut (.I0(GND_net), .I1(n8651[8]), .I2(n767), .I3(n26336), 
            .O(n8638[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_11 (.CI(n26336), .I0(n8651[8]), .I1(n767), .CO(n26337));
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3946));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4688_10_lut (.I0(GND_net), .I1(n8651[7]), .I2(n694), .I3(n26335), 
            .O(n8638[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17466_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17466_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17456_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17456_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4688_10 (.CI(n26335), .I0(n8651[7]), .I1(n694), .CO(n26336));
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27683_4_lut (.I0(n27), .I1(n15_adj_3948), .I2(n13_adj_3949), 
            .I3(n11_adj_3950), .O(n33357));
    defparam i27683_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_831_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3516[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3516[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3516[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4688_9_lut (.I0(GND_net), .I1(n8651[6]), .I2(n621), .I3(n26334), 
            .O(n8638[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_9 (.CI(n26334), .I0(n8651[6]), .I1(n621), .CO(n26335));
    SB_LUT4 duty_23__I_831_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3516[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3516[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3516[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4688_8_lut (.I0(GND_net), .I1(n8651[5]), .I2(n548), .I3(n26333), 
            .O(n8638[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_8 (.CI(n26333), .I0(n8651[5]), .I1(n548), .CO(n26334));
    SB_LUT4 add_4688_7_lut (.I0(GND_net), .I1(n8651[4]), .I2(n475), .I3(n26332), 
            .O(n8638[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_7 (.CI(n26332), .I0(n8651[4]), .I1(n475), .CO(n26333));
    SB_LUT4 duty_23__I_831_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3516[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3951));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4688_6_lut (.I0(GND_net), .I1(n8651[3]), .I2(n402), .I3(n26331), 
            .O(n8638[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_6 (.CI(n26331), .I0(n8651[3]), .I1(n402), .CO(n26332));
    SB_LUT4 add_4688_5_lut (.I0(GND_net), .I1(n8651[2]), .I2(n329), .I3(n26330), 
            .O(n8638[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3516[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_3952));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4688_5 (.CI(n26330), .I0(n8651[2]), .I1(n329), .CO(n26331));
    SB_LUT4 add_4688_4_lut (.I0(GND_net), .I1(n8651[1]), .I2(n256_adj_3953), 
            .I3(n26329), .O(n8638[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_4 (.CI(n26329), .I0(n8651[1]), .I1(n256_adj_3953), 
            .CO(n26330));
    SB_LUT4 add_4688_3_lut (.I0(GND_net), .I1(n8651[0]), .I2(n183), .I3(n26328), 
            .O(n8638[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_3 (.CI(n26328), .I0(n8651[0]), .I1(n183), .CO(n26329));
    SB_LUT4 add_4688_2_lut (.I0(GND_net), .I1(n41_adj_3954), .I2(n110), 
            .I3(GND_net), .O(n8638[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4688_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4688_2 (.CI(GND_net), .I0(n41_adj_3954), .I1(n110), .CO(n26328));
    SB_LUT4 add_4687_13_lut (.I0(GND_net), .I1(n8638[10]), .I2(n910), 
            .I3(n26327), .O(n8624[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3516[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3955));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4687_12_lut (.I0(GND_net), .I1(n8638[9]), .I2(n837), .I3(n26326), 
            .O(n8624[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3516[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3956));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3516[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3957));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4687_12 (.CI(n26326), .I0(n8638[9]), .I1(n837), .CO(n26327));
    SB_LUT4 duty_23__I_831_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3516[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3958));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3516[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_3959));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4687_11_lut (.I0(GND_net), .I1(n8638[8]), .I2(n764), .I3(n26325), 
            .O(n8624[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4687_11 (.CI(n26325), .I0(n8638[8]), .I1(n764), .CO(n26326));
    SB_LUT4 duty_23__I_831_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3516[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4687_10_lut (.I0(GND_net), .I1(n8638[7]), .I2(n691), .I3(n26324), 
            .O(n8624[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3516[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3960));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4687_10 (.CI(n26324), .I0(n8638[7]), .I1(n691), .CO(n26325));
    SB_LUT4 duty_23__I_831_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3516[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3961));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4687_9_lut (.I0(GND_net), .I1(n8638[6]), .I2(n618), .I3(n26323), 
            .O(n8624[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3516[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3516[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4687_9 (.CI(n26323), .I0(n8638[6]), .I1(n618), .CO(n26324));
    SB_LUT4 add_4687_8_lut (.I0(GND_net), .I1(n8638[5]), .I2(n545), .I3(n26322), 
            .O(n8624[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27647_4_lut (.I0(n21), .I1(n19), .I2(n17_adj_3961), .I3(n9_adj_3960), 
            .O(n33321));
    defparam i27647_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4687_8 (.CI(n26322), .I0(n8638[5]), .I1(n545), .CO(n26323));
    SB_LUT4 i27641_4_lut (.I0(n27_adj_3959), .I1(n15_adj_3958), .I2(n13_adj_3957), 
            .I3(n11_adj_3956), .O(n33315));
    defparam i27641_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_831_i12_3_lut (.I0(duty_23__N_3516[7]), .I1(duty_23__N_3516[16]), 
            .I2(n33), .I3(GND_net), .O(n12_adj_3962));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4687_7_lut (.I0(GND_net), .I1(n8638[4]), .I2(n472), .I3(n26321), 
            .O(n8624[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4687_7 (.CI(n26321), .I0(n8638[4]), .I1(n472), .CO(n26322));
    SB_LUT4 add_4687_6_lut (.I0(GND_net), .I1(n8638[3]), .I2(n399), .I3(n26320), 
            .O(n8624[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i10_3_lut (.I0(duty_23__N_3516[5]), .I1(duty_23__N_3516[6]), 
            .I2(n13_adj_3957), .I3(GND_net), .O(n10));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4687_6 (.CI(n26320), .I0(n8638[3]), .I1(n399), .CO(n26321));
    SB_LUT4 duty_23__I_831_i30_3_lut (.I0(n12_adj_3962), .I1(duty_23__N_3516[17]), 
            .I2(n35_adj_3955), .I3(GND_net), .O(n30));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4687_5_lut (.I0(GND_net), .I1(n8638[2]), .I2(n326), .I3(n26319), 
            .O(n8624[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27927_4_lut (.I0(n13_adj_3957), .I1(n11_adj_3956), .I2(n9_adj_3960), 
            .I3(n33331), .O(n33603));
    defparam i27927_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i27923_4_lut (.I0(n19), .I1(n17_adj_3961), .I2(n15_adj_3958), 
            .I3(n33603), .O(n33599));
    defparam i27923_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i28233_4_lut (.I0(n25_adj_3952), .I1(n23_adj_3951), .I2(n21), 
            .I3(n33599), .O(n33909));
    defparam i28233_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_4687_5 (.CI(n26319), .I0(n8638[2]), .I1(n326), .CO(n26320));
    SB_LUT4 i28075_4_lut (.I0(n31), .I1(n29), .I2(n27_adj_3959), .I3(n33909), 
            .O(n33751));
    defparam i28075_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28286_4_lut (.I0(n37), .I1(n35_adj_3955), .I2(n33), .I3(n33751), 
            .O(n33962));
    defparam i28286_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_831_i16_3_lut (.I0(duty_23__N_3516[9]), .I1(duty_23__N_3516[21]), 
            .I2(n43), .I3(GND_net), .O(n16_adj_3964));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28219_3_lut (.I0(n6_adj_3965), .I1(duty_23__N_3516[10]), .I2(n21), 
            .I3(GND_net), .O(n33895));   // verilog/motorControl.v(36[10:25])
    defparam i28219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28220_3_lut (.I0(n33895), .I1(duty_23__N_3516[11]), .I2(n23_adj_3951), 
            .I3(GND_net), .O(n33896));   // verilog/motorControl.v(36[10:25])
    defparam i28220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i8_3_lut (.I0(duty_23__N_3516[4]), .I1(duty_23__N_3516[8]), 
            .I2(n17_adj_3961), .I3(GND_net), .O(n8_adj_3966));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i24_3_lut (.I0(n16_adj_3964), .I1(duty_23__N_3516[22]), 
            .I2(n45), .I3(GND_net), .O(n24_adj_3967));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27627_4_lut (.I0(n43), .I1(n25_adj_3952), .I2(n23_adj_3951), 
            .I3(n33321), .O(n33301));
    defparam i27627_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_12_18 (.CI(n24917), .I0(n106[16]), .I1(n155[16]), .CO(n24918));
    SB_LUT4 i28093_4_lut (.I0(n24_adj_3967), .I1(n8_adj_3966), .I2(n45), 
            .I3(n33299), .O(n33769));   // verilog/motorControl.v(36[10:25])
    defparam i28093_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_563_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n2629[14]), .I3(n24854), .O(\PID_CONTROLLER.integral_23__N_3416 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28160_3_lut (.I0(n33896), .I1(duty_23__N_3516[12]), .I2(n25_adj_3952), 
            .I3(GND_net), .O(n33836));   // verilog/motorControl.v(36[10:25])
    defparam i28160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i4_4_lut (.I0(duty_23__N_3516[0]), .I1(duty_23__N_3516[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_3968));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i28209_3_lut (.I0(n4_adj_3968), .I1(duty_23__N_3516[13]), .I2(n27_adj_3959), 
            .I3(GND_net), .O(n33885));   // verilog/motorControl.v(36[10:25])
    defparam i28209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28210_3_lut (.I0(n33885), .I1(\duty_23__N_3516[14] ), .I2(n29), 
            .I3(GND_net), .O(n33886));   // verilog/motorControl.v(36[10:25])
    defparam i28210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27637_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n33315), 
            .O(n33311));
    defparam i27637_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28296_4_lut (.I0(n30), .I1(n10), .I2(n35_adj_3955), .I3(n33309), 
            .O(n33972));   // verilog/motorControl.v(36[10:25])
    defparam i28296_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28162_3_lut (.I0(n33886), .I1(duty_23__N_3516[15]), .I2(n31), 
            .I3(GND_net), .O(n33838));   // verilog/motorControl.v(36[10:25])
    defparam i28162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28345_4_lut (.I0(n33838), .I1(n33972), .I2(n35_adj_3955), 
            .I3(n33311), .O(n34021));   // verilog/motorControl.v(36[10:25])
    defparam i28345_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28346_3_lut (.I0(n34021), .I1(duty_23__N_3516[18]), .I2(n37), 
            .I3(GND_net), .O(n34022));   // verilog/motorControl.v(36[10:25])
    defparam i28346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28327_3_lut (.I0(n34022), .I1(duty_23__N_3516[19]), .I2(n39), 
            .I3(GND_net), .O(n34003));   // verilog/motorControl.v(36[10:25])
    defparam i28327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27629_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n33962), 
            .O(n33303));
    defparam i27629_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28249_4_lut (.I0(n33836), .I1(n33769), .I2(n45), .I3(n33301), 
            .O(n33925));   // verilog/motorControl.v(36[10:25])
    defparam i28249_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28315_3_lut (.I0(n34003), .I1(duty_23__N_3516[20]), .I2(n41), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(36[10:25])
    defparam i28315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28251_4_lut (.I0(n40), .I1(n33925), .I2(n45), .I3(n33303), 
            .O(n33927));   // verilog/motorControl.v(36[10:25])
    defparam i28251_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28252_3_lut (.I0(n33927), .I1(PWMLimit[23]), .I2(duty_23__N_3516[23]), 
            .I3(GND_net), .O(duty_23__N_3515));   // verilog/motorControl.v(36[10:25])
    defparam i28252_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n24916), .O(duty_23__N_3516[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_563_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n2629[4]), .I3(n24844), .O(\PID_CONTROLLER.integral_23__N_3416 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3516[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_3971));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3516[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3972));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3516[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_3974));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3516[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_3975));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3516[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_3976));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(\duty_23__N_3516[14] ), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3977));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3516[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_3978));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3516[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3979));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3516[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_3980));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3516[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3981));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3516[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_3983));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4687_4_lut (.I0(GND_net), .I1(n8638[1]), .I2(n253), .I3(n26318), 
            .O(n8624[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3516[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3984));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3516[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3985));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3516[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3986));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3516[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_3988));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3516[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3989));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3516[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3990));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3516[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3991));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3516[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_3993));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i27611_4_lut (.I0(n21_adj_3993), .I1(n19_adj_3991), .I2(n17_adj_3990), 
            .I3(n9_adj_3989), .O(n33285));
    defparam i27611_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i27604_4_lut (.I0(n27_adj_3988), .I1(n15_adj_3986), .I2(n13_adj_3985), 
            .I3(n11_adj_3984), .O(n33278));
    defparam i27604_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_3983), 
            .I3(GND_net), .O(n12_adj_3994));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_3985), 
            .I3(GND_net), .O(n10_adj_3995));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_3994), .I1(n257[17]), .I2(n35_adj_3981), 
            .I3(GND_net), .O(n30_adj_3996));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27894_4_lut (.I0(n13_adj_3985), .I1(n11_adj_3984), .I2(n9_adj_3989), 
            .I3(n33296), .O(n33570));
    defparam i27894_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i27890_4_lut (.I0(n19_adj_3991), .I1(n17_adj_3990), .I2(n15_adj_3986), 
            .I3(n33570), .O(n33566));
    defparam i27890_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i28225_4_lut (.I0(n25_adj_3980), .I1(n23_adj_3979), .I2(n21_adj_3993), 
            .I3(n33566), .O(n33901));
    defparam i28225_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28059_4_lut (.I0(n31_adj_3978), .I1(n29_adj_3977), .I2(n27_adj_3988), 
            .I3(n33901), .O(n33735));
    defparam i28059_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28284_4_lut (.I0(n37_adj_3976), .I1(n35_adj_3981), .I2(n33_adj_3983), 
            .I3(n33735), .O(n33960));
    defparam i28284_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_3975), 
            .I3(GND_net), .O(n16_adj_3997));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28205_3_lut (.I0(n6_adj_3998), .I1(n257[10]), .I2(n21_adj_3993), 
            .I3(GND_net), .O(n33881));   // verilog/motorControl.v(38[19:35])
    defparam i28205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28206_3_lut (.I0(n33881), .I1(n257[11]), .I2(n23_adj_3979), 
            .I3(GND_net), .O(n33882));   // verilog/motorControl.v(38[19:35])
    defparam i28206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_3990), 
            .I3(GND_net), .O(n8_adj_3999));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_3997), .I1(n257[22]), .I2(n45_adj_3974), 
            .I3(GND_net), .O(n24_adj_4000));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27589_4_lut (.I0(n43_adj_3975), .I1(n25_adj_3980), .I2(n23_adj_3979), 
            .I3(n33285), .O(n33263));
    defparam i27589_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28095_4_lut (.I0(n24_adj_4000), .I1(n8_adj_3999), .I2(n45_adj_3974), 
            .I3(n33261), .O(n33771));   // verilog/motorControl.v(38[19:35])
    defparam i28095_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28166_3_lut (.I0(n33882), .I1(n257[12]), .I2(n25_adj_3980), 
            .I3(GND_net), .O(n33842));   // verilog/motorControl.v(38[19:35])
    defparam i28166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3516[0]), .I1(n257[1]), 
            .I2(duty_23__N_3516[1]), .I3(n257[0]), .O(n4_adj_4001));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i28203_3_lut (.I0(n4_adj_4001), .I1(n257[13]), .I2(n27_adj_3988), 
            .I3(GND_net), .O(n33879));   // verilog/motorControl.v(38[19:35])
    defparam i28203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28204_3_lut (.I0(n33879), .I1(n257[14]), .I2(n29_adj_3977), 
            .I3(GND_net), .O(n33880));   // verilog/motorControl.v(38[19:35])
    defparam i28204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27600_4_lut (.I0(n33_adj_3983), .I1(n31_adj_3978), .I2(n29_adj_3977), 
            .I3(n33278), .O(n33274));
    defparam i27600_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28298_4_lut (.I0(n30_adj_3996), .I1(n10_adj_3995), .I2(n35_adj_3981), 
            .I3(n33272), .O(n33974));   // verilog/motorControl.v(38[19:35])
    defparam i28298_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28168_3_lut (.I0(n33880), .I1(n257[15]), .I2(n31_adj_3978), 
            .I3(GND_net), .O(n33844));   // verilog/motorControl.v(38[19:35])
    defparam i28168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28347_4_lut (.I0(n33844), .I1(n33974), .I2(n35_adj_3981), 
            .I3(n33274), .O(n34023));   // verilog/motorControl.v(38[19:35])
    defparam i28347_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28348_3_lut (.I0(n34023), .I1(n257[18]), .I2(n37_adj_3976), 
            .I3(GND_net), .O(n34024));   // verilog/motorControl.v(38[19:35])
    defparam i28348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28325_3_lut (.I0(n34024), .I1(n257[19]), .I2(n39_adj_3971), 
            .I3(GND_net), .O(n34001));   // verilog/motorControl.v(38[19:35])
    defparam i28325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27591_4_lut (.I0(n43_adj_3975), .I1(n41_adj_3972), .I2(n39_adj_3971), 
            .I3(n33960), .O(n33265));
    defparam i27591_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28255_4_lut (.I0(n33842), .I1(n33771), .I2(n45_adj_3974), 
            .I3(n33263), .O(n33931));   // verilog/motorControl.v(38[19:35])
    defparam i28255_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28317_3_lut (.I0(n34001), .I1(n257[20]), .I2(n41_adj_3972), 
            .I3(GND_net), .O(n40_adj_4002));   // verilog/motorControl.v(38[19:35])
    defparam i28317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28257_4_lut (.I0(n40_adj_4002), .I1(n33931), .I2(n45_adj_3974), 
            .I3(n33265), .O(n33933));   // verilog/motorControl.v(38[19:35])
    defparam i28257_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28258_3_lut (.I0(n33933), .I1(duty_23__N_3516[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(38[19:35])
    defparam i28258_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3516[0]), .I1(n257[0]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3491[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17457_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17467_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3954));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4687_4 (.CI(n26318), .I0(n8638[1]), .I1(n253), .CO(n26319));
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17458_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17458_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3937));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4687_3_lut (.I0(GND_net), .I1(n8638[0]), .I2(n180), .I3(n26317), 
            .O(n8624[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4687_3 (.CI(n26317), .I0(n8638[0]), .I1(n180), .CO(n26318));
    SB_LUT4 add_4687_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n8624[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4687_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4687_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n26317));
    SB_CARRY add_12_17 (.CI(n24916), .I0(n106[15]), .I1(n155[15]), .CO(n24917));
    SB_LUT4 add_4686_14_lut (.I0(GND_net), .I1(n8624[11]), .I2(n980), 
            .I3(n26316), .O(n8609[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4686_13_lut (.I0(GND_net), .I1(n8624[10]), .I2(n907), 
            .I3(n26315), .O(n8609[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_13 (.CI(n26315), .I0(n8624[10]), .I1(n907), .CO(n26316));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3392[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_4686_12_lut (.I0(GND_net), .I1(n8624[9]), .I2(n834), .I3(n26314), 
            .O(n8609[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4686_12 (.CI(n26314), .I0(n8624[9]), .I1(n834), .CO(n26315));
    SB_LUT4 add_4686_11_lut (.I0(GND_net), .I1(n8624[8]), .I2(n761), .I3(n26313), 
            .O(n8609[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_11 (.CI(n26313), .I0(n8624[8]), .I1(n761), .CO(n26314));
    SB_LUT4 add_4686_10_lut (.I0(GND_net), .I1(n8624[7]), .I2(n688), .I3(n26312), 
            .O(n8609[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_10 (.CI(n26312), .I0(n8624[7]), .I1(n688), .CO(n26313));
    SB_LUT4 add_4686_9_lut (.I0(GND_net), .I1(n8624[6]), .I2(n615), .I3(n26311), 
            .O(n8609[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_9 (.CI(n26311), .I0(n8624[6]), .I1(n615), .CO(n26312));
    SB_LUT4 add_4686_8_lut (.I0(GND_net), .I1(n8624[5]), .I2(n542), .I3(n26310), 
            .O(n8609[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_16 (.CI(n24854), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n2629[14]), .CO(n24855));
    SB_CARRY add_4686_8 (.CI(n26310), .I0(n8624[5]), .I1(n542), .CO(n26311));
    SB_LUT4 add_4686_7_lut (.I0(GND_net), .I1(n8624[4]), .I2(n469), .I3(n26309), 
            .O(n8609[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_7 (.CI(n26309), .I0(n8624[4]), .I1(n469), .CO(n26310));
    SB_LUT4 add_4686_6_lut (.I0(GND_net), .I1(n8624[3]), .I2(n396), .I3(n26308), 
            .O(n8609[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_6 (.CI(n26308), .I0(n8624[3]), .I1(n396), .CO(n26309));
    SB_LUT4 add_4686_5_lut (.I0(GND_net), .I1(n8624[2]), .I2(n323), .I3(n26307), 
            .O(n8609[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27692_4_lut (.I0(n21_adj_4005), .I1(n19_adj_4006), .I2(n17_adj_4007), 
            .I3(n9_adj_4008), .O(n33366));
    defparam i27692_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4686_5 (.CI(n26307), .I0(n8624[2]), .I1(n323), .CO(n26308));
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4686_4_lut (.I0(GND_net), .I1(n8624[1]), .I2(n250), .I3(n26306), 
            .O(n8609[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_4 (.CI(n26306), .I0(n8624[1]), .I1(n250), .CO(n26307));
    SB_LUT4 add_4686_3_lut (.I0(GND_net), .I1(n8624[0]), .I2(n177), .I3(n26305), 
            .O(n8609[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_3 (.CI(n26305), .I0(n8624[0]), .I1(n177), .CO(n26306));
    SB_LUT4 add_4686_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n8609[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4686_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4686_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n26305));
    SB_LUT4 add_4685_15_lut (.I0(GND_net), .I1(n8609[12]), .I2(n1050), 
            .I3(n26304), .O(n8593[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4685_14_lut (.I0(GND_net), .I1(n8609[11]), .I2(n977), 
            .I3(n26303), .O(n8593[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_14 (.CI(n26303), .I0(n8609[11]), .I1(n977), .CO(n26304));
    SB_LUT4 add_4685_13_lut (.I0(GND_net), .I1(n8609[10]), .I2(n904), 
            .I3(n26302), .O(n8593[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_4009), .I3(GND_net), 
            .O(n16_adj_4010));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i27659_2_lut (.I0(n43_adj_4009), .I1(n19_adj_4006), .I2(GND_net), 
            .I3(GND_net), .O(n33333));
    defparam i27659_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_4685_13 (.CI(n26302), .I0(n8609[10]), .I1(n904), .CO(n26303));
    SB_LUT4 add_4685_12_lut (.I0(GND_net), .I1(n8609[9]), .I2(n831), .I3(n26301), 
            .O(n8593[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_12 (.CI(n26301), .I0(n8609[9]), .I1(n831), .CO(n26302));
    SB_LUT4 add_4685_11_lut (.I0(GND_net), .I1(n8609[8]), .I2(n758), .I3(n26300), 
            .O(n8593[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_11 (.CI(n26300), .I0(n8609[8]), .I1(n758), .CO(n26301));
    SB_LUT4 add_4685_10_lut (.I0(GND_net), .I1(n8609[7]), .I2(n685), .I3(n26299), 
            .O(n8593[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_10 (.CI(n26299), .I0(n8609[7]), .I1(n685), .CO(n26300));
    SB_CARRY add_563_6 (.CI(n24844), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n2629[4]), .CO(n24845));
    SB_LUT4 add_4685_9_lut (.I0(GND_net), .I1(n8609[6]), .I2(n612), .I3(n26298), 
            .O(n8593[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_9 (.CI(n26298), .I0(n8609[6]), .I1(n612), .CO(n26299));
    SB_LUT4 add_4685_8_lut (.I0(GND_net), .I1(n8609[5]), .I2(n539), .I3(n26297), 
            .O(n8593[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n2629[3]), .I3(n24843), .O(\PID_CONTROLLER.integral_23__N_3416 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_8 (.CI(n26297), .I0(n8609[5]), .I1(n539), .CO(n26298));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4007), .I3(GND_net), 
            .O(n8_adj_4011));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_4685_7_lut (.I0(GND_net), .I1(n8609[4]), .I2(n466), .I3(n26296), 
            .O(n8593[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_7 (.CI(n26296), .I0(n8609[4]), .I1(n466), .CO(n26297));
    SB_LUT4 add_4685_6_lut (.I0(GND_net), .I1(n8609[3]), .I2(n393), .I3(n26295), 
            .O(n8593[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n2629[13]), .I3(n24853), .O(\PID_CONTROLLER.integral_23__N_3416 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_6 (.CI(n26295), .I0(n8609[3]), .I1(n393), .CO(n26296));
    SB_LUT4 add_4685_5_lut (.I0(GND_net), .I1(n8609[2]), .I2(n320), .I3(n26294), 
            .O(n8593[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_5 (.CI(n26294), .I0(n8609[2]), .I1(n320), .CO(n26295));
    SB_LUT4 add_4685_4_lut (.I0(GND_net), .I1(n8609[1]), .I2(n247), .I3(n26293), 
            .O(n8593[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4014));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4015));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4016));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4017));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_563_5 (.CI(n24843), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n2629[3]), .CO(n24844));
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4018));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4019));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4020));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4022));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4024));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4025));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4027));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17470_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17470_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4028));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4685_4 (.CI(n26293), .I0(n8609[1]), .I1(n247), .CO(n26294));
    SB_LUT4 add_4685_3_lut (.I0(GND_net), .I1(n8609[0]), .I2(n174), .I3(n26292), 
            .O(n8593[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4685_3 (.CI(n26292), .I0(n8609[0]), .I1(n174), .CO(n26293));
    SB_LUT4 add_4685_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8593[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4685_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17471_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4685_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n26292));
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4031));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4684_16_lut (.I0(GND_net), .I1(n8593[13]), .I2(n1120), 
            .I3(n26291), .O(n8576[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4033));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4034));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4010), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_4035), .I3(GND_net), 
            .O(n24_adj_4036));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_4684_15_lut (.I0(GND_net), .I1(n8593[12]), .I2(n1047), 
            .I3(n26290), .O(n8576[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4684_15 (.CI(n26290), .I0(n8593[12]), .I1(n1047), .CO(n26291));
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4037));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4684_14_lut (.I0(GND_net), .I1(n8593[11]), .I2(n974), 
            .I3(n26289), .O(n8576[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4684_14 (.CI(n26289), .I0(n8593[11]), .I1(n974), .CO(n26290));
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4039));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4040));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4042));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4043));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4684_13_lut (.I0(GND_net), .I1(n8593[10]), .I2(n901), 
            .I3(n26288), .O(n8576[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4045));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4684_13 (.CI(n26288), .I0(n8593[10]), .I1(n901), .CO(n26289));
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n24915), .O(\duty_23__N_3516[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4048));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4049));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1472 (.I0(n6_adj_4050), .I1(\Ki[4] ), .I2(n8708[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [18]), .O(n8701[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1472.LUT_INIT = 16'h965a;
    SB_CARRY add_12_16 (.CI(n24915), .I0(n106[14]), .I1(n155[14]), .CO(n24916));
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_4051));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20685_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3416 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [21]), .O(n8719[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20685_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_4684_12_lut (.I0(GND_net), .I1(n8593[9]), .I2(n828), .I3(n26287), 
            .O(n8576[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4684_12 (.CI(n26287), .I0(n8593[9]), .I1(n828), .CO(n26288));
    SB_LUT4 i27724_2_lut (.I0(n7_adj_4052), .I1(n5_adj_4053), .I2(GND_net), 
            .I3(GND_net), .O(n33398));
    defparam i27724_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i27974_4_lut (.I0(n13_adj_3949), .I1(n11_adj_3950), .I2(n9_adj_4008), 
            .I3(n33398), .O(n33650));
    defparam i27974_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i27970_4_lut (.I0(n19_adj_4006), .I1(n17_adj_4007), .I2(n15_adj_3948), 
            .I3(n33650), .O(n33646));
    defparam i27970_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i28261_4_lut (.I0(n25_adj_4054), .I1(n23_adj_4055), .I2(n21_adj_4005), 
            .I3(n33646), .O(n33937));
    defparam i28261_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28101_4_lut (.I0(n31_adj_4056), .I1(n29_adj_4057), .I2(n27), 
            .I3(n33937), .O(n33777));
    defparam i28101_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28288_4_lut (.I0(n37_adj_4058), .I1(n35_adj_4059), .I2(n33_adj_4060), 
            .I3(n33777), .O(n33964));
    defparam i28288_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_66_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n35239));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_66_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28005_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n35239), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4061), .O(n33681));
    defparam i28005_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_36_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n35209));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_36_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i27993_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n35209), 
            .I2(IntegralLimit[14]), .I3(n33681), .O(n33669));
    defparam i27993_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_4684_11_lut (.I0(GND_net), .I1(n8593[8]), .I2(n755), .I3(n26286), 
            .O(n8576[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1473 (.I0(n4_adj_4062), .I1(\Ki[3] ), .I2(n8714[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [19]), .O(n8708[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1473.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_3930));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4684_11 (.CI(n26286), .I0(n8593[8]), .I1(n755), .CO(n26287));
    SB_LUT4 add_4684_10_lut (.I0(GND_net), .I1(n8593[7]), .I2(n682), .I3(n26285), 
            .O(n8576[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1474 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3416 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [20]), .O(n12_adj_4063));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1474.LUT_INIT = 16'h9c50;
    SB_CARRY add_4684_10 (.CI(n26285), .I0(n8593[7]), .I1(n682), .CO(n26286));
    SB_LUT4 i20621_4_lut (.I0(n8708[2]), .I1(\Ki[4] ), .I2(n6_adj_4050), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [18]), .O(n8_adj_4064));   // verilog/motorControl.v(34[25:36])
    defparam i20621_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_4684_9_lut (.I0(GND_net), .I1(n8593[6]), .I2(n609), .I3(n26284), 
            .O(n8576[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4684_9 (.CI(n26284), .I0(n8593[6]), .I1(n609), .CO(n26285));
    SB_LUT4 add_4684_8_lut (.I0(GND_net), .I1(n8593[5]), .I2(n536), .I3(n26283), 
            .O(n8576[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4684_8 (.CI(n26283), .I0(n8593[5]), .I1(n536), .CO(n26284));
    SB_LUT4 add_4684_7_lut (.I0(GND_net), .I1(n8593[4]), .I2(n463), .I3(n26282), 
            .O(n8576[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_15 (.CI(n24853), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n2629[13]), .CO(n24854));
    SB_CARRY add_4684_7 (.CI(n26282), .I0(n8593[4]), .I1(n463), .CO(n26283));
    SB_LUT4 add_4684_6_lut (.I0(GND_net), .I1(n8593[3]), .I2(n390), .I3(n26281), 
            .O(n8576[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4684_6 (.CI(n26281), .I0(n8593[3]), .I1(n390), .CO(n26282));
    SB_LUT4 i1_4_lut_adj_1475 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3416 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [21]), .O(n11_adj_4065));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut_adj_1475.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_4684_5_lut (.I0(GND_net), .I1(n8593[2]), .I2(n317), .I3(n26280), 
            .O(n8576[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4684_5 (.CI(n26280), .I0(n8593[2]), .I1(n317), .CO(n26281));
    SB_LUT4 add_4684_4_lut (.I0(GND_net), .I1(n8593[1]), .I2(n244), .I3(n26279), 
            .O(n8576[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4684_4 (.CI(n26279), .I0(n8593[1]), .I1(n244), .CO(n26280));
    SB_LUT4 add_4684_3_lut (.I0(GND_net), .I1(n8593[0]), .I2(n171), .I3(n26278), 
            .O(n8576[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4684_3 (.CI(n26278), .I0(n8593[0]), .I1(n171), .CO(n26279));
    SB_LUT4 add_4684_2_lut (.I0(GND_net), .I1(n29_c), .I2(n98), .I3(GND_net), 
            .O(n8576[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4684_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4684_2 (.CI(GND_net), .I0(n29_c), .I1(n98), .CO(n26278));
    SB_LUT4 i20652_4_lut (.I0(n8714[1]), .I1(\Ki[3] ), .I2(n4_adj_4062), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [19]), .O(n6_adj_4066));   // verilog/motorControl.v(34[25:36])
    defparam i20652_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_4683_17_lut (.I0(GND_net), .I1(n8576[14]), .I2(GND_net), 
            .I3(n26277), .O(n8558[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4683_16_lut (.I0(GND_net), .I1(n8576[13]), .I2(n1117), 
            .I3(n26276), .O(n8558[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_16 (.CI(n26276), .I0(n8576[13]), .I1(n1117), .CO(n26277));
    SB_LUT4 add_4683_15_lut (.I0(GND_net), .I1(n8576[12]), .I2(n1044), 
            .I3(n26275), .O(n8558[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n24914), .O(duty_23__N_3516[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20687_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3416 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [21]), .O(n24782));   // verilog/motorControl.v(34[25:36])
    defparam i20687_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_4683_15 (.CI(n26275), .I0(n8576[12]), .I1(n1044), .CO(n26276));
    SB_LUT4 add_4683_14_lut (.I0(GND_net), .I1(n8576[11]), .I2(n971), 
            .I3(n26274), .O(n8558[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n2629[12]), .I3(n24852), .O(\PID_CONTROLLER.integral_23__N_3416 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_15 (.CI(n24914), .I0(n106[13]), .I1(n155[13]), .CO(n24915));
    SB_LUT4 i8_4_lut_adj_1476 (.I0(n6_adj_4066), .I1(n11_adj_4065), .I2(n8_adj_4064), 
            .I3(n12_adj_4063), .O(n18_adj_4067));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1477 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3416 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3416 [22]), .O(n13_adj_4068));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut_adj_1477.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1478 (.I0(n13_adj_4068), .I1(n18_adj_4067), .I2(n24782), 
            .I3(n4_adj_4069), .O(n31043));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_CARRY add_4683_14 (.CI(n26274), .I0(n8576[11]), .I1(n971), .CO(n26275));
    SB_LUT4 add_4683_13_lut (.I0(GND_net), .I1(n8576[10]), .I2(n898), 
            .I3(n26273), .O(n8558[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_13 (.CI(n26273), .I0(n8576[10]), .I1(n898), .CO(n26274));
    SB_LUT4 add_4683_12_lut (.I0(GND_net), .I1(n8576[9]), .I2(n825), .I3(n26272), 
            .O(n8558[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_12 (.CI(n26272), .I0(n8576[9]), .I1(n825), .CO(n26273));
    SB_LUT4 add_4683_11_lut (.I0(GND_net), .I1(n8576[8]), .I2(n752), .I3(n26271), 
            .O(n8558[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_11 (.CI(n26271), .I0(n8576[8]), .I1(n752), .CO(n26272));
    SB_LUT4 add_4683_10_lut (.I0(GND_net), .I1(n8576[7]), .I2(n679), .I3(n26270), 
            .O(n8558[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_10 (.CI(n26270), .I0(n8576[7]), .I1(n679), .CO(n26271));
    SB_LUT4 add_4683_9_lut (.I0(GND_net), .I1(n8576[6]), .I2(n606), .I3(n26269), 
            .O(n8558[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_9 (.CI(n26269), .I0(n8576[6]), .I1(n606), .CO(n26270));
    SB_LUT4 add_4683_8_lut (.I0(GND_net), .I1(n8576[5]), .I2(n533), .I3(n26268), 
            .O(n8558[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_8 (.CI(n26268), .I0(n8576[5]), .I1(n533), .CO(n26269));
    SB_LUT4 add_4683_7_lut (.I0(GND_net), .I1(n8576[4]), .I2(n460), .I3(n26267), 
            .O(n8558[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_7 (.CI(n26267), .I0(n8576[4]), .I1(n460), .CO(n26268));
    SB_LUT4 add_4683_6_lut (.I0(GND_net), .I1(n8576[3]), .I2(n387), .I3(n26266), 
            .O(n8558[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_6 (.CI(n26266), .I0(n8576[3]), .I1(n387), .CO(n26267));
    SB_LUT4 add_4683_5_lut (.I0(GND_net), .I1(n8576[2]), .I2(n314), .I3(n26265), 
            .O(n8558[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_5 (.CI(n26265), .I0(n8576[2]), .I1(n314), .CO(n26266));
    SB_LUT4 add_4683_4_lut (.I0(GND_net), .I1(n8576[1]), .I2(n241), .I3(n26264), 
            .O(n8558[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n24913), .O(duty_23__N_3516[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_4 (.CI(n26264), .I0(n8576[1]), .I1(n241), .CO(n26265));
    SB_LUT4 add_4683_3_lut (.I0(GND_net), .I1(n8576[0]), .I2(n168), .I3(n26263), 
            .O(n8558[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_3 (.CI(n26263), .I0(n8576[0]), .I1(n168), .CO(n26264));
    SB_LUT4 add_4683_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n8558[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4683_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4683_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n26263));
    SB_LUT4 add_4682_18_lut (.I0(GND_net), .I1(n8558[15]), .I2(GND_net), 
            .I3(n26262), .O(n8539[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n25053), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_14 (.CI(n24852), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n2629[12]), .CO(n24853));
    SB_LUT4 add_4682_17_lut (.I0(GND_net), .I1(n8558[14]), .I2(GND_net), 
            .I3(n26261), .O(n8539[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n2629[11]), .I3(n24851), .O(\PID_CONTROLLER.integral_23__N_3416 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n2629[2]), .I3(n24842), .O(\PID_CONTROLLER.integral_23__N_3416 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n25052), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_4 (.CI(n24842), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n2629[2]), .CO(n24843));
    SB_CARRY add_563_13 (.CI(n24851), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n2629[11]), .CO(n24852));
    SB_LUT4 add_563_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n2629[10]), .I3(n24850), .O(\PID_CONTROLLER.integral_23__N_3416 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n25052), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n25053));
    SB_LUT4 add_563_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n2629[1]), .I3(n24841), .O(\PID_CONTROLLER.integral_23__N_3416 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n24913), .I0(n106[12]), .I1(n155[12]), .CO(n24914));
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4682_17 (.CI(n26261), .I0(n8558[14]), .I1(GND_net), .CO(n26262));
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n24912), .O(duty_23__N_3516[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_12 (.CI(n24850), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n2629[10]), .CO(n24851));
    SB_CARRY add_12_13 (.CI(n24912), .I0(n106[11]), .I1(n155[11]), .CO(n24913));
    SB_LUT4 add_4682_16_lut (.I0(GND_net), .I1(n8558[13]), .I2(n1114), 
            .I3(n26260), .O(n8539[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_16 (.CI(n26260), .I0(n8558[13]), .I1(n1114), .CO(n26261));
    SB_LUT4 add_4682_15_lut (.I0(GND_net), .I1(n8558[12]), .I2(n1041), 
            .I3(n26259), .O(n8539[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_15 (.CI(n26259), .I0(n8558[12]), .I1(n1041), .CO(n26260));
    SB_LUT4 add_4682_14_lut (.I0(GND_net), .I1(n8558[11]), .I2(n968), 
            .I3(n26258), .O(n8539[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_14 (.CI(n26258), .I0(n8558[11]), .I1(n968), .CO(n26259));
    SB_LUT4 add_4682_13_lut (.I0(GND_net), .I1(n8558[10]), .I2(n895), 
            .I3(n26257), .O(n8539[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_13 (.CI(n26257), .I0(n8558[10]), .I1(n895), .CO(n26258));
    SB_LUT4 add_4682_12_lut (.I0(GND_net), .I1(n8558[9]), .I2(n822), .I3(n26256), 
            .O(n8539[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_12 (.CI(n26256), .I0(n8558[9]), .I1(n822), .CO(n26257));
    SB_LUT4 add_4682_11_lut (.I0(GND_net), .I1(n8558[8]), .I2(n749), .I3(n26255), 
            .O(n8539[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_11 (.CI(n26255), .I0(n8558[8]), .I1(n749), .CO(n26256));
    SB_LUT4 add_4682_10_lut (.I0(GND_net), .I1(n8558[7]), .I2(n676), .I3(n26254), 
            .O(n8539[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_10 (.CI(n26254), .I0(n8558[7]), .I1(n676), .CO(n26255));
    SB_LUT4 add_563_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n2629[9]), .I3(n24849), .O(\PID_CONTROLLER.integral_23__N_3416 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4682_9_lut (.I0(GND_net), .I1(n8558[6]), .I2(n603), .I3(n26253), 
            .O(n8539[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_9 (.CI(n26253), .I0(n8558[6]), .I1(n603), .CO(n26254));
    SB_LUT4 add_4682_8_lut (.I0(GND_net), .I1(n8558[5]), .I2(n530), .I3(n26252), 
            .O(n8539[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_8 (.CI(n26252), .I0(n8558[5]), .I1(n530), .CO(n26253));
    SB_LUT4 add_4682_7_lut (.I0(GND_net), .I1(n8558[4]), .I2(n457), .I3(n26251), 
            .O(n8539[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n25051), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4072));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4073));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_31_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n35204));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4074));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4075));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27740_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n33414));
    defparam i27740_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_54_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n35227));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_54_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4076));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4074), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_4077));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28189_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n35222), 
            .I2(IntegralLimit[11]), .I3(n33679), .O(n33865));
    defparam i28189_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4078));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4682_7 (.CI(n26251), .I0(n8558[4]), .I1(n457), .CO(n26252));
    SB_LUT4 add_4682_6_lut (.I0(GND_net), .I1(n8558[3]), .I2(n384), .I3(n26250), 
            .O(n8539[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_6 (.CI(n26250), .I0(n8558[3]), .I1(n384), .CO(n26251));
    SB_LUT4 i27748_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n35216), 
            .I2(IntegralLimit[13]), .I3(n33865), .O(n33422));
    defparam i27748_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4079));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4682_5_lut (.I0(GND_net), .I1(n8558[2]), .I2(n311), .I3(n26249), 
            .O(n8539[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_5 (.CI(n26249), .I0(n8558[2]), .I1(n311), .CO(n26250));
    SB_CARRY add_563_9 (.CI(n24847), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n2629[7]), .CO(n24848));
    SB_LUT4 add_4682_4_lut (.I0(GND_net), .I1(n8558[1]), .I2(n238), .I3(n26248), 
            .O(n8539[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_4 (.CI(n26248), .I0(n8558[1]), .I1(n238), .CO(n26249));
    SB_LUT4 add_4682_3_lut (.I0(GND_net), .I1(n8558[0]), .I2(n165), .I3(n26247), 
            .O(n8539[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_3 (.CI(n26247), .I0(n8558[0]), .I1(n165), .CO(n26248));
    SB_LUT4 add_4682_2_lut (.I0(GND_net), .I1(n23_adj_4080), .I2(n92), 
            .I3(GND_net), .O(n8539[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_23 (.CI(n25051), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n25052));
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4081));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4082));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4083));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4084));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4085));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4086));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4087));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4089));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4090));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4091));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4093));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4094));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4095));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4097));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4682_2 (.CI(GND_net), .I0(n23_adj_4080), .I1(n92), .CO(n26247));
    SB_LUT4 add_4681_19_lut (.I0(GND_net), .I1(n8539[16]), .I2(GND_net), 
            .I3(n26246), .O(n8519[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n24911), .O(duty_23__N_3516[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n25050), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_22 (.CI(n25050), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n25051));
    SB_CARRY add_563_3 (.CI(n24841), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n2629[1]), .CO(n24842));
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n25049), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n25049), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n25050));
    SB_LUT4 add_4681_18_lut (.I0(GND_net), .I1(n8539[15]), .I2(GND_net), 
            .I3(n26245), .O(n8519[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_18 (.CI(n26245), .I0(n8539[15]), .I1(GND_net), .CO(n26246));
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n25048), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4681_17_lut (.I0(GND_net), .I1(n8539[14]), .I2(GND_net), 
            .I3(n26244), .O(n8519[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_34_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n35207));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_34_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_563_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n2629[8]), .I3(n24848), .O(\PID_CONTROLLER.integral_23__N_3416 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n2629[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3416 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_17 (.CI(n26244), .I0(n8539[14]), .I1(GND_net), .CO(n26245));
    SB_CARRY add_12_12 (.CI(n24911), .I0(n106[10]), .I1(n155[10]), .CO(n24912));
    SB_CARRY sub_3_add_2_20 (.CI(n25048), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n25049));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n24910), 
            .O(duty_23__N_3516[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28827_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34501));   // verilog/motorControl.v(29[14] 48[8])
    defparam i28827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_11 (.CI(n24910), .I0(n106[9]), .I1(n155[9]), .CO(n24911));
    SB_CARRY add_563_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n2629[0]), .CO(n24841));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n24909), 
            .O(duty_23__N_3516[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28117_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n35207), 
            .I2(IntegralLimit[15]), .I3(n33422), .O(n33793));
    defparam i28117_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_4681_16_lut (.I0(GND_net), .I1(n8539[13]), .I2(n1111), 
            .I3(n26243), .O(n8519[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_60_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n35233));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_60_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_10 (.CI(n24909), .I0(n106[8]), .I1(n155[8]), .CO(n24910));
    SB_CARRY add_563_10 (.CI(n24848), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n2629[8]), .CO(n24849));
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4681_16 (.CI(n26243), .I0(n8539[13]), .I1(n1111), .CO(n26244));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n25047), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_19 (.CI(n25047), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n25048));
    SB_LUT4 add_4681_15_lut (.I0(GND_net), .I1(n8539[12]), .I2(n1038), 
            .I3(n26242), .O(n8519[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_15 (.CI(n26242), .I0(n8539[12]), .I1(n1038), .CO(n26243));
    SB_LUT4 add_4681_14_lut (.I0(GND_net), .I1(n8539[11]), .I2(n965), 
            .I3(n26241), .O(n8519[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_14 (.CI(n26241), .I0(n8539[11]), .I1(n965), .CO(n26242));
    SB_LUT4 add_4681_13_lut (.I0(GND_net), .I1(n8539[10]), .I2(n892), 
            .I3(n26240), .O(n8519[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_13 (.CI(n26240), .I0(n8539[10]), .I1(n892), .CO(n26241));
    SB_LUT4 add_4681_12_lut (.I0(GND_net), .I1(n8539[9]), .I2(n819), .I3(n26239), 
            .O(n8519[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_12 (.CI(n26239), .I0(n8539[9]), .I1(n819), .CO(n26240));
    SB_LUT4 add_4681_11_lut (.I0(GND_net), .I1(n8539[8]), .I2(n746), .I3(n26238), 
            .O(n8519[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_11 (.CI(n26238), .I0(n8539[8]), .I1(n746), .CO(n26239));
    SB_LUT4 add_4681_10_lut (.I0(GND_net), .I1(n8539[7]), .I2(n673), .I3(n26237), 
            .O(n8519[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_10 (.CI(n26237), .I0(n8539[7]), .I1(n673), .CO(n26238));
    SB_LUT4 add_4681_9_lut (.I0(GND_net), .I1(n8539[6]), .I2(n600), .I3(n26236), 
            .O(n8519[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n24908), 
            .O(duty_23__N_3516[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28266_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n35233), 
            .I2(IntegralLimit[17]), .I3(n33793), .O(n33942));
    defparam i28266_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_4681_9 (.CI(n26236), .I0(n8539[6]), .I1(n600), .CO(n26237));
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4681_8_lut (.I0(GND_net), .I1(n8539[5]), .I2(n527), .I3(n26235), 
            .O(n8519[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_8 (.CI(n26235), .I0(n8539[5]), .I1(n527), .CO(n26236));
    SB_LUT4 add_4681_7_lut (.I0(GND_net), .I1(n8539[4]), .I2(n454), .I3(n26234), 
            .O(n8519[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_7 (.CI(n26234), .I0(n8539[4]), .I1(n454), .CO(n26235));
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[23]), 
            .I3(n25122), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[22]), 
            .I3(n25121), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n25121), .I0(GND_net), .I1(n1_adj_4337[22]), 
            .CO(n25122));
    SB_LUT4 add_4681_6_lut (.I0(GND_net), .I1(n8539[3]), .I2(n381), .I3(n26233), 
            .O(n8519[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[21]), 
            .I3(n25120), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_6 (.CI(n26233), .I0(n8539[3]), .I1(n381), .CO(n26234));
    SB_LUT4 add_4681_5_lut (.I0(GND_net), .I1(n8539[2]), .I2(n308), .I3(n26232), 
            .O(n8519[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_5 (.CI(n26232), .I0(n8539[2]), .I1(n308), .CO(n26233));
    SB_LUT4 add_4681_4_lut (.I0(GND_net), .I1(n8539[1]), .I2(n235), .I3(n26231), 
            .O(n8519[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_4 (.CI(n26231), .I0(n8539[1]), .I1(n235), .CO(n26232));
    SB_LUT4 add_4681_3_lut (.I0(GND_net), .I1(n8539[0]), .I2(n162), .I3(n26230), 
            .O(n8519[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_3 (.CI(n26230), .I0(n8539[0]), .I1(n162), .CO(n26231));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n25046), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4681_2_lut (.I0(GND_net), .I1(n20_adj_4104), .I2(n89), 
            .I3(GND_net), .O(n8519[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4681_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4681_2 (.CI(GND_net), .I0(n20_adj_4104), .I1(n89), .CO(n26230));
    SB_LUT4 add_4680_20_lut (.I0(GND_net), .I1(n8519[17]), .I2(GND_net), 
            .I3(n26229), .O(n8498[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4680_19_lut (.I0(GND_net), .I1(n8519[16]), .I2(GND_net), 
            .I3(n26228), .O(n8498[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_19 (.CI(n26228), .I0(n8519[16]), .I1(GND_net), .CO(n26229));
    SB_LUT4 add_4680_18_lut (.I0(GND_net), .I1(n8519[15]), .I2(GND_net), 
            .I3(n26227), .O(n8498[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_18 (.CI(n26227), .I0(n8519[15]), .I1(GND_net), .CO(n26228));
    SB_LUT4 add_4680_17_lut (.I0(GND_net), .I1(n8519[14]), .I2(GND_net), 
            .I3(n26226), .O(n8498[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_17 (.CI(n26226), .I0(n8519[14]), .I1(GND_net), .CO(n26227));
    SB_LUT4 add_4680_16_lut (.I0(GND_net), .I1(n8519[13]), .I2(n1108), 
            .I3(n26225), .O(n8498[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_16 (.CI(n26225), .I0(n8519[13]), .I1(n1108), .CO(n26226));
    SB_LUT4 add_4680_15_lut (.I0(GND_net), .I1(n8519[12]), .I2(n1035), 
            .I3(n26224), .O(n8498[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_15 (.CI(n26224), .I0(n8519[12]), .I1(n1035), .CO(n26225));
    SB_LUT4 add_4680_14_lut (.I0(GND_net), .I1(n8519[11]), .I2(n962), 
            .I3(n26223), .O(n8498[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n25120), .I0(GND_net), .I1(n1_adj_4337[21]), 
            .CO(n25121));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[20]), 
            .I3(n25119), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n25119), .I0(GND_net), .I1(n1_adj_4337[20]), 
            .CO(n25120));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[19]), 
            .I3(n25118), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n25118), .I0(GND_net), .I1(n1_adj_4337[19]), 
            .CO(n25119));
    SB_CARRY sub_3_add_2_18 (.CI(n25046), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n25047));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[18]), 
            .I3(n25117), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n25117), .I0(GND_net), .I1(n1_adj_4337[18]), 
            .CO(n25118));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[17]), 
            .I3(n25116), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n25045), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_9 (.CI(n24908), .I0(n106[7]), .I1(n155[7]), .CO(n24909));
    SB_CARRY unary_minus_16_add_3_19 (.CI(n25116), .I0(GND_net), .I1(n1_adj_4337[17]), 
            .CO(n25117));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[16]), 
            .I3(n25115), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_25_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n35198));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28320_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n35198), 
            .I2(IntegralLimit[19]), .I3(n33942), .O(n33996));
    defparam i28320_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_22_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n35195));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_22_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4111));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i27726_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n33400));
    defparam i27726_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4111), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4112));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4113));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28137_3_lut (.I0(n6_adj_4113), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n33813));   // verilog/motorControl.v(31[10:34])
    defparam i28137_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28138_3_lut (.I0(n33813), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n33814));   // verilog/motorControl.v(31[10:34])
    defparam i28138_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i27728_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n35216), 
            .I2(IntegralLimit[21]), .I3(n33675), .O(n33402));
    defparam i27728_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i28089_4_lut (.I0(n24_adj_4112), .I1(n8_adj_4114), .I2(n35193), 
            .I3(n33400), .O(n33765));   // verilog/motorControl.v(31[10:34])
    defparam i28089_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i27944_3_lut (.I0(n33814), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n33620));   // verilog/motorControl.v(31[10:34])
    defparam i27944_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3467 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4115), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4116));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i28129_3_lut (.I0(n4_adj_4116), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n33805));   // verilog/motorControl.v(31[38:63])
    defparam i28129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28130_3_lut (.I0(n33805), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4057), .I3(GND_net), .O(n33806));   // verilog/motorControl.v(31[38:63])
    defparam i28130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33_adj_4060), .I3(GND_net), 
            .O(n12_adj_4117));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i27671_2_lut (.I0(n33_adj_4060), .I1(n15_adj_3948), .I2(GND_net), 
            .I3(GND_net), .O(n33345));
    defparam i27671_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_3949), .I3(GND_net), 
            .O(n10_adj_4118));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4117), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4059), .I3(GND_net), 
            .O(n30_adj_4119));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_4680_14 (.CI(n26223), .I0(n8519[11]), .I1(n962), .CO(n26224));
    SB_LUT4 add_4680_13_lut (.I0(GND_net), .I1(n8519[10]), .I2(n889), 
            .I3(n26222), .O(n8498[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_13 (.CI(n26222), .I0(n8519[10]), .I1(n889), .CO(n26223));
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n25115), .I0(GND_net), .I1(n1_adj_4337[16]), 
            .CO(n25116));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[15]), 
            .I3(n25114), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4680_12_lut (.I0(GND_net), .I1(n8519[9]), .I2(n816), .I3(n26221), 
            .O(n8498[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_12 (.CI(n26221), .I0(n8519[9]), .I1(n816), .CO(n26222));
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4680_11_lut (.I0(GND_net), .I1(n8519[8]), .I2(n743), .I3(n26220), 
            .O(n8498[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n25114), .I0(GND_net), .I1(n1_adj_4337[15]), 
            .CO(n25115));
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4680_11 (.CI(n26220), .I0(n8519[8]), .I1(n743), .CO(n26221));
    SB_LUT4 add_4680_10_lut (.I0(GND_net), .I1(n8519[7]), .I2(n670), .I3(n26219), 
            .O(n8498[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_10 (.CI(n26219), .I0(n8519[7]), .I1(n670), .CO(n26220));
    SB_CARRY sub_3_add_2_17 (.CI(n25045), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n25046));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[14]), 
            .I3(n25113), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4680_9_lut (.I0(GND_net), .I1(n8519[6]), .I2(n597), .I3(n26218), 
            .O(n8498[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17459_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4680_9 (.CI(n26218), .I0(n8519[6]), .I1(n597), .CO(n26219));
    SB_LUT4 add_4680_8_lut (.I0(GND_net), .I1(n8519[5]), .I2(n524), .I3(n26217), 
            .O(n8498[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_8 (.CI(n26217), .I0(n8519[5]), .I1(n524), .CO(n26218));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n25113), .I0(GND_net), .I1(n1_adj_4337[14]), 
            .CO(n25114));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[13]), 
            .I3(n25112), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n24907), 
            .O(duty_23__N_3516[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4680_7_lut (.I0(GND_net), .I1(n8519[4]), .I2(n451), .I3(n26216), 
            .O(n8498[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_7 (.CI(n26216), .I0(n8519[4]), .I1(n451), .CO(n26217));
    SB_LUT4 add_4680_6_lut (.I0(GND_net), .I1(n8519[3]), .I2(n378), .I3(n26215), 
            .O(n8498[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_6 (.CI(n26215), .I0(n8519[3]), .I1(n378), .CO(n26216));
    SB_LUT4 add_4680_5_lut (.I0(GND_net), .I1(n8519[2]), .I2(n305), .I3(n26214), 
            .O(n8498[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_5 (.CI(n26214), .I0(n8519[2]), .I1(n305), .CO(n26215));
    SB_LUT4 add_4680_4_lut (.I0(GND_net), .I1(n8519[1]), .I2(n232), .I3(n26213), 
            .O(n8498[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_4 (.CI(n26213), .I0(n8519[1]), .I1(n232), .CO(n26214));
    SB_LUT4 add_4680_3_lut (.I0(GND_net), .I1(n8519[0]), .I2(n159), .I3(n26212), 
            .O(n8498[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n8422[0]), 
            .I3(n24625), .O(n8417[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i27677_4_lut (.I0(n33_adj_4060), .I1(n31_adj_4056), .I2(n29_adj_4057), 
            .I3(n33357), .O(n33351));
    defparam i27677_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28294_4_lut (.I0(n30_adj_4119), .I1(n10_adj_4118), .I2(n35_adj_4059), 
            .I3(n33345), .O(n33970));   // verilog/motorControl.v(31[38:63])
    defparam i28294_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i27957_3_lut (.I0(n33806), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_4056), .I3(GND_net), .O(n33633));   // verilog/motorControl.v(31[38:63])
    defparam i27957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28343_4_lut (.I0(n33633), .I1(n33970), .I2(n35_adj_4059), 
            .I3(n33351), .O(n34019));   // verilog/motorControl.v(31[38:63])
    defparam i28343_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28344_3_lut (.I0(n34019), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37_adj_4058), .I3(GND_net), .O(n34020));   // verilog/motorControl.v(31[38:63])
    defparam i28344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28329_3_lut (.I0(n34020), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_4121), .I3(GND_net), .O(n34005));   // verilog/motorControl.v(31[38:63])
    defparam i28329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4052), .I3(GND_net), 
            .O(n6_adj_4122));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i28155_3_lut (.I0(n6_adj_4122), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4005), .I3(GND_net), .O(n33831));   // verilog/motorControl.v(31[38:63])
    defparam i28155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28156_3_lut (.I0(n33831), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4055), .I3(GND_net), .O(n33832));   // verilog/motorControl.v(31[38:63])
    defparam i28156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27661_4_lut (.I0(n43_adj_4009), .I1(n25_adj_4054), .I2(n23_adj_4055), 
            .I3(n33366), .O(n33335));
    defparam i27661_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28091_4_lut (.I0(n24_adj_4036), .I1(n8_adj_4011), .I2(n45_adj_4035), 
            .I3(n33333), .O(n33767));   // verilog/motorControl.v(31[38:63])
    defparam i28091_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4680_3 (.CI(n26212), .I0(n8519[0]), .I1(n159), .CO(n26213));
    SB_LUT4 add_4680_2_lut (.I0(GND_net), .I1(n17_adj_3946), .I2(n86), 
            .I3(GND_net), .O(n8498[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4680_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4680_2 (.CI(GND_net), .I0(n17_adj_3946), .I1(n86), .CO(n26212));
    SB_LUT4 add_4679_21_lut (.I0(GND_net), .I1(n8498[18]), .I2(GND_net), 
            .I3(n26211), .O(n8476[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4679_20_lut (.I0(GND_net), .I1(n8498[17]), .I2(GND_net), 
            .I3(n26210), .O(n8476[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_20 (.CI(n26210), .I0(n8498[17]), .I1(GND_net), .CO(n26211));
    SB_LUT4 add_4679_19_lut (.I0(GND_net), .I1(n8498[16]), .I2(GND_net), 
            .I3(n26209), .O(n8476[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_19 (.CI(n26209), .I0(n8498[16]), .I1(GND_net), .CO(n26210));
    SB_LUT4 add_4679_18_lut (.I0(GND_net), .I1(n8498[15]), .I2(GND_net), 
            .I3(n26208), .O(n8476[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_18 (.CI(n26208), .I0(n8498[15]), .I1(GND_net), .CO(n26209));
    SB_LUT4 add_4679_17_lut (.I0(GND_net), .I1(n8498[14]), .I2(GND_net), 
            .I3(n26207), .O(n8476[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_17 (.CI(n26207), .I0(n8498[14]), .I1(GND_net), .CO(n26208));
    SB_LUT4 i17075_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17075_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17461_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n25044), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4679_16_lut (.I0(GND_net), .I1(n8498[13]), .I2(n1105), 
            .I3(n26206), .O(n8476[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27766_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n33440));
    defparam i27766_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n25112), .I0(GND_net), .I1(n1_adj_4337[13]), 
            .CO(n25113));
    SB_CARRY add_12_8 (.CI(n24907), .I0(n106[6]), .I1(n155[6]), .CO(n24908));
    SB_LUT4 i27955_3_lut (.I0(n33832), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4054), .I3(GND_net), .O(n33631));   // verilog/motorControl.v(31[38:63])
    defparam i27955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27663_4_lut (.I0(n43_adj_4009), .I1(n41_adj_4124), .I2(n39_adj_4121), 
            .I3(n33964), .O(n33337));
    defparam i27663_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28243_4_lut (.I0(n33631), .I1(n33767), .I2(n45_adj_4035), 
            .I3(n33335), .O(n33919));   // verilog/motorControl.v(31[38:63])
    defparam i28243_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4679_16 (.CI(n26206), .I0(n8498[13]), .I1(n1105), .CO(n26207));
    SB_CARRY sub_3_add_2_16 (.CI(n25044), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n25045));
    SB_LUT4 add_4679_15_lut (.I0(GND_net), .I1(n8498[12]), .I2(n1032), 
            .I3(n26205), .O(n8476[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_15 (.CI(n26205), .I0(n8498[12]), .I1(n1032), .CO(n26206));
    SB_LUT4 add_4679_14_lut (.I0(GND_net), .I1(n8498[11]), .I2(n959), 
            .I3(n26204), .O(n8476[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28313_3_lut (.I0(n34005), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4124), .I3(GND_net), .O(n40_adj_4125));   // verilog/motorControl.v(31[38:63])
    defparam i28313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28245_4_lut (.I0(n40_adj_4125), .I1(n33919), .I2(n45_adj_4035), 
            .I3(n33337), .O(n33921));   // verilog/motorControl.v(31[38:63])
    defparam i28245_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4126));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_4679_14 (.CI(n26204), .I0(n8498[11]), .I1(n959), .CO(n26205));
    SB_LUT4 i28135_3_lut (.I0(n4_adj_4126), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n33811));   // verilog/motorControl.v(31[10:34])
    defparam i28135_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4679_13_lut (.I0(GND_net), .I1(n8498[10]), .I2(n886), 
            .I3(n26203), .O(n8476[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_13 (.CI(n26203), .I0(n8498[10]), .I1(n886), .CO(n26204));
    SB_LUT4 i28136_3_lut (.I0(n33811), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n33812));   // verilog/motorControl.v(31[10:34])
    defparam i28136_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i27742_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n35204), 
            .I2(IntegralLimit[16]), .I3(n33669), .O(n33416));
    defparam i27742_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i28278_4_lut (.I0(n30_adj_4077), .I1(n10_adj_4076), .I2(n35227), 
            .I3(n33414), .O(n33954));   // verilog/motorControl.v(31[10:34])
    defparam i28278_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i27946_3_lut (.I0(n33812), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n33622));   // verilog/motorControl.v(31[10:34])
    defparam i27946_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28330_4_lut (.I0(n33622), .I1(n33954), .I2(n35227), .I3(n33416), 
            .O(n34006));   // verilog/motorControl.v(31[10:34])
    defparam i28330_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4679_12_lut (.I0(GND_net), .I1(n8498[9]), .I2(n813), .I3(n26202), 
            .O(n8476[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28331_3_lut (.I0(n34006), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n34007));   // verilog/motorControl.v(31[10:34])
    defparam i28331_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28305_3_lut (.I0(n34007), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n33981));   // verilog/motorControl.v(31[10:34])
    defparam i28305_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i27733_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n35195), 
            .I2(IntegralLimit[21]), .I3(n33996), .O(n33407));
    defparam i27733_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_20_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n35193));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28239_4_lut (.I0(n33620), .I1(n33765), .I2(n35193), .I3(n33402), 
            .O(n33915));   // verilog/motorControl.v(31[10:34])
    defparam i28239_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i27952_3_lut (.I0(n33981), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n33628));   // verilog/motorControl.v(31[10:34])
    defparam i27952_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28246_3_lut (.I0(n33921), .I1(\PID_CONTROLLER.integral_23__N_3467 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3466 ));   // verilog/motorControl.v(31[38:63])
    defparam i28246_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28290_4_lut (.I0(n33628), .I1(n33915), .I2(n35193), .I3(n33407), 
            .O(n33966));   // verilog/motorControl.v(31[10:34])
    defparam i28290_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_830_4_lut  (.I0(n33966), .I1(\PID_CONTROLLER.integral_23__N_3466 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3464 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_830_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n25043), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n25043), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n25044));
    SB_CARRY add_4679_12 (.CI(n26202), .I0(n8498[9]), .I1(n813), .CO(n26203));
    SB_LUT4 add_4679_11_lut (.I0(GND_net), .I1(n8498[8]), .I2(n740), .I3(n26201), 
            .O(n8476[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n25042), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_11 (.CI(n26201), .I0(n8498[8]), .I1(n740), .CO(n26202));
    SB_LUT4 add_4679_10_lut (.I0(GND_net), .I1(n8498[7]), .I2(n667), .I3(n26200), 
            .O(n8476[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_10 (.CI(n26200), .I0(n8498[7]), .I1(n667), .CO(n26201));
    SB_LUT4 add_4679_9_lut (.I0(GND_net), .I1(n8498[6]), .I2(n594), .I3(n26199), 
            .O(n8476[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_9 (.CI(n26199), .I0(n8498[6]), .I1(n594), .CO(n26200));
    SB_LUT4 add_4679_8_lut (.I0(GND_net), .I1(n8498[5]), .I2(n521), .I3(n26198), 
            .O(n8476[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_8 (.CI(n26198), .I0(n8498[5]), .I1(n521), .CO(n26199));
    SB_LUT4 i17468_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4679_7_lut (.I0(GND_net), .I1(n8498[4]), .I2(n448), .I3(n26197), 
            .O(n8476[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_7 (.CI(n26197), .I0(n8498[4]), .I1(n448), .CO(n26198));
    SB_LUT4 add_4679_6_lut (.I0(GND_net), .I1(n8498[3]), .I2(n375), .I3(n26196), 
            .O(n8476[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_6 (.CI(n26196), .I0(n8498[3]), .I1(n375), .CO(n26197));
    SB_LUT4 add_4679_5_lut (.I0(GND_net), .I1(n8498[2]), .I2(n302), .I3(n26195), 
            .O(n8476[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_5 (.CI(n26195), .I0(n8498[2]), .I1(n302), .CO(n26196));
    SB_LUT4 add_4679_4_lut (.I0(GND_net), .I1(n8498[1]), .I2(n229), .I3(n26194), 
            .O(n8476[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_4 (.CI(n26194), .I0(n8498[1]), .I1(n229), .CO(n26195));
    SB_LUT4 add_4679_3_lut (.I0(GND_net), .I1(n8498[0]), .I2(n156), .I3(n26193), 
            .O(n8476[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_3 (.CI(n26193), .I0(n8498[0]), .I1(n156), .CO(n26194));
    SB_LUT4 add_4679_2_lut (.I0(GND_net), .I1(n14_adj_3939), .I2(n83), 
            .I3(GND_net), .O(n8476[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4679_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4679_2 (.CI(GND_net), .I0(n14_adj_3939), .I1(n83), .CO(n26193));
    SB_LUT4 add_4678_22_lut (.I0(GND_net), .I1(n8476[19]), .I2(GND_net), 
            .I3(n26192), .O(n8453[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4678_21_lut (.I0(GND_net), .I1(n8476[18]), .I2(GND_net), 
            .I3(n26191), .O(n8453[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_21 (.CI(n26191), .I0(n8476[18]), .I1(GND_net), .CO(n26192));
    SB_LUT4 add_4678_20_lut (.I0(GND_net), .I1(n8476[17]), .I2(GND_net), 
            .I3(n26190), .O(n8453[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_20 (.CI(n26190), .I0(n8476[17]), .I1(GND_net), .CO(n26191));
    SB_LUT4 add_4678_19_lut (.I0(GND_net), .I1(n8476[16]), .I2(GND_net), 
            .I3(n26189), .O(n8453[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_19 (.CI(n26189), .I0(n8476[16]), .I1(GND_net), .CO(n26190));
    SB_LUT4 add_4678_18_lut (.I0(GND_net), .I1(n8476[15]), .I2(GND_net), 
            .I3(n26188), .O(n8453[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_18 (.CI(n26188), .I0(n8476[15]), .I1(GND_net), .CO(n26189));
    SB_LUT4 add_4678_17_lut (.I0(GND_net), .I1(n8476[14]), .I2(GND_net), 
            .I3(n26187), .O(n8453[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_17 (.CI(n26187), .I0(n8476[14]), .I1(GND_net), .CO(n26188));
    SB_LUT4 add_4678_16_lut (.I0(GND_net), .I1(n8476[13]), .I2(n1102), 
            .I3(n26186), .O(n8453[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_16 (.CI(n26186), .I0(n8476[13]), .I1(n1102), .CO(n26187));
    SB_LUT4 add_4678_15_lut (.I0(GND_net), .I1(n8476[12]), .I2(n1029), 
            .I3(n26185), .O(n8453[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_15 (.CI(n26185), .I0(n8476[12]), .I1(n1029), .CO(n26186));
    SB_LUT4 add_4678_14_lut (.I0(GND_net), .I1(n8476[11]), .I2(n956), 
            .I3(n26184), .O(n8453[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_14 (.CI(n26184), .I0(n8476[11]), .I1(n956), .CO(n26185));
    SB_LUT4 add_4678_13_lut (.I0(GND_net), .I1(n8476[10]), .I2(n883), 
            .I3(n26183), .O(n8453[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_13 (.CI(n26183), .I0(n8476[10]), .I1(n883), .CO(n26184));
    SB_LUT4 add_4678_12_lut (.I0(GND_net), .I1(n8476[9]), .I2(n810), .I3(n26182), 
            .O(n8453[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_12 (.CI(n26182), .I0(n8476[9]), .I1(n810), .CO(n26183));
    SB_LUT4 add_4678_11_lut (.I0(GND_net), .I1(n8476[8]), .I2(n737), .I3(n26181), 
            .O(n8453[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_11 (.CI(n26181), .I0(n8476[8]), .I1(n737), .CO(n26182));
    SB_LUT4 add_4678_10_lut (.I0(GND_net), .I1(n8476[7]), .I2(n664), .I3(n26180), 
            .O(n8453[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_10 (.CI(n26180), .I0(n8476[7]), .I1(n664), .CO(n26181));
    SB_LUT4 add_4678_9_lut (.I0(GND_net), .I1(n8476[6]), .I2(n591), .I3(n26179), 
            .O(n8453[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_9 (.CI(n26179), .I0(n8476[6]), .I1(n591), .CO(n26180));
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3392[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_4678_8_lut (.I0(GND_net), .I1(n8476[5]), .I2(n518), .I3(n26178), 
            .O(n8453[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20542_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n24625));   // verilog/motorControl.v(34[16:22])
    defparam i20542_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4080));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20540_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n8417[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20540_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i17460_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17460_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4678_8 (.CI(n26178), .I0(n8476[5]), .I1(n518), .CO(n26179));
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_563_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n2629[7]), .I3(n24847), .O(\PID_CONTROLLER.integral_23__N_3416 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4678_7_lut (.I0(GND_net), .I1(n8476[4]), .I2(n445), .I3(n26177), 
            .O(n8453[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_7 (.CI(n26177), .I0(n8476[4]), .I1(n445), .CO(n26178));
    SB_LUT4 i2_3_lut_4_lut_adj_1479 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n8411[0]), 
            .I3(n24548), .O(n8404[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1479.LUT_INIT = 16'h8778;
    SB_LUT4 i20509_2_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(\Kp[1] ), 
            .I3(n1[19]), .O(n8411[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20509_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i20483_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n24548), 
            .I3(n8411[0]), .O(n4_adj_4128));   // verilog/motorControl.v(34[16:22])
    defparam i20483_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_4678_6_lut (.I0(GND_net), .I1(n8476[3]), .I2(n372), .I3(n26176), 
            .O(n8453[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_6 (.CI(n26176), .I0(n8476[3]), .I1(n372), .CO(n26177));
    SB_LUT4 add_4678_5_lut (.I0(GND_net), .I1(n8476[2]), .I2(n299), .I3(n26175), 
            .O(n8453[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_5 (.CI(n26175), .I0(n8476[2]), .I1(n299), .CO(n26176));
    SB_LUT4 add_4678_4_lut (.I0(GND_net), .I1(n8476[1]), .I2(n226), .I3(n26174), 
            .O(n8453[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n24906), 
            .O(duty_23__N_3516[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20472_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n24548));   // verilog/motorControl.v(34[16:22])
    defparam i20472_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_4678_4 (.CI(n26174), .I0(n8476[1]), .I1(n226), .CO(n26175));
    SB_LUT4 add_4678_3_lut (.I0(GND_net), .I1(n8476[0]), .I2(n153), .I3(n26173), 
            .O(n8453[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n25042), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n25043));
    SB_CARRY add_4678_3 (.CI(n26173), .I0(n8476[0]), .I1(n153), .CO(n26174));
    SB_LUT4 add_4678_2_lut (.I0(GND_net), .I1(n11_adj_3934), .I2(n80), 
            .I3(GND_net), .O(n8453[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_2 (.CI(GND_net), .I0(n11_adj_3934), .I1(n80), .CO(n26173));
    SB_LUT4 i20470_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n8404[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20470_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3416 [23]), 
            .I1(n8429[21]), .I2(GND_net), .I3(n26172), .O(n6842[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n8429[20]), .I2(GND_net), 
            .I3(n26171), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n24906), .I0(n106[5]), .I1(n155[5]), .CO(n24907));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n25041), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n26171), .I0(n8429[20]), .I1(GND_net), 
            .CO(n26172));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n8429[19]), .I2(GND_net), 
            .I3(n26170), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n26170), .I0(n8429[19]), .I1(GND_net), 
            .CO(n26171));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n8429[18]), .I2(GND_net), 
            .I3(n26169), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n26169), .I0(n8429[18]), .I1(GND_net), 
            .CO(n26170));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n8429[17]), .I2(GND_net), 
            .I3(n26168), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[12]), 
            .I3(n25111), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n25111), .I0(GND_net), .I1(n1_adj_4337[12]), 
            .CO(n25112));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n24905), 
            .O(duty_23__N_3516[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n26168), .I0(n8429[17]), .I1(GND_net), 
            .CO(n26169));
    SB_CARRY sub_3_add_2_13 (.CI(n25041), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n25042));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n8429[16]), .I2(GND_net), 
            .I3(n26167), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n26167), .I0(n8429[16]), .I1(GND_net), 
            .CO(n26168));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n8429[15]), .I2(GND_net), 
            .I3(n26166), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n26166), .I0(n8429[15]), .I1(GND_net), 
            .CO(n26167));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n8429[14]), .I2(GND_net), 
            .I3(n26165), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n26165), .I0(n8429[14]), .I1(GND_net), 
            .CO(n26166));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n8429[13]), .I2(n1096), 
            .I3(n26164), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n25040), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[11]), 
            .I3(n25110), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n26164), .I0(n8429[13]), .I1(n1096), 
            .CO(n26165));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n8429[12]), .I2(n1023), 
            .I3(n26163), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n26163), .I0(n8429[12]), .I1(n1023), 
            .CO(n26164));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n8429[11]), .I2(n950), 
            .I3(n26162), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n26162), .I0(n8429[11]), .I1(n950), 
            .CO(n26163));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n8429[10]), .I2(n877), 
            .I3(n26161), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n26161), .I0(n8429[10]), .I1(n877), 
            .CO(n26162));
    SB_CARRY sub_3_add_2_12 (.CI(n25040), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n25041));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n8429[9]), .I2(n804), 
            .I3(n26160), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n26160), .I0(n8429[9]), .I1(n804), 
            .CO(n26161));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n8429[8]), .I2(n731), 
            .I3(n26159), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n26159), .I0(n8429[8]), .I1(n731), 
            .CO(n26160));
    SB_LUT4 i27763_3_lut (.I0(n11_adj_4061), .I1(n9_adj_4132), .I2(n33440), 
            .I3(GND_net), .O(n33437));
    defparam i27763_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n25039), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n8429[7]), .I2(n658), 
            .I3(n26158), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n26158), .I0(n8429[7]), .I1(n658), 
            .CO(n26159));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n8429[6]), .I2(n585), 
            .I3(n26157), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n26157), .I0(n8429[6]), .I1(n585), 
            .CO(n26158));
    SB_LUT4 i20522_3_lut_4_lut (.I0(n62_adj_4133), .I1(n131_adj_4134), .I2(n204), 
            .I3(n8417[0]), .O(n4_adj_3913));   // verilog/motorControl.v(34[16:22])
    defparam i20522_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n8429[5]), .I2(n512), 
            .I3(n26156), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1480 (.I0(n62_adj_4133), .I1(n131_adj_4134), 
            .I2(n8417[0]), .I3(n204), .O(n8411[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1480.LUT_INIT = 16'h8778;
    SB_CARRY mult_11_add_1225_8 (.CI(n26156), .I0(n8429[5]), .I1(n512), 
            .CO(n26157));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n8429[4]), .I2(n439), 
            .I3(n26155), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n25110), .I0(GND_net), .I1(n1_adj_4337[11]), 
            .CO(n25111));
    SB_CARRY mult_11_add_1225_7 (.CI(n26155), .I0(n8429[4]), .I1(n439), 
            .CO(n26156));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n8429[3]), .I2(n366), 
            .I3(n26154), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n26154), .I0(n8429[3]), .I1(n366), 
            .CO(n26155));
    SB_CARRY add_12_6 (.CI(n24905), .I0(n106[4]), .I1(n155[4]), .CO(n24906));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n8429[2]), .I2(n293), 
            .I3(n26153), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n26153), .I0(n8429[2]), .I1(n293), 
            .CO(n26154));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n8429[1]), .I2(n220), 
            .I3(n26152), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n26152), .I0(n8429[1]), .I1(n220), 
            .CO(n26153));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n8429[0]), .I2(n147), 
            .I3(n26151), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n26151), .I0(n8429[0]), .I1(n147), 
            .CO(n26152));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_3927), .I2(n74), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_3927), .I1(n74), 
            .CO(n26151));
    SB_LUT4 add_4677_23_lut (.I0(GND_net), .I1(n8453[20]), .I2(GND_net), 
            .I3(n26150), .O(n8429[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[10]), 
            .I3(n25109), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_22_lut (.I0(GND_net), .I1(n8453[19]), .I2(GND_net), 
            .I3(n26149), .O(n8429[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_22 (.CI(n26149), .I0(n8453[19]), .I1(GND_net), .CO(n26150));
    SB_CARRY unary_minus_16_add_3_12 (.CI(n25109), .I0(GND_net), .I1(n1_adj_4337[10]), 
            .CO(n25110));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[9]), 
            .I3(n25108), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n25108), .I0(GND_net), .I1(n1_adj_4337[9]), 
            .CO(n25109));
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n24904), 
            .O(duty_23__N_3516[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_11 (.CI(n25039), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n25040));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n25038), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[8]), 
            .I3(n25107), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_5 (.CI(n24904), .I0(n106[3]), .I1(n155[3]), .CO(n24905));
    SB_CARRY unary_minus_16_add_3_10 (.CI(n25107), .I0(GND_net), .I1(n1_adj_4337[8]), 
            .CO(n25108));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[7]), 
            .I3(n25106), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n24903), 
            .O(duty_23__N_3516[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n25038), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n25039));
    SB_LUT4 add_4677_21_lut (.I0(GND_net), .I1(n8453[18]), .I2(GND_net), 
            .I3(n26148), .O(n8429[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_21 (.CI(n26148), .I0(n8453[18]), .I1(GND_net), .CO(n26149));
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n25037), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_20_lut (.I0(GND_net), .I1(n8453[17]), .I2(GND_net), 
            .I3(n26147), .O(n8429[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_20 (.CI(n26147), .I0(n8453[17]), .I1(GND_net), .CO(n26148));
    SB_LUT4 add_4677_19_lut (.I0(GND_net), .I1(n8453[16]), .I2(GND_net), 
            .I3(n26146), .O(n8429[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_19 (.CI(n26146), .I0(n8453[16]), .I1(GND_net), .CO(n26147));
    SB_LUT4 add_4677_18_lut (.I0(GND_net), .I1(n8453[15]), .I2(GND_net), 
            .I3(n26145), .O(n8429[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_18 (.CI(n26145), .I0(n8453[15]), .I1(GND_net), .CO(n26146));
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4677_17_lut (.I0(GND_net), .I1(n8453[14]), .I2(GND_net), 
            .I3(n26144), .O(n8429[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_17 (.CI(n26144), .I0(n8453[14]), .I1(GND_net), .CO(n26145));
    SB_LUT4 add_4677_16_lut (.I0(GND_net), .I1(n8453[13]), .I2(n1099), 
            .I3(n26143), .O(n8429[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_16 (.CI(n26143), .I0(n8453[13]), .I1(n1099), .CO(n26144));
    SB_LUT4 add_4677_15_lut (.I0(GND_net), .I1(n8453[12]), .I2(n1026), 
            .I3(n26142), .O(n8429[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_15 (.CI(n26142), .I0(n8453[12]), .I1(n1026), .CO(n26143));
    SB_LUT4 add_4677_14_lut (.I0(GND_net), .I1(n8453[11]), .I2(n953), 
            .I3(n26141), .O(n8429[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_14 (.CI(n26141), .I0(n8453[11]), .I1(n953), .CO(n26142));
    SB_LUT4 add_4677_13_lut (.I0(GND_net), .I1(n8453[10]), .I2(n880), 
            .I3(n26140), .O(n8429[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_13 (.CI(n26140), .I0(n8453[10]), .I1(n880), .CO(n26141));
    SB_LUT4 add_4677_12_lut (.I0(GND_net), .I1(n8453[9]), .I2(n807), .I3(n26139), 
            .O(n8429[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_12 (.CI(n26139), .I0(n8453[9]), .I1(n807), .CO(n26140));
    SB_LUT4 add_4677_11_lut (.I0(GND_net), .I1(n8453[8]), .I2(n734), .I3(n26138), 
            .O(n8429[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_11 (.CI(n26138), .I0(n8453[8]), .I1(n734), .CO(n26139));
    SB_LUT4 add_4677_10_lut (.I0(GND_net), .I1(n8453[7]), .I2(n661), .I3(n26137), 
            .O(n8429[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_10 (.CI(n26137), .I0(n8453[7]), .I1(n661), .CO(n26138));
    SB_LUT4 add_4677_9_lut (.I0(GND_net), .I1(n8453[6]), .I2(n588), .I3(n26136), 
            .O(n8429[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_9 (.CI(n26136), .I0(n8453[6]), .I1(n588), .CO(n26137));
    SB_LUT4 add_4677_8_lut (.I0(GND_net), .I1(n8453[5]), .I2(n515), .I3(n26135), 
            .O(n8429[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_8 (.CI(n26135), .I0(n8453[5]), .I1(n515), .CO(n26136));
    SB_LUT4 add_4677_7_lut (.I0(GND_net), .I1(n8453[4]), .I2(n442), .I3(n26134), 
            .O(n8429[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_7 (.CI(n26134), .I0(n8453[4]), .I1(n442), .CO(n26135));
    SB_LUT4 add_4677_6_lut (.I0(GND_net), .I1(n8453[3]), .I2(n369), .I3(n26133), 
            .O(n8429[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_6 (.CI(n26133), .I0(n8453[3]), .I1(n369), .CO(n26134));
    SB_LUT4 add_4677_5_lut (.I0(GND_net), .I1(n8453[2]), .I2(n296), .I3(n26132), 
            .O(n8429[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_5 (.CI(n26132), .I0(n8453[2]), .I1(n296), .CO(n26133));
    SB_LUT4 add_4677_4_lut (.I0(GND_net), .I1(n8453[1]), .I2(n223), .I3(n26131), 
            .O(n8429[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_4 (.CI(n26131), .I0(n8453[1]), .I1(n223), .CO(n26132));
    SB_LUT4 add_4677_3_lut (.I0(GND_net), .I1(n8453[0]), .I2(n150), .I3(n26130), 
            .O(n8429[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_3 (.CI(n26130), .I0(n8453[0]), .I1(n150), .CO(n26131));
    SB_LUT4 add_4677_2_lut (.I0(GND_net), .I1(n8_adj_3918), .I2(n77), 
            .I3(GND_net), .O(n8429[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_2 (.CI(GND_net), .I0(n8_adj_3918), .I1(n77), .CO(n26130));
    SB_LUT4 add_4671_7_lut (.I0(GND_net), .I1(n30955), .I2(n490), .I3(n26129), 
            .O(n8396[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4671_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4671_6_lut (.I0(GND_net), .I1(n8404[3]), .I2(n417_adj_4136), 
            .I3(n26128), .O(n8396[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4671_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4671_6 (.CI(n26128), .I0(n8404[3]), .I1(n417_adj_4136), 
            .CO(n26129));
    SB_LUT4 add_4671_5_lut (.I0(GND_net), .I1(n8404[2]), .I2(n344_adj_4137), 
            .I3(n26127), .O(n8396[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4671_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4671_5 (.CI(n26127), .I0(n8404[2]), .I1(n344_adj_4137), 
            .CO(n26128));
    SB_LUT4 add_4671_4_lut (.I0(GND_net), .I1(n8404[1]), .I2(n271_adj_4138), 
            .I3(n26126), .O(n8396[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4671_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4671_4 (.CI(n26126), .I0(n8404[1]), .I1(n271_adj_4138), 
            .CO(n26127));
    SB_LUT4 add_4671_3_lut (.I0(GND_net), .I1(n8404[0]), .I2(n198_adj_4139), 
            .I3(n26125), .O(n8396[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4671_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4671_3 (.CI(n26125), .I0(n8404[0]), .I1(n198_adj_4139), 
            .CO(n26126));
    SB_LUT4 add_4671_2_lut (.I0(GND_net), .I1(n56_adj_4140), .I2(n125_adj_4141), 
            .I3(GND_net), .O(n8396[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4671_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4671_2 (.CI(GND_net), .I0(n56_adj_4140), .I1(n125_adj_4141), 
            .CO(n26125));
    SB_LUT4 add_4670_8_lut (.I0(GND_net), .I1(n8396[5]), .I2(n560_adj_4142), 
            .I3(n26124), .O(n8387[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4670_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4670_7_lut (.I0(GND_net), .I1(n8396[4]), .I2(n487_adj_4143), 
            .I3(n26123), .O(n8387[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4670_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4670_7 (.CI(n26123), .I0(n8396[4]), .I1(n487_adj_4143), 
            .CO(n26124));
    SB_LUT4 add_4670_6_lut (.I0(GND_net), .I1(n8396[3]), .I2(n414_adj_4144), 
            .I3(n26122), .O(n8387[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4670_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4670_6 (.CI(n26122), .I0(n8396[3]), .I1(n414_adj_4144), 
            .CO(n26123));
    SB_LUT4 add_4670_5_lut (.I0(GND_net), .I1(n8396[2]), .I2(n341_adj_4145), 
            .I3(n26121), .O(n8387[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4670_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4670_5 (.CI(n26121), .I0(n8396[2]), .I1(n341_adj_4145), 
            .CO(n26122));
    SB_LUT4 add_4670_4_lut (.I0(GND_net), .I1(n8396[1]), .I2(n268_adj_4146), 
            .I3(n26120), .O(n8387[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4670_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4670_4 (.CI(n26120), .I0(n8396[1]), .I1(n268_adj_4146), 
            .CO(n26121));
    SB_LUT4 add_4670_3_lut (.I0(GND_net), .I1(n8396[0]), .I2(n195_adj_4147), 
            .I3(n26119), .O(n8387[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4670_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4670_3 (.CI(n26119), .I0(n8396[0]), .I1(n195_adj_4147), 
            .CO(n26120));
    SB_CARRY unary_minus_16_add_3_9 (.CI(n25106), .I0(GND_net), .I1(n1_adj_4337[7]), 
            .CO(n25107));
    SB_LUT4 add_4670_2_lut (.I0(GND_net), .I1(n53_adj_4148), .I2(n122_adj_4149), 
            .I3(GND_net), .O(n8387[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4670_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4670_2 (.CI(GND_net), .I0(n53_adj_4148), .I1(n122_adj_4149), 
            .CO(n26119));
    SB_CARRY sub_3_add_2_9 (.CI(n25037), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n25038));
    SB_CARRY add_12_4 (.CI(n24903), .I0(n106[2]), .I1(n155[2]), .CO(n24904));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n25036), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_9_lut (.I0(GND_net), .I1(n8387[6]), .I2(n630_adj_4150), 
            .I3(n26118), .O(n8377[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_8_lut (.I0(GND_net), .I1(n8387[5]), .I2(n557_adj_4151), 
            .I3(n26117), .O(n8377[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_8 (.CI(n26117), .I0(n8387[5]), .I1(n557_adj_4151), 
            .CO(n26118));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[6]), 
            .I3(n25105), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n24902), 
            .O(duty_23__N_3516[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_7_lut (.I0(GND_net), .I1(n8387[4]), .I2(n484_adj_4154), 
            .I3(n26116), .O(n8377[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_7 (.CI(n26116), .I0(n8387[4]), .I1(n484_adj_4154), 
            .CO(n26117));
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4155));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4156));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_8 (.CI(n25036), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n25037));
    SB_CARRY unary_minus_16_add_3_8 (.CI(n25105), .I0(GND_net), .I1(n1_adj_4337[6]), 
            .CO(n25106));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[5]), 
            .I3(n25104), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n25104), .I0(GND_net), .I1(n1_adj_4337[5]), 
            .CO(n25105));
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4158));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n25035), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_7 (.CI(n25035), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n25036));
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n25034), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_3 (.CI(n24902), .I0(n106[1]), .I1(n155[1]), .CO(n24903));
    SB_LUT4 add_4669_6_lut (.I0(GND_net), .I1(n8387[3]), .I2(n411_adj_4159), 
            .I3(n26115), .O(n8377[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_6 (.CI(n26115), .I0(n8387[3]), .I1(n411_adj_4159), 
            .CO(n26116));
    SB_LUT4 add_4669_5_lut (.I0(GND_net), .I1(n8387[2]), .I2(n338_adj_4160), 
            .I3(n26114), .O(n8377[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_5 (.CI(n26114), .I0(n8387[2]), .I1(n338_adj_4160), 
            .CO(n26115));
    SB_CARRY sub_3_add_2_6 (.CI(n25034), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n25035));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[4]), 
            .I3(n25103), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n25103), .I0(GND_net), .I1(n1_adj_4337[4]), 
            .CO(n25104));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3516[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n25033), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_5 (.CI(n25033), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n25034));
    SB_LUT4 add_4669_4_lut (.I0(GND_net), .I1(n8387[1]), .I2(n265_adj_4162), 
            .I3(n26113), .O(n8377[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[3]), 
            .I3(n25102), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n24902));
    SB_CARRY unary_minus_16_add_3_5 (.CI(n25102), .I0(GND_net), .I1(n1_adj_4337[3]), 
            .CO(n25103));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[2]), 
            .I3(n25101), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_4 (.CI(n26113), .I0(n8387[1]), .I1(n265_adj_4162), 
            .CO(n26114));
    SB_LUT4 add_4669_3_lut (.I0(GND_net), .I1(n8387[0]), .I2(n192_adj_4165), 
            .I3(n26112), .O(n8377[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_3 (.CI(n26112), .I0(n8387[0]), .I1(n192_adj_4165), 
            .CO(n26113));
    SB_LUT4 add_4669_2_lut (.I0(GND_net), .I1(n50_adj_4166), .I2(n119_adj_4167), 
            .I3(GND_net), .O(n8377[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_2 (.CI(GND_net), .I0(n50_adj_4166), .I1(n119_adj_4167), 
            .CO(n26112));
    SB_LUT4 add_4668_10_lut (.I0(GND_net), .I1(n8377[7]), .I2(n700_adj_4168), 
            .I3(n26111), .O(n8366[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4668_9_lut (.I0(GND_net), .I1(n8377[6]), .I2(n627_adj_4169), 
            .I3(n26110), .O(n8366[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4668_9 (.CI(n26110), .I0(n8377[6]), .I1(n627_adj_4169), 
            .CO(n26111));
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n25032), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4668_8_lut (.I0(GND_net), .I1(n8377[5]), .I2(n554_adj_4170), 
            .I3(n26109), .O(n8366[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4668_8 (.CI(n26109), .I0(n8377[5]), .I1(n554_adj_4170), 
            .CO(n26110));
    SB_CARRY unary_minus_16_add_3_4 (.CI(n25101), .I0(GND_net), .I1(n1_adj_4337[2]), 
            .CO(n25102));
    SB_LUT4 add_4668_7_lut (.I0(GND_net), .I1(n8377[4]), .I2(n481_adj_4171), 
            .I3(n26108), .O(n8366[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4668_7 (.CI(n26108), .I0(n8377[4]), .I1(n481_adj_4171), 
            .CO(n26109));
    SB_LUT4 add_4668_6_lut (.I0(GND_net), .I1(n8377[3]), .I2(n408_adj_4172), 
            .I3(n26107), .O(n8366[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4668_6 (.CI(n26107), .I0(n8377[3]), .I1(n408_adj_4172), 
            .CO(n26108));
    SB_LUT4 add_4668_5_lut (.I0(GND_net), .I1(n8377[2]), .I2(n335_adj_4173), 
            .I3(n26106), .O(n8366[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4668_5 (.CI(n26106), .I0(n8377[2]), .I1(n335_adj_4173), 
            .CO(n26107));
    SB_LUT4 add_4668_4_lut (.I0(GND_net), .I1(n8377[1]), .I2(n262_adj_4174), 
            .I3(n26105), .O(n8366[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4337[1]), 
            .I3(n25100), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4668_4 (.CI(n26105), .I0(n8377[1]), .I1(n262_adj_4174), 
            .CO(n26106));
    SB_CARRY sub_3_add_2_4 (.CI(n25032), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n25033));
    SB_CARRY unary_minus_16_add_3_3 (.CI(n25100), .I0(GND_net), .I1(n1_adj_4337[1]), 
            .CO(n25101));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n25031), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n25031), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n25032));
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n18701), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4668_3_lut (.I0(GND_net), .I1(n8377[0]), .I2(n189_adj_4176), 
            .I3(n26104), .O(n8366[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n18701), 
            .CO(n25100));
    SB_CARRY add_4668_3 (.CI(n26104), .I0(n8377[0]), .I1(n189_adj_4176), 
            .CO(n26105));
    SB_LUT4 add_4668_2_lut (.I0(GND_net), .I1(n47_adj_4177), .I2(n116_adj_4178), 
            .I3(GND_net), .O(n8366[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4668_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4668_2 (.CI(GND_net), .I0(n47_adj_4177), .I1(n116_adj_4178), 
            .CO(n26104));
    SB_LUT4 add_4667_11_lut (.I0(GND_net), .I1(n8366[8]), .I2(n770_adj_4179), 
            .I3(n26103), .O(n8354[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4338[23]), 
            .I3(n25099), .O(\PID_CONTROLLER.integral_23__N_3467 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4667_10_lut (.I0(GND_net), .I1(n8366[7]), .I2(n697_adj_4181), 
            .I3(n26102), .O(n8354[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_10 (.CI(n26102), .I0(n8366[7]), .I1(n697_adj_4181), 
            .CO(n26103));
    SB_LUT4 add_4667_9_lut (.I0(GND_net), .I1(n8366[6]), .I2(n624_adj_4182), 
            .I3(n26101), .O(n8354[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_9 (.CI(n26101), .I0(n8366[6]), .I1(n624_adj_4182), 
            .CO(n26102));
    SB_LUT4 add_4667_8_lut (.I0(GND_net), .I1(n8366[5]), .I2(n551_adj_4183), 
            .I3(n26100), .O(n8354[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_8 (.CI(n26100), .I0(n8366[5]), .I1(n551_adj_4183), 
            .CO(n26101));
    SB_LUT4 add_4667_7_lut (.I0(GND_net), .I1(n8366[4]), .I2(n478_adj_4184), 
            .I3(n26099), .O(n8354[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_7 (.CI(n26099), .I0(n8366[4]), .I1(n478_adj_4184), 
            .CO(n26100));
    SB_LUT4 add_4667_6_lut (.I0(GND_net), .I1(n8366[3]), .I2(n405_adj_4185), 
            .I3(n26098), .O(n8354[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_6 (.CI(n26098), .I0(n8366[3]), .I1(n405_adj_4185), 
            .CO(n26099));
    SB_LUT4 add_4667_5_lut (.I0(GND_net), .I1(n8366[2]), .I2(n332_adj_4186), 
            .I3(n26097), .O(n8354[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_5 (.CI(n26097), .I0(n8366[2]), .I1(n332_adj_4186), 
            .CO(n26098));
    SB_LUT4 add_4667_4_lut (.I0(GND_net), .I1(n8366[1]), .I2(n259_adj_4187), 
            .I3(n26096), .O(n8354[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28123_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n35239), 
            .I2(IntegralLimit[7]), .I3(n33437), .O(n33799));
    defparam i28123_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_4667_4 (.CI(n26096), .I0(n8366[1]), .I1(n259_adj_4187), 
            .CO(n26097));
    SB_LUT4 add_4667_3_lut (.I0(GND_net), .I1(n8366[0]), .I2(n186_adj_4188), 
            .I3(n26095), .O(n8354[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n25031));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4338[22]), .I3(n25098), .O(n45_adj_4035)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n25098), .I0(GND_net), .I1(n1_adj_4338[22]), 
            .CO(n25099));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4338[21]), .I3(n25097), .O(n43_adj_4009)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4667_3 (.CI(n26095), .I0(n8366[0]), .I1(n186_adj_4188), 
            .CO(n26096));
    SB_LUT4 add_4667_2_lut (.I0(GND_net), .I1(n44_adj_4191), .I2(n113_adj_4192), 
            .I3(GND_net), .O(n8354[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_2 (.CI(GND_net), .I0(n44_adj_4191), .I1(n113_adj_4192), 
            .CO(n26095));
    SB_LUT4 add_4666_12_lut (.I0(GND_net), .I1(n8354[9]), .I2(n840_adj_4193), 
            .I3(n26094), .O(n8341[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4666_11_lut (.I0(GND_net), .I1(n8354[8]), .I2(n767_adj_4194), 
            .I3(n26093), .O(n8341[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_11 (.CI(n26093), .I0(n8354[8]), .I1(n767_adj_4194), 
            .CO(n26094));
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4195));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4666_10_lut (.I0(GND_net), .I1(n8354[7]), .I2(n694_adj_4196), 
            .I3(n26092), .O(n8341[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28003_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4197), 
            .I2(IntegralLimit[9]), .I3(n33799), .O(n33679));
    defparam i28003_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_4666_10 (.CI(n26092), .I0(n8354[7]), .I1(n694_adj_4196), 
            .CO(n26093));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n25097), .I0(GND_net), .I1(n1_adj_4338[21]), 
            .CO(n25098));
    SB_LUT4 add_4666_9_lut (.I0(GND_net), .I1(n8354[6]), .I2(n621_adj_4198), 
            .I3(n26091), .O(n8341[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_9 (.CI(n26091), .I0(n8354[6]), .I1(n621_adj_4198), 
            .CO(n26092));
    SB_LUT4 add_4666_8_lut (.I0(GND_net), .I1(n8354[5]), .I2(n548_adj_4199), 
            .I3(n26090), .O(n8341[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_8 (.CI(n26090), .I0(n8354[5]), .I1(n548_adj_4199), 
            .CO(n26091));
    SB_LUT4 add_4666_7_lut (.I0(GND_net), .I1(n8354[4]), .I2(n475_adj_4200), 
            .I3(n26089), .O(n8341[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_7 (.CI(n26089), .I0(n8354[4]), .I1(n475_adj_4200), 
            .CO(n26090));
    SB_LUT4 add_4666_6_lut (.I0(GND_net), .I1(n8354[3]), .I2(n402_adj_4201), 
            .I3(n26088), .O(n8341[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_6 (.CI(n26088), .I0(n8354[3]), .I1(n402_adj_4201), 
            .CO(n26089));
    SB_LUT4 add_4666_5_lut (.I0(GND_net), .I1(n8354[2]), .I2(n329_adj_4202), 
            .I3(n26087), .O(n8341[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_5 (.CI(n26087), .I0(n8354[2]), .I1(n329_adj_4202), 
            .CO(n26088));
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4203));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4666_4_lut (.I0(GND_net), .I1(n8354[1]), .I2(n256_adj_4204), 
            .I3(n26086), .O(n8341[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_4 (.CI(n26086), .I0(n8354[1]), .I1(n256_adj_4204), 
            .CO(n26087));
    SB_LUT4 add_4666_3_lut (.I0(GND_net), .I1(n8354[0]), .I2(n183_adj_4205), 
            .I3(n26085), .O(n8341[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_3 (.CI(n26085), .I0(n8354[0]), .I1(n183_adj_4205), 
            .CO(n26086));
    SB_LUT4 add_4666_2_lut (.I0(GND_net), .I1(n41_adj_4206), .I2(n110_adj_4207), 
            .I3(GND_net), .O(n8341[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4666_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4666_2 (.CI(GND_net), .I0(n41_adj_4206), .I1(n110_adj_4207), 
            .CO(n26085));
    SB_LUT4 add_4665_13_lut (.I0(GND_net), .I1(n8341[10]), .I2(n910_adj_4208), 
            .I3(n26084), .O(n8327[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4665_12_lut (.I0(GND_net), .I1(n8341[9]), .I2(n837_adj_4209), 
            .I3(n26083), .O(n8327[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_12 (.CI(n26083), .I0(n8341[9]), .I1(n837_adj_4209), 
            .CO(n26084));
    SB_LUT4 add_4665_11_lut (.I0(GND_net), .I1(n8341[8]), .I2(n764_adj_4210), 
            .I3(n26082), .O(n8327[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_11 (.CI(n26082), .I0(n8341[8]), .I1(n764_adj_4210), 
            .CO(n26083));
    SB_LUT4 add_4665_10_lut (.I0(GND_net), .I1(n8341[7]), .I2(n691_adj_4211), 
            .I3(n26081), .O(n8327[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_10 (.CI(n26081), .I0(n8341[7]), .I1(n691_adj_4211), 
            .CO(n26082));
    SB_LUT4 add_4665_9_lut (.I0(GND_net), .I1(n8341[6]), .I2(n618_adj_4212), 
            .I3(n26080), .O(n8327[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_9 (.CI(n26080), .I0(n8341[6]), .I1(n618_adj_4212), 
            .CO(n26081));
    SB_LUT4 add_4665_8_lut (.I0(GND_net), .I1(n8341[5]), .I2(n545_adj_4213), 
            .I3(n26079), .O(n8327[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4214));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4665_8 (.CI(n26079), .I0(n8341[5]), .I1(n545_adj_4213), 
            .CO(n26080));
    SB_LUT4 add_4665_7_lut (.I0(GND_net), .I1(n8341[4]), .I2(n472_adj_4215), 
            .I3(n26078), .O(n8327[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_7 (.CI(n26078), .I0(n8341[4]), .I1(n472_adj_4215), 
            .CO(n26079));
    SB_LUT4 add_4665_6_lut (.I0(GND_net), .I1(n8341[3]), .I2(n399_adj_4216), 
            .I3(n26077), .O(n8327[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_6 (.CI(n26077), .I0(n8341[3]), .I1(n399_adj_4216), 
            .CO(n26078));
    SB_LUT4 add_4665_5_lut (.I0(GND_net), .I1(n8341[2]), .I2(n326_adj_4217), 
            .I3(n26076), .O(n8327[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_5 (.CI(n26076), .I0(n8341[2]), .I1(n326_adj_4217), 
            .CO(n26077));
    SB_LUT4 add_4665_4_lut (.I0(GND_net), .I1(n8341[1]), .I2(n253_adj_4218), 
            .I3(n26075), .O(n8327[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_4 (.CI(n26075), .I0(n8341[1]), .I1(n253_adj_4218), 
            .CO(n26076));
    SB_LUT4 add_4665_3_lut (.I0(GND_net), .I1(n8341[0]), .I2(n180_adj_4219), 
            .I3(n26074), .O(n8327[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_3 (.CI(n26074), .I0(n8341[0]), .I1(n180_adj_4219), 
            .CO(n26075));
    SB_LUT4 add_4665_2_lut (.I0(GND_net), .I1(n38_adj_4220), .I2(n107_adj_4221), 
            .I3(GND_net), .O(n8327[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4665_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4665_2 (.CI(GND_net), .I0(n38_adj_4220), .I1(n107_adj_4221), 
            .CO(n26074));
    SB_LUT4 add_4664_14_lut (.I0(GND_net), .I1(n8327[11]), .I2(n980_adj_4222), 
            .I3(n26073), .O(n8312[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4664_13_lut (.I0(GND_net), .I1(n8327[10]), .I2(n907_adj_4223), 
            .I3(n26072), .O(n8312[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_13 (.CI(n26072), .I0(n8327[10]), .I1(n907_adj_4223), 
            .CO(n26073));
    SB_LUT4 add_4664_12_lut (.I0(GND_net), .I1(n8327[9]), .I2(n834_adj_4224), 
            .I3(n26071), .O(n8312[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_12 (.CI(n26071), .I0(n8327[9]), .I1(n834_adj_4224), 
            .CO(n26072));
    SB_LUT4 add_4664_11_lut (.I0(GND_net), .I1(n8327[8]), .I2(n761_adj_4225), 
            .I3(n26070), .O(n8312[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_11 (.CI(n26070), .I0(n8327[8]), .I1(n761_adj_4225), 
            .CO(n26071));
    SB_LUT4 add_4664_10_lut (.I0(GND_net), .I1(n8327[7]), .I2(n688_adj_4226), 
            .I3(n26069), .O(n8312[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_10 (.CI(n26069), .I0(n8327[7]), .I1(n688_adj_4226), 
            .CO(n26070));
    SB_LUT4 add_4664_9_lut (.I0(GND_net), .I1(n8327[6]), .I2(n615_adj_4227), 
            .I3(n26068), .O(n8312[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_9 (.CI(n26068), .I0(n8327[6]), .I1(n615_adj_4227), 
            .CO(n26069));
    SB_LUT4 add_4664_8_lut (.I0(GND_net), .I1(n8327[5]), .I2(n542_adj_4228), 
            .I3(n26067), .O(n8312[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_8 (.CI(n26067), .I0(n8327[5]), .I1(n542_adj_4228), 
            .CO(n26068));
    SB_LUT4 add_4664_7_lut (.I0(GND_net), .I1(n8327[4]), .I2(n469_adj_4229), 
            .I3(n26066), .O(n8312[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_7 (.CI(n26066), .I0(n8327[4]), .I1(n469_adj_4229), 
            .CO(n26067));
    SB_LUT4 add_4664_6_lut (.I0(GND_net), .I1(n8327[3]), .I2(n396_adj_4230), 
            .I3(n26065), .O(n8312[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_6 (.CI(n26065), .I0(n8327[3]), .I1(n396_adj_4230), 
            .CO(n26066));
    SB_LUT4 add_4664_5_lut (.I0(GND_net), .I1(n8327[2]), .I2(n323_adj_4231), 
            .I3(n26064), .O(n8312[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_5 (.CI(n26064), .I0(n8327[2]), .I1(n323_adj_4231), 
            .CO(n26065));
    SB_LUT4 add_4664_4_lut (.I0(GND_net), .I1(n8327[1]), .I2(n250_adj_4232), 
            .I3(n26063), .O(n8312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_4 (.CI(n26063), .I0(n8327[1]), .I1(n250_adj_4232), 
            .CO(n26064));
    SB_LUT4 add_4664_3_lut (.I0(GND_net), .I1(n8327[0]), .I2(n177_adj_4233), 
            .I3(n26062), .O(n8312[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4338[20]), .I3(n25096), .O(n41_adj_4124)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4664_3 (.CI(n26062), .I0(n8327[0]), .I1(n177_adj_4233), 
            .CO(n26063));
    SB_LUT4 add_4664_2_lut (.I0(GND_net), .I1(n35_adj_4235), .I2(n104_adj_4236), 
            .I3(GND_net), .O(n8312[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4664_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4664_2 (.CI(GND_net), .I0(n35_adj_4235), .I1(n104_adj_4236), 
            .CO(n26062));
    SB_LUT4 add_4663_15_lut (.I0(GND_net), .I1(n8312[12]), .I2(n1050_adj_4237), 
            .I3(n26061), .O(n8296[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4663_14_lut (.I0(GND_net), .I1(n8312[11]), .I2(n977_adj_4238), 
            .I3(n26060), .O(n8296[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_14 (.CI(n26060), .I0(n8312[11]), .I1(n977_adj_4238), 
            .CO(n26061));
    SB_LUT4 add_4663_13_lut (.I0(GND_net), .I1(n8312[10]), .I2(n904_adj_4239), 
            .I3(n26059), .O(n8296[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_13 (.CI(n26059), .I0(n8312[10]), .I1(n904_adj_4239), 
            .CO(n26060));
    SB_LUT4 add_4663_12_lut (.I0(GND_net), .I1(n8312[9]), .I2(n831_adj_4240), 
            .I3(n26058), .O(n8296[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_12 (.CI(n26058), .I0(n8312[9]), .I1(n831_adj_4240), 
            .CO(n26059));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n25096), .I0(GND_net), .I1(n1_adj_4338[20]), 
            .CO(n25097));
    SB_LUT4 add_4663_11_lut (.I0(GND_net), .I1(n8312[8]), .I2(n758_adj_4241), 
            .I3(n26057), .O(n8296[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_11 (.CI(n26057), .I0(n8312[8]), .I1(n758_adj_4241), 
            .CO(n26058));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4338[19]), .I3(n25095), .O(n39_adj_4121)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4663_10_lut (.I0(GND_net), .I1(n8312[7]), .I2(n685_adj_4243), 
            .I3(n26056), .O(n8296[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_10 (.CI(n26056), .I0(n8312[7]), .I1(n685_adj_4243), 
            .CO(n26057));
    SB_LUT4 add_4663_9_lut (.I0(GND_net), .I1(n8312[6]), .I2(n612_adj_4244), 
            .I3(n26055), .O(n8296[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_9 (.CI(n26055), .I0(n8312[6]), .I1(n612_adj_4244), 
            .CO(n26056));
    SB_LUT4 add_4663_8_lut (.I0(GND_net), .I1(n8312[5]), .I2(n539_adj_4245), 
            .I3(n26054), .O(n8296[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_8 (.CI(n26054), .I0(n8312[5]), .I1(n539_adj_4245), 
            .CO(n26055));
    SB_CARRY unary_minus_5_add_3_21 (.CI(n25095), .I0(GND_net), .I1(n1_adj_4338[19]), 
            .CO(n25096));
    SB_LUT4 add_4663_7_lut (.I0(GND_net), .I1(n8312[4]), .I2(n466_adj_4246), 
            .I3(n26053), .O(n8296[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_7 (.CI(n26053), .I0(n8312[4]), .I1(n466_adj_4246), 
            .CO(n26054));
    SB_LUT4 add_4663_6_lut (.I0(GND_net), .I1(n8312[3]), .I2(n393_adj_4247), 
            .I3(n26052), .O(n8296[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_6 (.CI(n26052), .I0(n8312[3]), .I1(n393_adj_4247), 
            .CO(n26053));
    SB_LUT4 add_4663_5_lut (.I0(GND_net), .I1(n8312[2]), .I2(n320_adj_4248), 
            .I3(n26051), .O(n8296[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_5 (.CI(n26051), .I0(n8312[2]), .I1(n320_adj_4248), 
            .CO(n26052));
    SB_LUT4 add_4663_4_lut (.I0(GND_net), .I1(n8312[1]), .I2(n247_adj_4249), 
            .I3(n26050), .O(n8296[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_4 (.CI(n26050), .I0(n8312[1]), .I1(n247_adj_4249), 
            .CO(n26051));
    SB_LUT4 add_4663_3_lut (.I0(GND_net), .I1(n8312[0]), .I2(n174_adj_4250), 
            .I3(n26049), .O(n8296[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4663_3 (.CI(n26049), .I0(n8312[0]), .I1(n174_adj_4250), 
            .CO(n26050));
    SB_LUT4 add_4663_2_lut (.I0(GND_net), .I1(n32_adj_4251), .I2(n101_adj_4252), 
            .I3(GND_net), .O(n8296[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4663_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4663_2 (.CI(GND_net), .I0(n32_adj_4251), .I1(n101_adj_4252), 
            .CO(n26049));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4338[18]), .I3(n25094), .O(n37_adj_4058)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4662_16_lut (.I0(GND_net), .I1(n8296[13]), .I2(n1120_adj_4255), 
            .I3(n26048), .O(n8279[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n25094), .I0(GND_net), .I1(n1_adj_4338[18]), 
            .CO(n25095));
    SB_LUT4 add_4662_15_lut (.I0(GND_net), .I1(n8296[12]), .I2(n1047_adj_4256), 
            .I3(n26047), .O(n8279[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n2629[6]), .I3(n24846), .O(\PID_CONTROLLER.integral_23__N_3416 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_15 (.CI(n26047), .I0(n8296[12]), .I1(n1047_adj_4256), 
            .CO(n26048));
    SB_LUT4 add_4662_14_lut (.I0(GND_net), .I1(n8296[11]), .I2(n974_adj_4257), 
            .I3(n26046), .O(n8279[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n2629[23]), .I3(n24863), .O(\PID_CONTROLLER.integral_23__N_3416 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4258));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4662_14 (.CI(n26046), .I0(n8296[11]), .I1(n974_adj_4257), 
            .CO(n26047));
    SB_LUT4 add_4662_13_lut (.I0(GND_net), .I1(n8296[10]), .I2(n901_adj_4259), 
            .I3(n26045), .O(n8279[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_13 (.CI(n26045), .I0(n8296[10]), .I1(n901_adj_4259), 
            .CO(n26046));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4338[17]), .I3(n25093), .O(n35_adj_4059)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4662_12_lut (.I0(GND_net), .I1(n8296[9]), .I2(n828_adj_4261), 
            .I3(n26044), .O(n8279[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_12 (.CI(n26044), .I0(n8296[9]), .I1(n828_adj_4261), 
            .CO(n26045));
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3392[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_4662_11_lut (.I0(GND_net), .I1(n8296[8]), .I2(n755_adj_4262), 
            .I3(n26043), .O(n8279[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_11 (.CI(n26043), .I0(n8296[8]), .I1(n755_adj_4262), 
            .CO(n26044));
    SB_CARRY unary_minus_5_add_3_19 (.CI(n25093), .I0(GND_net), .I1(n1_adj_4338[17]), 
            .CO(n25094));
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4263));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4662_10_lut (.I0(GND_net), .I1(n8296[7]), .I2(n682_adj_4264), 
            .I3(n26042), .O(n8279[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_10 (.CI(n26042), .I0(n8296[7]), .I1(n682_adj_4264), 
            .CO(n26043));
    SB_LUT4 add_563_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n2629[22]), .I3(n24862), .O(\PID_CONTROLLER.integral_23__N_3416 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4265));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4662_9_lut (.I0(GND_net), .I1(n8296[6]), .I2(n609_adj_4266), 
            .I3(n26041), .O(n8279[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4267));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4268));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4662_9 (.CI(n26041), .I0(n8296[6]), .I1(n609_adj_4266), 
            .CO(n26042));
    SB_LUT4 add_4662_8_lut (.I0(GND_net), .I1(n8296[5]), .I2(n536_adj_4269), 
            .I3(n26040), .O(n8279[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_8 (.CI(n26040), .I0(n8296[5]), .I1(n536_adj_4269), 
            .CO(n26041));
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4270));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4662_7_lut (.I0(GND_net), .I1(n8296[4]), .I2(n463_adj_4271), 
            .I3(n26039), .O(n8279[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_49_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n35222));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_49_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_563_24 (.CI(n24862), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n2629[22]), .CO(n24863));
    SB_CARRY add_4662_7 (.CI(n26039), .I0(n8296[4]), .I1(n463_adj_4271), 
            .CO(n26040));
    SB_CARRY add_563_11 (.CI(n24849), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n2629[9]), .CO(n24850));
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3392[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3392[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3392[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3392[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3392[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3392[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3392[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3392[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3392[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3392[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3392[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3392[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3392[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3392[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3392[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3392[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3392[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3392[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3392[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3392[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3392[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3416 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i28001_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4197), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4132), .O(n33677));
    defparam i28001_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_4662_6_lut (.I0(GND_net), .I1(n8296[3]), .I2(n390_adj_4272), 
            .I3(n26038), .O(n8279[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_6 (.CI(n26038), .I0(n8296[3]), .I1(n390_adj_4272), 
            .CO(n26039));
    SB_LUT4 add_4662_5_lut (.I0(GND_net), .I1(n8296[2]), .I2(n317_adj_4273), 
            .I3(n26037), .O(n8279[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_5 (.CI(n26037), .I0(n8296[2]), .I1(n317_adj_4273), 
            .CO(n26038));
    SB_LUT4 add_4662_4_lut (.I0(GND_net), .I1(n8296[1]), .I2(n244_adj_4274), 
            .I3(n26036), .O(n8279[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_4 (.CI(n26036), .I0(n8296[1]), .I1(n244_adj_4274), 
            .CO(n26037));
    SB_LUT4 add_4662_3_lut (.I0(GND_net), .I1(n8296[0]), .I2(n171_adj_4275), 
            .I3(n26035), .O(n8279[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_3 (.CI(n26035), .I0(n8296[0]), .I1(n171_adj_4275), 
            .CO(n26036));
    SB_LUT4 add_4662_2_lut (.I0(GND_net), .I1(n29_adj_4276), .I2(n98_adj_4277), 
            .I3(GND_net), .O(n8279[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4662_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4662_2 (.CI(GND_net), .I0(n29_adj_4276), .I1(n98_adj_4277), 
            .CO(n26035));
    SB_LUT4 add_4661_17_lut (.I0(GND_net), .I1(n8279[14]), .I2(GND_net), 
            .I3(n26034), .O(n8261[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4661_16_lut (.I0(GND_net), .I1(n8279[13]), .I2(n1117_adj_4278), 
            .I3(n26033), .O(n8261[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_16 (.CI(n26033), .I0(n8279[13]), .I1(n1117_adj_4278), 
            .CO(n26034));
    SB_LUT4 add_4661_15_lut (.I0(GND_net), .I1(n8279[12]), .I2(n1044_adj_4279), 
            .I3(n26032), .O(n8261[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_15 (.CI(n26032), .I0(n8279[12]), .I1(n1044_adj_4279), 
            .CO(n26033));
    SB_LUT4 add_4661_14_lut (.I0(GND_net), .I1(n8279[11]), .I2(n971_adj_4280), 
            .I3(n26031), .O(n8261[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_14 (.CI(n26031), .I0(n8279[11]), .I1(n971_adj_4280), 
            .CO(n26032));
    SB_LUT4 add_4661_13_lut (.I0(GND_net), .I1(n8279[10]), .I2(n898_adj_4281), 
            .I3(n26030), .O(n8261[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_13 (.CI(n26030), .I0(n8279[10]), .I1(n898_adj_4281), 
            .CO(n26031));
    SB_LUT4 add_4661_12_lut (.I0(GND_net), .I1(n8279[9]), .I2(n825_adj_4282), 
            .I3(n26029), .O(n8261[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_12 (.CI(n26029), .I0(n8279[9]), .I1(n825_adj_4282), 
            .CO(n26030));
    SB_LUT4 add_4661_11_lut (.I0(GND_net), .I1(n8279[8]), .I2(n752_adj_4283), 
            .I3(n26028), .O(n8261[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_11 (.CI(n26028), .I0(n8279[8]), .I1(n752_adj_4283), 
            .CO(n26029));
    SB_LUT4 add_4661_10_lut (.I0(GND_net), .I1(n8279[7]), .I2(n679_adj_4284), 
            .I3(n26027), .O(n8261[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_10 (.CI(n26027), .I0(n8279[7]), .I1(n679_adj_4284), 
            .CO(n26028));
    SB_LUT4 add_4661_9_lut (.I0(GND_net), .I1(n8279[6]), .I2(n606_adj_4285), 
            .I3(n26026), .O(n8261[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_9 (.CI(n26026), .I0(n8279[6]), .I1(n606_adj_4285), 
            .CO(n26027));
    SB_LUT4 add_4661_8_lut (.I0(GND_net), .I1(n8279[5]), .I2(n533_adj_4286), 
            .I3(n26025), .O(n8261[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_8 (.CI(n26025), .I0(n8279[5]), .I1(n533_adj_4286), 
            .CO(n26026));
    SB_LUT4 add_4661_7_lut (.I0(GND_net), .I1(n8279[4]), .I2(n460_adj_4287), 
            .I3(n26024), .O(n8261[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_7 (.CI(n26024), .I0(n8279[4]), .I1(n460_adj_4287), 
            .CO(n26025));
    SB_LUT4 add_4661_6_lut (.I0(GND_net), .I1(n8279[3]), .I2(n387_adj_4288), 
            .I3(n26023), .O(n8261[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_6 (.CI(n26023), .I0(n8279[3]), .I1(n387_adj_4288), 
            .CO(n26024));
    SB_LUT4 add_4661_5_lut (.I0(GND_net), .I1(n8279[2]), .I2(n314_adj_4289), 
            .I3(n26022), .O(n8261[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_5 (.CI(n26022), .I0(n8279[2]), .I1(n314_adj_4289), 
            .CO(n26023));
    SB_LUT4 add_4661_4_lut (.I0(GND_net), .I1(n8279[1]), .I2(n241_adj_4290), 
            .I3(n26021), .O(n8261[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4661_4 (.CI(n26021), .I0(n8279[1]), .I1(n241_adj_4290), 
            .CO(n26022));
    SB_LUT4 add_4661_3_lut (.I0(GND_net), .I1(n8279[0]), .I2(n168_adj_4291), 
            .I3(n26020), .O(n8261[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4338[16]), .I3(n25092), .O(n33_adj_4060)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4661_3 (.CI(n26020), .I0(n8279[0]), .I1(n168_adj_4291), 
            .CO(n26021));
    SB_LUT4 add_4661_2_lut (.I0(GND_net), .I1(n26_adj_4293), .I2(n95_adj_4294), 
            .I3(GND_net), .O(n8261[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4661_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n25092), .I0(GND_net), .I1(n1_adj_4338[16]), 
            .CO(n25093));
    SB_CARRY add_4661_2 (.CI(GND_net), .I0(n26_adj_4293), .I1(n95_adj_4294), 
            .CO(n26020));
    SB_LUT4 add_4660_18_lut (.I0(GND_net), .I1(n8261[15]), .I2(GND_net), 
            .I3(n26019), .O(n8242[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4660_17_lut (.I0(GND_net), .I1(n8261[14]), .I2(GND_net), 
            .I3(n26018), .O(n8242[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n2629[21]), .I3(n24861), .O(\PID_CONTROLLER.integral_23__N_3416 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_17 (.CI(n26018), .I0(n8261[14]), .I1(GND_net), .CO(n26019));
    SB_LUT4 add_4660_16_lut (.I0(GND_net), .I1(n8261[13]), .I2(n1114_adj_4295), 
            .I3(n26017), .O(n8242[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4338[15]), .I3(n25091), .O(n31_adj_4056)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4660_16 (.CI(n26017), .I0(n8261[13]), .I1(n1114_adj_4295), 
            .CO(n26018));
    SB_LUT4 add_4660_15_lut (.I0(GND_net), .I1(n8261[12]), .I2(n1041_adj_4297), 
            .I3(n26016), .O(n8242[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_15 (.CI(n26016), .I0(n8261[12]), .I1(n1041_adj_4297), 
            .CO(n26017));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n25091), .I0(GND_net), .I1(n1_adj_4338[15]), 
            .CO(n25092));
    SB_LUT4 add_4660_14_lut (.I0(GND_net), .I1(n8261[11]), .I2(n968_adj_4298), 
            .I3(n26015), .O(n8242[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_14 (.CI(n26015), .I0(n8261[11]), .I1(n968_adj_4298), 
            .CO(n26016));
    SB_LUT4 add_4660_13_lut (.I0(GND_net), .I1(n8261[10]), .I2(n895_adj_4299), 
            .I3(n26014), .O(n8242[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_13 (.CI(n26014), .I0(n8261[10]), .I1(n895_adj_4299), 
            .CO(n26015));
    SB_LUT4 add_4660_12_lut (.I0(GND_net), .I1(n8261[9]), .I2(n822_adj_4300), 
            .I3(n26013), .O(n8242[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_12 (.CI(n26013), .I0(n8261[9]), .I1(n822_adj_4300), 
            .CO(n26014));
    SB_LUT4 add_4660_11_lut (.I0(GND_net), .I1(n8261[8]), .I2(n749_adj_4301), 
            .I3(n26012), .O(n8242[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_11 (.CI(n26012), .I0(n8261[8]), .I1(n749_adj_4301), 
            .CO(n26013));
    SB_LUT4 add_4660_10_lut (.I0(GND_net), .I1(n8261[7]), .I2(n676_adj_4302), 
            .I3(n26011), .O(n8242[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4338[14]), .I3(n25090), .O(n29_adj_4057)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4660_10 (.CI(n26011), .I0(n8261[7]), .I1(n676_adj_4302), 
            .CO(n26012));
    SB_CARRY unary_minus_5_add_3_16 (.CI(n25090), .I0(GND_net), .I1(n1_adj_4338[14]), 
            .CO(n25091));
    SB_LUT4 add_4660_9_lut (.I0(GND_net), .I1(n8261[6]), .I2(n603_adj_4304), 
            .I3(n26010), .O(n8242[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_9 (.CI(n26010), .I0(n8261[6]), .I1(n603_adj_4304), 
            .CO(n26011));
    SB_LUT4 add_4660_8_lut (.I0(GND_net), .I1(n8261[5]), .I2(n530_adj_4305), 
            .I3(n26009), .O(n8242[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_8 (.CI(n26009), .I0(n8261[5]), .I1(n530_adj_4305), 
            .CO(n26010));
    SB_LUT4 add_4660_7_lut (.I0(GND_net), .I1(n8261[4]), .I2(n457_adj_4306), 
            .I3(n26008), .O(n8242[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_7 (.CI(n26008), .I0(n8261[4]), .I1(n457_adj_4306), 
            .CO(n26009));
    SB_LUT4 add_4660_6_lut (.I0(GND_net), .I1(n8261[3]), .I2(n384_adj_4307), 
            .I3(n26007), .O(n8242[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4338[13]), .I3(n25089), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4660_6 (.CI(n26007), .I0(n8261[3]), .I1(n384_adj_4307), 
            .CO(n26008));
    SB_LUT4 add_4660_5_lut (.I0(GND_net), .I1(n8261[2]), .I2(n311_adj_4309), 
            .I3(n26006), .O(n8242[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_5 (.CI(n26006), .I0(n8261[2]), .I1(n311_adj_4309), 
            .CO(n26007));
    SB_LUT4 add_4660_4_lut (.I0(GND_net), .I1(n8261[1]), .I2(n238_adj_4310), 
            .I3(n26005), .O(n8242[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_4 (.CI(n26005), .I0(n8261[1]), .I1(n238_adj_4310), 
            .CO(n26006));
    SB_LUT4 add_4660_3_lut (.I0(GND_net), .I1(n8261[0]), .I2(n165_adj_4311), 
            .I3(n26004), .O(n8242[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4660_3 (.CI(n26004), .I0(n8261[0]), .I1(n165_adj_4311), 
            .CO(n26005));
    SB_LUT4 add_4660_2_lut (.I0(GND_net), .I1(n23_adj_4312), .I2(n92_adj_4313), 
            .I3(GND_net), .O(n8242[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4660_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_23 (.CI(n24861), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n2629[21]), .CO(n24862));
    SB_CARRY add_4660_2 (.CI(GND_net), .I0(n23_adj_4312), .I1(n92_adj_4313), 
            .CO(n26004));
    SB_LUT4 add_4659_19_lut (.I0(GND_net), .I1(n8242[16]), .I2(GND_net), 
            .I3(n26003), .O(n8222[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_18_lut (.I0(GND_net), .I1(n8242[15]), .I2(GND_net), 
            .I3(n26002), .O(n8222[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_18 (.CI(n26002), .I0(n8242[15]), .I1(GND_net), .CO(n26003));
    SB_LUT4 add_4659_17_lut (.I0(GND_net), .I1(n8242[14]), .I2(GND_net), 
            .I3(n26001), .O(n8222[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_17 (.CI(n26001), .I0(n8242[14]), .I1(GND_net), .CO(n26002));
    SB_LUT4 add_4659_16_lut (.I0(GND_net), .I1(n8242[13]), .I2(n1111_adj_4314), 
            .I3(n26000), .O(n8222[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_16 (.CI(n26000), .I0(n8242[13]), .I1(n1111_adj_4314), 
            .CO(n26001));
    SB_LUT4 add_4659_15_lut (.I0(GND_net), .I1(n8242[12]), .I2(n1038_adj_4315), 
            .I3(n25999), .O(n8222[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_15 (.CI(n25999), .I0(n8242[12]), .I1(n1038_adj_4315), 
            .CO(n26000));
    SB_LUT4 add_4659_14_lut (.I0(GND_net), .I1(n8242[11]), .I2(n965_adj_4316), 
            .I3(n25998), .O(n8222[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_14 (.CI(n25998), .I0(n8242[11]), .I1(n965_adj_4316), 
            .CO(n25999));
    SB_LUT4 add_4659_13_lut (.I0(GND_net), .I1(n8242[10]), .I2(n892_adj_4317), 
            .I3(n25997), .O(n8222[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_13 (.CI(n25997), .I0(n8242[10]), .I1(n892_adj_4317), 
            .CO(n25998));
    SB_LUT4 add_4659_12_lut (.I0(GND_net), .I1(n8242[9]), .I2(n819_adj_4318), 
            .I3(n25996), .O(n8222[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_12 (.CI(n25996), .I0(n8242[9]), .I1(n819_adj_4318), 
            .CO(n25997));
    SB_CARRY unary_minus_5_add_3_15 (.CI(n25089), .I0(GND_net), .I1(n1_adj_4338[13]), 
            .CO(n25090));
    SB_LUT4 add_4659_11_lut (.I0(GND_net), .I1(n8242[8]), .I2(n746_adj_4319), 
            .I3(n25995), .O(n8222[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_11 (.CI(n25995), .I0(n8242[8]), .I1(n746_adj_4319), 
            .CO(n25996));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4338[12]), .I3(n25088), .O(n25_adj_4054)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4659_10_lut (.I0(GND_net), .I1(n8242[7]), .I2(n673_adj_4321), 
            .I3(n25994), .O(n8222[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_10 (.CI(n25994), .I0(n8242[7]), .I1(n673_adj_4321), 
            .CO(n25995));
    SB_LUT4 add_563_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n2629[20]), .I3(n24860), .O(\PID_CONTROLLER.integral_23__N_3416 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_9_lut (.I0(GND_net), .I1(n8242[6]), .I2(n600_adj_4322), 
            .I3(n25993), .O(n8222[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_9 (.CI(n25993), .I0(n8242[6]), .I1(n600_adj_4322), 
            .CO(n25994));
    SB_LUT4 add_4659_8_lut (.I0(GND_net), .I1(n8242[5]), .I2(n527_adj_4323), 
            .I3(n25992), .O(n8222[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n25088), .I0(GND_net), .I1(n1_adj_4338[12]), 
            .CO(n25089));
    SB_CARRY add_4659_8 (.CI(n25992), .I0(n8242[5]), .I1(n527_adj_4323), 
            .CO(n25993));
    SB_LUT4 add_4659_7_lut (.I0(GND_net), .I1(n8242[4]), .I2(n454_adj_4324), 
            .I3(n25991), .O(n8222[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_7 (.CI(n25991), .I0(n8242[4]), .I1(n454_adj_4324), 
            .CO(n25992));
    SB_LUT4 add_4659_6_lut (.I0(GND_net), .I1(n8242[3]), .I2(n381_adj_4325), 
            .I3(n25990), .O(n8222[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_6 (.CI(n25990), .I0(n8242[3]), .I1(n381_adj_4325), 
            .CO(n25991));
    SB_LUT4 add_4659_5_lut (.I0(GND_net), .I1(n8242[2]), .I2(n308_adj_4326), 
            .I3(n25989), .O(n8222[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_22 (.CI(n24860), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n2629[20]), .CO(n24861));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4338[11]), .I3(n25087), .O(n23_adj_4055)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n25087), .I0(GND_net), .I1(n1_adj_4338[11]), 
            .CO(n25088));
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4659_5 (.CI(n25989), .I0(n8242[2]), .I1(n308_adj_4326), 
            .CO(n25990));
    SB_LUT4 add_4659_4_lut (.I0(GND_net), .I1(n8242[1]), .I2(n235_adj_4329), 
            .I3(n25988), .O(n8222[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_4 (.CI(n25988), .I0(n8242[1]), .I1(n235_adj_4329), 
            .CO(n25989));
    SB_LUT4 add_4659_3_lut (.I0(GND_net), .I1(n8242[0]), .I2(n162_adj_4330), 
            .I3(n25987), .O(n8222[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_3 (.CI(n25987), .I0(n8242[0]), .I1(n162_adj_4330), 
            .CO(n25988));
    SB_LUT4 add_4659_2_lut (.I0(GND_net), .I1(n20_adj_4331), .I2(n89_adj_4332), 
            .I3(GND_net), .O(n8222[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_2 (.CI(GND_net), .I0(n20_adj_4331), .I1(n89_adj_4332), 
            .CO(n25987));
    SB_LUT4 add_4658_20_lut (.I0(GND_net), .I1(n8222[17]), .I2(GND_net), 
            .I3(n25986), .O(n8201[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4658_19_lut (.I0(GND_net), .I1(n8222[16]), .I2(GND_net), 
            .I3(n25985), .O(n8201[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_19 (.CI(n25985), .I0(n8222[16]), .I1(GND_net), .CO(n25986));
    SB_LUT4 add_4658_18_lut (.I0(GND_net), .I1(n8222[15]), .I2(GND_net), 
            .I3(n25984), .O(n8201[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_18 (.CI(n25984), .I0(n8222[15]), .I1(GND_net), .CO(n25985));
    SB_LUT4 add_4658_17_lut (.I0(GND_net), .I1(n8222[14]), .I2(GND_net), 
            .I3(n25983), .O(n8201[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_17 (.CI(n25983), .I0(n8222[14]), .I1(GND_net), .CO(n25984));
    SB_LUT4 add_4658_16_lut (.I0(GND_net), .I1(n8222[13]), .I2(n1108_adj_4333), 
            .I3(n25982), .O(n8201[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_16 (.CI(n25982), .I0(n8222[13]), .I1(n1108_adj_4333), 
            .CO(n25983));
    SB_LUT4 add_4658_15_lut (.I0(GND_net), .I1(n8222[12]), .I2(n1035_adj_4334), 
            .I3(n25981), .O(n8201[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n2629[19]), .I3(n24859), .O(\PID_CONTROLLER.integral_23__N_3416 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_15 (.CI(n25981), .I0(n8222[12]), .I1(n1035_adj_4334), 
            .CO(n25982));
    SB_LUT4 add_4658_14_lut (.I0(GND_net), .I1(n8222[11]), .I2(n962_adj_4335), 
            .I3(n25980), .O(n8201[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4338[10]), .I3(n25086), .O(n21_adj_4005)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n25086), .I0(GND_net), .I1(n1_adj_4338[10]), 
            .CO(n25087));
    SB_CARRY add_563_21 (.CI(n24859), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n2629[19]), .CO(n24860));
    SB_CARRY add_4658_14 (.CI(n25980), .I0(n8222[11]), .I1(n962_adj_4335), 
            .CO(n25981));
    SB_LUT4 add_4658_13_lut (.I0(GND_net), .I1(n8222[10]), .I2(n889_adj_4270), 
            .I3(n25979), .O(n8201[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_13 (.CI(n25979), .I0(n8222[10]), .I1(n889_adj_4270), 
            .CO(n25980));
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4658_12_lut (.I0(GND_net), .I1(n8222[9]), .I2(n816_adj_4268), 
            .I3(n25978), .O(n8201[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_12 (.CI(n25978), .I0(n8222[9]), .I1(n816_adj_4268), 
            .CO(n25979));
    SB_LUT4 add_4658_11_lut (.I0(GND_net), .I1(n8222[8]), .I2(n743_adj_4267), 
            .I3(n25977), .O(n8201[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_11 (.CI(n25977), .I0(n8222[8]), .I1(n743_adj_4267), 
            .CO(n25978));
    SB_LUT4 add_4658_10_lut (.I0(GND_net), .I1(n8222[7]), .I2(n670_adj_4265), 
            .I3(n25976), .O(n8201[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_10 (.CI(n25976), .I0(n8222[7]), .I1(n670_adj_4265), 
            .CO(n25977));
    SB_LUT4 add_4658_9_lut (.I0(GND_net), .I1(n8222[6]), .I2(n597_adj_4263), 
            .I3(n25975), .O(n8201[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_9 (.CI(n25975), .I0(n8222[6]), .I1(n597_adj_4263), 
            .CO(n25976));
    SB_LUT4 add_4658_8_lut (.I0(GND_net), .I1(n8222[5]), .I2(n524_adj_4258), 
            .I3(n25974), .O(n8201[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_8 (.CI(n25974), .I0(n8222[5]), .I1(n524_adj_4258), 
            .CO(n25975));
    SB_LUT4 add_4658_7_lut (.I0(GND_net), .I1(n8222[4]), .I2(n451_adj_4253), 
            .I3(n25973), .O(n8201[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_7 (.CI(n25973), .I0(n8222[4]), .I1(n451_adj_4253), 
            .CO(n25974));
    SB_LUT4 add_4658_6_lut (.I0(GND_net), .I1(n8222[3]), .I2(n378_adj_4214), 
            .I3(n25972), .O(n8201[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_6 (.CI(n25972), .I0(n8222[3]), .I1(n378_adj_4214), 
            .CO(n25973));
    SB_LUT4 add_4658_5_lut (.I0(GND_net), .I1(n8222[2]), .I2(n305_adj_4203), 
            .I3(n25971), .O(n8201[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_5 (.CI(n25971), .I0(n8222[2]), .I1(n305_adj_4203), 
            .CO(n25972));
    SB_LUT4 add_4658_4_lut (.I0(GND_net), .I1(n8222[1]), .I2(n232_adj_4195), 
            .I3(n25970), .O(n8201[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_4 (.CI(n25970), .I0(n8222[1]), .I1(n232_adj_4195), 
            .CO(n25971));
    SB_LUT4 add_4658_3_lut (.I0(GND_net), .I1(n8222[0]), .I2(n159_adj_4158), 
            .I3(n25969), .O(n8201[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_3 (.CI(n25969), .I0(n8222[0]), .I1(n159_adj_4158), 
            .CO(n25970));
    SB_LUT4 add_4658_2_lut (.I0(GND_net), .I1(n17_adj_4156), .I2(n86_adj_4155), 
            .I3(GND_net), .O(n8201[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4658_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4658_2 (.CI(GND_net), .I0(n17_adj_4156), .I1(n86_adj_4155), 
            .CO(n25969));
    SB_LUT4 add_4657_21_lut (.I0(GND_net), .I1(n8201[18]), .I2(GND_net), 
            .I3(n25968), .O(n8179[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4338[9]), .I3(n25085), .O(n19_adj_4006)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17472_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17472_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4334));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4657_20_lut (.I0(GND_net), .I1(n8201[17]), .I2(GND_net), 
            .I3(n25967), .O(n8179[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_20 (.CI(n25967), .I0(n8201[17]), .I1(GND_net), .CO(n25968));
    SB_LUT4 add_4657_19_lut (.I0(GND_net), .I1(n8201[16]), .I2(GND_net), 
            .I3(n25966), .O(n8179[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_19 (.CI(n25966), .I0(n8201[16]), .I1(GND_net), .CO(n25967));
    SB_LUT4 add_4657_18_lut (.I0(GND_net), .I1(n8201[15]), .I2(GND_net), 
            .I3(n25965), .O(n8179[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_18 (.CI(n25965), .I0(n8201[15]), .I1(GND_net), .CO(n25966));
    SB_LUT4 add_4657_17_lut (.I0(GND_net), .I1(n8201[14]), .I2(GND_net), 
            .I3(n25964), .O(n8179[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_17 (.CI(n25964), .I0(n8201[14]), .I1(GND_net), .CO(n25965));
    SB_LUT4 add_4657_16_lut (.I0(GND_net), .I1(n8201[13]), .I2(n1105_adj_4097), 
            .I3(n25963), .O(n8179[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_16 (.CI(n25963), .I0(n8201[13]), .I1(n1105_adj_4097), 
            .CO(n25964));
    SB_LUT4 add_4657_15_lut (.I0(GND_net), .I1(n8201[12]), .I2(n1032_adj_4096), 
            .I3(n25962), .O(n8179[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_15 (.CI(n25962), .I0(n8201[12]), .I1(n1032_adj_4096), 
            .CO(n25963));
    SB_LUT4 add_4657_14_lut (.I0(GND_net), .I1(n8201[11]), .I2(n959_adj_4095), 
            .I3(n25961), .O(n8179[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_14 (.CI(n25961), .I0(n8201[11]), .I1(n959_adj_4095), 
            .CO(n25962));
    SB_LUT4 add_4657_13_lut (.I0(GND_net), .I1(n8201[10]), .I2(n886_adj_4094), 
            .I3(n25960), .O(n8179[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_13 (.CI(n25960), .I0(n8201[10]), .I1(n886_adj_4094), 
            .CO(n25961));
    SB_LUT4 add_4657_12_lut (.I0(GND_net), .I1(n8201[9]), .I2(n813_adj_4093), 
            .I3(n25959), .O(n8179[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_12 (.CI(n25959), .I0(n8201[9]), .I1(n813_adj_4093), 
            .CO(n25960));
    SB_LUT4 add_4657_11_lut (.I0(GND_net), .I1(n8201[8]), .I2(n740_adj_4091), 
            .I3(n25958), .O(n8179[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_11 (.CI(n25958), .I0(n8201[8]), .I1(n740_adj_4091), 
            .CO(n25959));
    SB_LUT4 add_4657_10_lut (.I0(GND_net), .I1(n8201[7]), .I2(n667_adj_4090), 
            .I3(n25957), .O(n8179[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_10 (.CI(n25957), .I0(n8201[7]), .I1(n667_adj_4090), 
            .CO(n25958));
    SB_LUT4 add_4657_9_lut (.I0(GND_net), .I1(n8201[6]), .I2(n594_adj_4089), 
            .I3(n25956), .O(n8179[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_9 (.CI(n25956), .I0(n8201[6]), .I1(n594_adj_4089), 
            .CO(n25957));
    SB_LUT4 add_4657_8_lut (.I0(GND_net), .I1(n8201[5]), .I2(n521_adj_4087), 
            .I3(n25955), .O(n8179[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_8 (.CI(n25955), .I0(n8201[5]), .I1(n521_adj_4087), 
            .CO(n25956));
    SB_LUT4 add_4657_7_lut (.I0(GND_net), .I1(n8201[4]), .I2(n448_adj_4086), 
            .I3(n25954), .O(n8179[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_7 (.CI(n25954), .I0(n8201[4]), .I1(n448_adj_4086), 
            .CO(n25955));
    SB_LUT4 add_4657_6_lut (.I0(GND_net), .I1(n8201[3]), .I2(n375_adj_4085), 
            .I3(n25953), .O(n8179[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_6 (.CI(n25953), .I0(n8201[3]), .I1(n375_adj_4085), 
            .CO(n25954));
    SB_LUT4 add_4657_5_lut (.I0(GND_net), .I1(n8201[2]), .I2(n302_adj_4084), 
            .I3(n25952), .O(n8179[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_5 (.CI(n25952), .I0(n8201[2]), .I1(n302_adj_4084), 
            .CO(n25953));
    SB_LUT4 add_4657_4_lut (.I0(GND_net), .I1(n8201[1]), .I2(n229_adj_4083), 
            .I3(n25951), .O(n8179[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_4 (.CI(n25951), .I0(n8201[1]), .I1(n229_adj_4083), 
            .CO(n25952));
    SB_LUT4 add_4657_3_lut (.I0(GND_net), .I1(n8201[0]), .I2(n156_adj_4082), 
            .I3(n25950), .O(n8179[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_3 (.CI(n25950), .I0(n8201[0]), .I1(n156_adj_4082), 
            .CO(n25951));
    SB_LUT4 add_4657_2_lut (.I0(GND_net), .I1(n14_adj_4081), .I2(n83_adj_4079), 
            .I3(GND_net), .O(n8179[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4657_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4657_2 (.CI(GND_net), .I0(n14_adj_4081), .I1(n83_adj_4079), 
            .CO(n25950));
    SB_LUT4 add_4656_22_lut (.I0(GND_net), .I1(n8179[19]), .I2(GND_net), 
            .I3(n25949), .O(n8156[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4656_21_lut (.I0(GND_net), .I1(n8179[18]), .I2(GND_net), 
            .I3(n25948), .O(n8156[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_21 (.CI(n25948), .I0(n8179[18]), .I1(GND_net), .CO(n25949));
    SB_LUT4 add_4656_20_lut (.I0(GND_net), .I1(n8179[17]), .I2(GND_net), 
            .I3(n25947), .O(n8156[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_20 (.CI(n25947), .I0(n8179[17]), .I1(GND_net), .CO(n25948));
    SB_LUT4 add_4656_19_lut (.I0(GND_net), .I1(n8179[16]), .I2(GND_net), 
            .I3(n25946), .O(n8156[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_19 (.CI(n25946), .I0(n8179[16]), .I1(GND_net), .CO(n25947));
    SB_LUT4 add_4656_18_lut (.I0(GND_net), .I1(n8179[15]), .I2(GND_net), 
            .I3(n25945), .O(n8156[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_18 (.CI(n25945), .I0(n8179[15]), .I1(GND_net), .CO(n25946));
    SB_LUT4 add_4656_17_lut (.I0(GND_net), .I1(n8179[14]), .I2(GND_net), 
            .I3(n25944), .O(n8156[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_17 (.CI(n25944), .I0(n8179[14]), .I1(GND_net), .CO(n25945));
    SB_LUT4 add_4656_16_lut (.I0(GND_net), .I1(n8179[13]), .I2(n1102_adj_4078), 
            .I3(n25943), .O(n8156[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_16 (.CI(n25943), .I0(n8179[13]), .I1(n1102_adj_4078), 
            .CO(n25944));
    SB_LUT4 add_4656_15_lut (.I0(GND_net), .I1(n8179[12]), .I2(n1029_adj_4075), 
            .I3(n25942), .O(n8156[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_15 (.CI(n25942), .I0(n8179[12]), .I1(n1029_adj_4075), 
            .CO(n25943));
    SB_LUT4 add_4656_14_lut (.I0(GND_net), .I1(n8179[11]), .I2(n956_adj_4073), 
            .I3(n25941), .O(n8156[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_14 (.CI(n25941), .I0(n8179[11]), .I1(n956_adj_4073), 
            .CO(n25942));
    SB_LUT4 add_4656_13_lut (.I0(GND_net), .I1(n8179[10]), .I2(n883_adj_4072), 
            .I3(n25940), .O(n8156[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_13 (.CI(n25940), .I0(n8179[10]), .I1(n883_adj_4072), 
            .CO(n25941));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n25085), .I0(GND_net), .I1(n1_adj_4338[9]), 
            .CO(n25086));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4338[8]), .I3(n25084), .O(n17_adj_4007)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4656_12_lut (.I0(GND_net), .I1(n8179[9]), .I2(n810_adj_4049), 
            .I3(n25939), .O(n8156[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_12 (.CI(n25939), .I0(n8179[9]), .I1(n810_adj_4049), 
            .CO(n25940));
    SB_LUT4 add_4656_11_lut (.I0(GND_net), .I1(n8179[8]), .I2(n737_adj_4048), 
            .I3(n25938), .O(n8156[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_11 (.CI(n25938), .I0(n8179[8]), .I1(n737_adj_4048), 
            .CO(n25939));
    SB_LUT4 add_4656_10_lut (.I0(GND_net), .I1(n8179[7]), .I2(n664_adj_4047), 
            .I3(n25937), .O(n8156[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_10 (.CI(n25937), .I0(n8179[7]), .I1(n664_adj_4047), 
            .CO(n25938));
    SB_LUT4 add_4656_9_lut (.I0(GND_net), .I1(n8179[6]), .I2(n591_adj_4045), 
            .I3(n25936), .O(n8156[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_9 (.CI(n25936), .I0(n8179[6]), .I1(n591_adj_4045), 
            .CO(n25937));
    SB_LUT4 add_4656_8_lut (.I0(GND_net), .I1(n8179[5]), .I2(n518_adj_4044), 
            .I3(n25935), .O(n8156[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_8 (.CI(n25935), .I0(n8179[5]), .I1(n518_adj_4044), 
            .CO(n25936));
    SB_LUT4 add_4656_7_lut (.I0(GND_net), .I1(n8179[4]), .I2(n445_adj_4043), 
            .I3(n25934), .O(n8156[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_7 (.CI(n25934), .I0(n8179[4]), .I1(n445_adj_4043), 
            .CO(n25935));
    SB_LUT4 add_4656_6_lut (.I0(GND_net), .I1(n8179[3]), .I2(n372_adj_4042), 
            .I3(n25933), .O(n8156[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_6 (.CI(n25933), .I0(n8179[3]), .I1(n372_adj_4042), 
            .CO(n25934));
    SB_LUT4 add_4656_5_lut (.I0(GND_net), .I1(n8179[2]), .I2(n299_adj_4041), 
            .I3(n25932), .O(n8156[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_5 (.CI(n25932), .I0(n8179[2]), .I1(n299_adj_4041), 
            .CO(n25933));
    SB_LUT4 add_4656_4_lut (.I0(GND_net), .I1(n8179[1]), .I2(n226_adj_4040), 
            .I3(n25931), .O(n8156[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_4 (.CI(n25931), .I0(n8179[1]), .I1(n226_adj_4040), 
            .CO(n25932));
    SB_LUT4 add_4656_3_lut (.I0(GND_net), .I1(n8179[0]), .I2(n153_adj_4039), 
            .I3(n25930), .O(n8156[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_3 (.CI(n25930), .I0(n8179[0]), .I1(n153_adj_4039), 
            .CO(n25931));
    SB_LUT4 add_4656_2_lut (.I0(GND_net), .I1(n11_adj_4038), .I2(n80_adj_4037), 
            .I3(GND_net), .O(n8156[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_2 (.CI(GND_net), .I0(n11_adj_4038), .I1(n80_adj_4037), 
            .CO(n25930));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n8132[21]), .I2(GND_net), 
            .I3(n25929), .O(n6838[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n8132[20]), .I2(GND_net), 
            .I3(n25928), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n25928), .I0(n8132[20]), .I1(GND_net), 
            .CO(n25929));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n8132[19]), .I2(GND_net), 
            .I3(n25927), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n25927), .I0(n8132[19]), .I1(GND_net), 
            .CO(n25928));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n8132[18]), .I2(GND_net), 
            .I3(n25926), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n25926), .I0(n8132[18]), .I1(GND_net), 
            .CO(n25927));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n8132[17]), .I2(GND_net), 
            .I3(n25925), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n25925), .I0(n8132[17]), .I1(GND_net), 
            .CO(n25926));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n8132[16]), .I2(GND_net), 
            .I3(n25924), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n25924), .I0(n8132[16]), .I1(GND_net), 
            .CO(n25925));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n8132[15]), .I2(GND_net), 
            .I3(n25923), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n25923), .I0(n8132[15]), .I1(GND_net), 
            .CO(n25924));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n8132[14]), .I2(GND_net), 
            .I3(n25922), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n25922), .I0(n8132[14]), .I1(GND_net), 
            .CO(n25923));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n8132[13]), .I2(n1096_adj_4034), 
            .I3(n25921), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n25921), .I0(n8132[13]), .I1(n1096_adj_4034), 
            .CO(n25922));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n8132[12]), .I2(n1023_adj_4033), 
            .I3(n25920), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n25920), .I0(n8132[12]), .I1(n1023_adj_4033), 
            .CO(n25921));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n8132[11]), .I2(n950_adj_4032), 
            .I3(n25919), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n25919), .I0(n8132[11]), .I1(n950_adj_4032), 
            .CO(n25920));
    SB_CARRY unary_minus_5_add_3_10 (.CI(n25084), .I0(GND_net), .I1(n1_adj_4338[8]), 
            .CO(n25085));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n8132[10]), .I2(n877_adj_4031), 
            .I3(n25918), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4338[7]), .I3(n25083), .O(n15_adj_3948)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_563_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n2629[18]), .I3(n24858), .O(\PID_CONTROLLER.integral_23__N_3416 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n25918), .I0(n8132[10]), .I1(n877_adj_4031), 
            .CO(n25919));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n25083), .I0(GND_net), .I1(n1_adj_4338[7]), 
            .CO(n25084));
    SB_CARRY add_563_20 (.CI(n24858), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n2629[18]), .CO(n24859));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4338[6]), .I3(n25082), .O(n13_adj_3949)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n6838[0]), .I2(n6842[0]), 
            .I3(n24924), .O(duty_23__N_3516[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n25082), .I0(GND_net), .I1(n1_adj_4338[6]), 
            .CO(n25083));
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4333));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4331));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4330));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n8132[9]), .I2(n804_adj_4028), 
            .I3(n25917), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n25917), .I0(n8132[9]), .I1(n804_adj_4028), 
            .CO(n25918));
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_563_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n2629[17]), .I3(n24857), .O(\PID_CONTROLLER.integral_23__N_3416 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4338[5]), .I3(n25081), .O(n11_adj_3950)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n8132[8]), .I2(n731_adj_4027), 
            .I3(n25916), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n25916), .I0(n8132[8]), .I1(n731_adj_4027), 
            .CO(n25917));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n25081), .I0(GND_net), .I1(n1_adj_4338[5]), 
            .CO(n25082));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4338[4]), .I3(n25080), .O(n9_adj_4008)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n8132[7]), .I2(n658_adj_4025), 
            .I3(n25915), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n25915), .I0(n8132[7]), .I1(n658_adj_4025), 
            .CO(n25916));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n8132[6]), .I2(n585_adj_4024), 
            .I3(n25914), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n24923), .O(duty_23__N_3516[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n25914), .I0(n8132[6]), .I1(n585_adj_4024), 
            .CO(n25915));
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_563_19 (.CI(n24857), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n2629[17]), .CO(n24858));
    SB_CARRY unary_minus_5_add_3_6 (.CI(n25080), .I0(GND_net), .I1(n1_adj_4338[4]), 
            .CO(n25081));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4338[3]), .I3(n25079), .O(n7_adj_4052)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n25079), .I0(GND_net), .I1(n1_adj_4338[3]), 
            .CO(n25080));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n8132[5]), .I2(n512_adj_4022), 
            .I3(n25913), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4338[2]), .I3(n25078), .O(n5_adj_4053)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_10_add_1225_8 (.CI(n25913), .I0(n8132[5]), .I1(n512_adj_4022), 
            .CO(n25914));
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4325));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20613_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [18]), 
            .I2(n4_adj_4336), .I3(n8708[1]), .O(n6_adj_4050));   // verilog/motorControl.v(34[25:36])
    defparam i20613_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n8132[4]), .I2(n439_adj_4020), 
            .I3(n25912), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4324));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_7 (.CI(n25912), .I0(n8132[4]), .I1(n439_adj_4020), 
            .CO(n25913));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n8132[3]), .I2(n366_adj_4019), 
            .I3(n25911), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n25078), .I0(GND_net), .I1(n1_adj_4338[2]), 
            .CO(n25079));
    SB_CARRY mult_10_add_1225_6 (.CI(n25911), .I0(n8132[3]), .I1(n366_adj_4019), 
            .CO(n25912));
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [18]), 
            .I2(n8708[1]), .I3(n4_adj_4336), .O(n8701[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n8132[2]), .I2(n293_adj_4018), 
            .I3(n25910), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n25910), .I0(n8132[2]), .I1(n293_adj_4018), 
            .CO(n25911));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n8132[1]), .I2(n220_adj_4017), 
            .I3(n25909), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n25909), .I0(n8132[1]), .I1(n220_adj_4017), 
            .CO(n25910));
    SB_LUT4 i2_3_lut_4_lut_adj_1482 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [18]), 
            .I2(n8708[0]), .I3(n24680), .O(n8701[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1482.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n8132[0]), .I2(n147_adj_4016), 
            .I3(n25908), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n25908), .I0(n8132[0]), .I1(n147_adj_4016), 
            .CO(n25909));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4015), .I2(n74_adj_4014), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4338[1]), .I3(n25077), .O(n3_adj_4115)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4322));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17473_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17473_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n25077), .I0(GND_net), .I1(n1_adj_4338[1]), 
            .CO(n25078));
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4321));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4319));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4318));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4317));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4316));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20605_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [18]), 
            .I2(n24680), .I3(n8708[0]), .O(n4_adj_4336));   // verilog/motorControl.v(34[25:36])
    defparam i20605_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4315));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4015), .I1(n74_adj_4014), 
            .CO(n25908));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4338[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3467 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_24 (.CI(n24923), .I0(n106[22]), .I1(n155[22]), .CO(n24924));
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4338[0]), 
            .CO(n25077));
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4313));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4655_23_lut (.I0(GND_net), .I1(n8156[20]), .I2(GND_net), 
            .I3(n25901), .O(n8132[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4655_22_lut (.I0(GND_net), .I1(n8156[19]), .I2(GND_net), 
            .I3(n25900), .O(n8132[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_22 (.CI(n25900), .I0(n8156[19]), .I1(GND_net), .CO(n25901));
    SB_LUT4 add_4655_21_lut (.I0(GND_net), .I1(n8156[18]), .I2(GND_net), 
            .I3(n25899), .O(n8132[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_21 (.CI(n25899), .I0(n8156[18]), .I1(GND_net), .CO(n25900));
    SB_LUT4 add_4655_20_lut (.I0(GND_net), .I1(n8156[17]), .I2(GND_net), 
            .I3(n25898), .O(n8132[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_20 (.CI(n25898), .I0(n8156[17]), .I1(GND_net), .CO(n25899));
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4312));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4655_19_lut (.I0(GND_net), .I1(n8156[16]), .I2(GND_net), 
            .I3(n25897), .O(n8132[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_19 (.CI(n25897), .I0(n8156[16]), .I1(GND_net), .CO(n25898));
    SB_LUT4 add_4655_18_lut (.I0(GND_net), .I1(n8156[15]), .I2(GND_net), 
            .I3(n25896), .O(n8132[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4655_18 (.CI(n25896), .I0(n8156[15]), .I1(GND_net), .CO(n25897));
    SB_LUT4 add_4655_17_lut (.I0(GND_net), .I1(n8156[14]), .I2(GND_net), 
            .I3(n25895), .O(n8132[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20594_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3416 [18]), .I3(\Ki[1] ), 
            .O(n24680));   // verilog/motorControl.v(34[25:36])
    defparam i20594_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_4655_17 (.CI(n25895), .I0(n8156[14]), .I1(GND_net), .CO(n25896));
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4310));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20592_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3416 [18]), .I3(\Ki[1] ), 
            .O(n8701[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20592_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_4655_16_lut (.I0(GND_net), .I1(n8156[13]), .I2(n1099_adj_3945), 
            .I3(n25894), .O(n8132[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_16 (.CI(n25894), .I0(n8156[13]), .I1(n1099_adj_3945), 
            .CO(n25895));
    SB_LUT4 add_4655_15_lut (.I0(GND_net), .I1(n8156[12]), .I2(n1026_adj_3944), 
            .I3(n25893), .O(n8132[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4309));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4655_15 (.CI(n25893), .I0(n8156[12]), .I1(n1026_adj_3944), 
            .CO(n25894));
    SB_LUT4 add_4655_14_lut (.I0(GND_net), .I1(n8156[11]), .I2(n953_adj_3943), 
            .I3(n25892), .O(n8132[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_14 (.CI(n25892), .I0(n8156[11]), .I1(n953_adj_3943), 
            .CO(n25893));
    SB_LUT4 add_4655_13_lut (.I0(GND_net), .I1(n8156[10]), .I2(n880_adj_3942), 
            .I3(n25891), .O(n8132[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_13 (.CI(n25891), .I0(n8156[10]), .I1(n880_adj_3942), 
            .CO(n25892));
    SB_LUT4 add_4655_12_lut (.I0(GND_net), .I1(n8156[9]), .I2(n807_adj_3941), 
            .I3(n25890), .O(n8132[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_12 (.CI(n25890), .I0(n8156[9]), .I1(n807_adj_3941), 
            .CO(n25891));
    SB_LUT4 add_4655_11_lut (.I0(GND_net), .I1(n8156[8]), .I2(n734_adj_3940), 
            .I3(n25889), .O(n8132[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_11 (.CI(n25889), .I0(n8156[8]), .I1(n734_adj_3940), 
            .CO(n25890));
    SB_LUT4 add_4655_10_lut (.I0(GND_net), .I1(n8156[7]), .I2(n661_adj_3938), 
            .I3(n25888), .O(n8132[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4655_10 (.CI(n25888), .I0(n8156[7]), .I1(n661_adj_3938), 
            .CO(n25889));
    SB_LUT4 add_4655_9_lut (.I0(GND_net), .I1(n8156[6]), .I2(n588_adj_3936), 
            .I3(n25887), .O(n8132[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_9 (.CI(n25887), .I0(n8156[6]), .I1(n588_adj_3936), 
            .CO(n25888));
    SB_LUT4 add_4655_8_lut (.I0(GND_net), .I1(n8156[5]), .I2(n515_adj_3935), 
            .I3(n25886), .O(n8132[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_8 (.CI(n25886), .I0(n8156[5]), .I1(n515_adj_3935), 
            .CO(n25887));
    SB_LUT4 add_4655_7_lut (.I0(GND_net), .I1(n8156[4]), .I2(n442_adj_3932), 
            .I3(n25885), .O(n8132[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4307));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4655_7 (.CI(n25885), .I0(n8156[4]), .I1(n442_adj_3932), 
            .CO(n25886));
    SB_LUT4 add_4655_6_lut (.I0(GND_net), .I1(n8156[3]), .I2(n369_adj_3929), 
            .I3(n25884), .O(n8132[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4306));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4655_6 (.CI(n25884), .I0(n8156[3]), .I1(n369_adj_3929), 
            .CO(n25885));
    SB_LUT4 add_4655_5_lut (.I0(GND_net), .I1(n8156[2]), .I2(n296_adj_3928), 
            .I3(n25883), .O(n8132[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_5 (.CI(n25883), .I0(n8156[2]), .I1(n296_adj_3928), 
            .CO(n25884));
    SB_LUT4 add_4655_4_lut (.I0(GND_net), .I1(n8156[1]), .I2(n223_adj_3925), 
            .I3(n25882), .O(n8132[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_4 (.CI(n25882), .I0(n8156[1]), .I1(n223_adj_3925), 
            .CO(n25883));
    SB_LUT4 add_4655_3_lut (.I0(GND_net), .I1(n8156[0]), .I2(n150_adj_3924), 
            .I3(n25881), .O(n8132[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_3 (.CI(n25881), .I0(n8156[0]), .I1(n150_adj_3924), 
            .CO(n25882));
    SB_LUT4 add_4655_2_lut (.I0(GND_net), .I1(n8_adj_3922), .I2(n77_adj_3921), 
            .I3(GND_net), .O(n8132[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4655_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4655_2 (.CI(GND_net), .I0(n8_adj_3922), .I1(n77_adj_3921), 
            .CO(n25881));
    SB_LUT4 i20675_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [20]), 
            .I2(n24757), .I3(n8719[0]), .O(n4_adj_4069));   // verilog/motorControl.v(34[25:36])
    defparam i20675_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n24922), .O(duty_23__N_3516[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1483 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [20]), 
            .I2(n8719[0]), .I3(n24757), .O(n8714[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1483.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1484 (.I0(n62), .I1(n131), .I2(n8714[0]), 
            .I3(n204_adj_4051), .O(n8708[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1484.LUT_INIT = 16'h8778;
    SB_LUT4 i20644_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204_adj_4051), 
            .I3(n8714[0]), .O(n4_adj_4062));   // verilog/motorControl.v(34[25:36])
    defparam i20644_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i20662_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3416 [20]), .I3(\Ki[1] ), 
            .O(n8714[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20662_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_563_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n2629[16]), .I3(n24856), .O(\PID_CONTROLLER.integral_23__N_3416 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4304));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_23 (.CI(n24922), .I0(n106[21]), .I1(n155[21]), .CO(n24923));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n24921), .O(duty_23__N_3516[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20664_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3416 [20]), .I3(\Ki[1] ), 
            .O(n24757));   // verilog/motorControl.v(34[25:36])
    defparam i20664_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_22 (.CI(n24921), .I0(n106[20]), .I1(n155[20]), .CO(n24922));
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n24920), .O(duty_23__N_3516[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4301));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4300));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_21 (.CI(n24920), .I0(n106[19]), .I1(n155[19]), .CO(n24921));
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4298));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n24919), .O(duty_23__N_3516[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_18 (.CI(n24856), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n2629[16]), .CO(n24857));
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4297));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_20 (.CI(n24919), .I0(n106[18]), .I1(n155[18]), .CO(n24920));
    SB_LUT4 add_563_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n2629[15]), .I3(n24855), .O(\PID_CONTROLLER.integral_23__N_3416 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4114));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4295));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17474_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17474_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4294));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4291));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4290));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n24918), .O(duty_23__N_3516[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4289));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4288));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4287));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4286));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4285));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4284));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4283));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4282));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4281));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4280));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4279));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4278));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4277));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4276));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4275));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4274));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4273));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4272));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3516[23]), .I1(n257[23]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3491[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3516[22]), .I1(n257[22]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3491[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3516[21]), .I1(n257[21]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3491[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3516[20]), .I1(n257[20]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3491[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3516[19]), .I1(n257[19]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3491[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3516[18]), .I1(n257[18]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3491[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3516[17]), .I1(n257[17]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3491[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3516[16]), .I1(n257[16]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3491[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3516[15]), .I1(n257[15]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3491[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(\duty_23__N_3516[14] ), .I1(n257[14]), 
            .I2(n256), .I3(GND_net), .O(duty_23__N_3491[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3491[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3516[13]), .I1(n257[13]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3491[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3516[12]), .I1(n257[12]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3491[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3516[11]), .I1(n257[11]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3491[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3516[10]), .I1(n257[10]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3491[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3516[9]), .I1(n257[9]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3491[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3516[8]), .I1(n257[8]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3491[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3516[7]), .I1(n257[7]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3491[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3516[6]), .I1(n257[6]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3491[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3516[5]), .I1(n257[5]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3491[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3516[4]), .I1(n257[4]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3491[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3516[3]), .I1(n257[3]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3491[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4271));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4269));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4266));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17475_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4264));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4262));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3516[2]), .I1(n257[2]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3491[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3491[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3392[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27622_3_lut_4_lut (.I0(duty_23__N_3516[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3516[2]), .O(n33296));   // verilog/motorControl.v(38[19:35])
    defparam i27622_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4261));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4259));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17476_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17476_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4257));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4256));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4255));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4252));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4251));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3516[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_3998));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4249));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4248));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4247));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4246));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4245));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4244));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4243));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4241));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4240));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4239));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4237));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4236));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4233));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4231));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4230));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4229));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4228));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4227));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4226));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4225));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27657_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3516[3]), 
            .I2(PWMLimit[2]), .I3(duty_23__N_3516[2]), .O(n33331));   // verilog/motorControl.v(36[10:25])
    defparam i27657_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_831_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3516[3]), 
            .I2(duty_23__N_3516[2]), .I3(GND_net), .O(n6_adj_3965));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4224));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4222));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4221));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4219));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4218));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4217));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4216));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4215));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4213));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4212));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4211));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4210));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4209));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4132));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4208));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4207));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4061));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4197));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4206));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4205));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4204));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4202));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4201));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4200));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4199));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4198));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4196));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4194));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4193));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4192));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4191));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4188));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4187));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4186));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4185));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4184));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4182));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4181));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4338[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4179));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4178));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4177));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4176));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20553_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n24625), 
            .I3(n8422[0]), .O(n4_adj_3917));   // verilog/motorControl.v(34[16:22])
    defparam i20553_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i20631_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3416 [19]), 
            .O(n8708[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20631_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4174));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20491_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4128), 
            .I3(n8411[1]), .O(n6_adj_3914));   // verilog/motorControl.v(34[16:22])
    defparam i20491_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4173));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27587_2_lut_4_lut (.I0(duty_23__N_3516[21]), .I1(n257[21]), 
            .I2(duty_23__N_3516[9]), .I3(n257[9]), .O(n33261));
    defparam i27587_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4172));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4171));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27598_2_lut_4_lut (.I0(duty_23__N_3516[16]), .I1(n257[16]), 
            .I2(duty_23__N_3516[7]), .I3(n257[7]), .O(n33272));
    defparam i27598_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i2_3_lut_4_lut_adj_1485 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n8411[1]), 
            .I3(n4_adj_4128), .O(n8404[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1485.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4170));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27625_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3516[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3516[9]), .O(n33299));
    defparam i27625_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4169));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4168));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4167));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4166));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27635_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3516[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3516[7]), .O(n33309));
    defparam i27635_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3416 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4160));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4154));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4337[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4151));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4150));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4149));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4148));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4147));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4146));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4145));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4144));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4143));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4142));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4141));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4140));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17469_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3464 ), 
            .I2(GND_net), .I3(GND_net), .O(n2629[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4139));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4138));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4137));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4136));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1486 (.I0(n6_adj_3914), .I1(\Kp[4] ), .I2(n8411[2]), 
            .I3(n1[18]), .O(n8404[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1486.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_4134));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4133));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_out_frame[23] , \data_out_frame[24] , GND_net, \data_out_frame[25] , 
            \data_out_frame[20] , \data_out_frame[18] , \data_out_frame[17] , 
            \data_out_frame[15] , setpoint, clk32MHz, \data_out_frame[5] , 
            \data_out_frame[11] , \data_out_frame[8] , \data_out_frame[7] , 
            \data_out_frame[14] , \data_out_frame[16] , \data_out_frame[19] , 
            \data_in_frame[3] , \data_out_frame[13] , \data_out_frame[6] , 
            \data_out_frame[10] , \data_out_frame[9] , \data_out_frame[12] , 
            n63, n771, n63_adj_3, \FRAME_MATCHER.i_31__N_2364 , n29497, 
            \FRAME_MATCHER.state[0] , \data_in_frame[1] , \data_in_frame[2] , 
            n12869, n2329, n4452, \data_in[0] , \data_in[2] , \data_in[3] , 
            \data_in[1] , \FRAME_MATCHER.i_31__N_2370 , PWMLimit, \duty_23__N_3516[14] , 
            n29, rx_data, \data_in_frame[13] , \data_in_frame[18] , 
            \FRAME_MATCHER.state[3] , tx_active, \FRAME_MATCHER.state[2] , 
            rx_data_ready, n16911, \data_in_frame[21] , n16910, n16909, 
            \data_in_frame[4] , \data_in_frame[7] , \data_in_frame[6] , 
            \data_in_frame[8] , n4218, n16908, n16907, \data_in_frame[9] , 
            \data_in_frame[9][5] , \data_in_frame[9][4] , \data_in_frame[9][3] , 
            \data_in_frame[9][2] , \data_in_frame[9][1] , \data_in_frame[9][0] , 
            n16906, n78, n16905, n16904, n16903, control_mode, n16902, 
            \data_in_frame[10] , \data_in_frame[5] , n16901, \data_in_frame[15] , 
            \data_in_frame[11] , \data_in_frame[12] , \data_in_frame[14] , 
            n16900, n16899, n12944, \data_in_frame[10][1] , n2, DE_c, 
            n8868, n16898, n16897, n16896, n16894, n16893, n16892, 
            n16891, n16890, n16889, n16888, n16887, n16886, n16885, 
            n16884, n16882, n16881, n16880, n16879, n16878, n16877, 
            n16876, n16875, n16874, n35073, n28937, n16867, VCC_net, 
            n17373, IntegralLimit, n17372, n17371, n17370, n17369, 
            n17368, n17367, n17335, n17334, n17333, n17332, n17331, 
            n17330, n17329, n17328, n17327, n17326, n17325, n17324, 
            n17323, n17322, n17321, n17320, n17314, n17313, n17312, 
            n17311, n17310, n17309, n17308, n17307, n17306, n17305, 
            n17304, n17303, n17302, n17301, n17300, n17299, n17298, 
            n17297, n17296, n17295, n17294, n17293, n17292, n17291, 
            n17290, n17289, n17288, n17287, n17286, n17285, n17284, 
            n17283, \Kp[1] , n17282, \Kp[2] , n17281, \Kp[3] , n17280, 
            \Kp[4] , n17279, \Kp[5] , n17278, \Kp[6] , n17277, \Kp[7] , 
            n17276, \Kp[8] , n17275, \Kp[9] , n17274, \Kp[10] , 
            n17273, \Kp[11] , n17272, \Kp[12] , n17271, \Kp[13] , 
            n17270, \Kp[14] , n17269, \Kp[15] , n17268, \Ki[1] , 
            n17267, \Ki[2] , n17266, \Ki[3] , n17265, \Ki[4] , n17264, 
            \Ki[5] , n17263, \Ki[6] , n17262, \Ki[7] , n17261, \Ki[8] , 
            n17260, \Ki[9] , n17259, \Ki[10] , n17258, \Ki[11] , 
            n17257, \Ki[12] , n17256, \Ki[13] , n17255, \Ki[14] , 
            n17254, \Ki[15] , n17253, n17252, n17251, n17250, n17249, 
            n17248, n17247, n17246, n17245, n17244, n17243, n17242, 
            n17241, n17240, n17239, n17238, n17237, n17236, n17235, 
            n17234, n17233, n17232, n4216, n122, n5, n35368, n17231, 
            n17230, n17229, n17228, n17227, n17226, n17225, n17224, 
            n17223, n17222, n17221, n17220, n17219, n17218, n17217, 
            n17216, n17215, n17214, n17213, n17212, n17211, n17210, 
            n17209, n17208, n17207, n17206, n17205, n17204, n17203, 
            n17202, n17201, n17200, n17199, n17198, n17197, n17196, 
            n17195, n17194, n17193, n17192, n17191, n17190, n17189, 
            n17188, n17187, n17186, n17185, n17184, n17183, n17182, 
            n17181, n17180, n17179, n17178, n17177, n17176, n17175, 
            n17174, n17173, n17172, n17171, n17170, n17169, n17168, 
            n17167, n17166, n17165, n17164, n17163, n17162, n17161, 
            n17160, n17159, n17158, n17157, n17156, n17155, n17154, 
            n17153, n17152, n17151, n17150, n17149, n17148, n17147, 
            n17146, n17145, n17144, n17143, n17142, n17141, n17140, 
            n17139, n17138, n17137, n17136, n17135, n17134, n17133, 
            n17132, n17131, n17130, n17129, n17128, n17127, n17126, 
            n17125, n17124, n17123, n17122, n17121, n17120, n17119, 
            n17118, n17117, n17116, n29535, n17115, n17114, n17113, 
            n17112, n17111, LED_c, n17110, n29532, n17109, n17108, 
            n17107, n17106, n17105, n17104, n17103, n17102, n17101, 
            neopxl_color, n17100, n17099, n17098, n17097, n17096, 
            n17095, n17094, n17093, n17092, n17091, n17090, n17089, 
            n17088, n17087, n17086, n17085, n17084, n17083, n17082, 
            n17081, n17080, n17079, n16865, n16864, \Ki[0] , n16863, 
            \Kp[0] , n16862, n16853, n17031, n17030, n17029, n17028, 
            n17027, n17026, n17025, n17024, n17023, n17022, n17021, 
            n17020, n17019, n17018, n17017, n17016, n16967, n16966, 
            n16965, n16964, n16963, n16962, n16961, n16960, n16959, 
            n16958, n16957, n16956, n16955, n16954, n16953, n16952, 
            n16935, n16934, n16933, n16932, n16931, n16930, n16929, 
            n16928, n18701, n29541, n29542, n29538, n29539, n6, 
            \r_SM_Main[1] , tx_o, n4, n16871, n8947, tx_enable, 
            n16710, n16802, n21215, n4_adj_4, r_Rx_Data, n4_adj_5, 
            \r_Bit_Index[0] , n15595, RX_N_2, n15590, n4_adj_6, n17376, 
            n17380, n16861, n16860, n16859, n16858, n16857, n16856, 
            n16855) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[24] ;
    input GND_net;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[15] ;
    output [23:0]setpoint;
    input clk32MHz;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[12] ;
    output n63;
    output n771;
    input n63_adj_3;
    output \FRAME_MATCHER.i_31__N_2364 ;
    output n29497;
    output \FRAME_MATCHER.state[0] ;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[2] ;
    output n12869;
    output n2329;
    output n4452;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[1] ;
    output \FRAME_MATCHER.i_31__N_2370 ;
    output [23:0]PWMLimit;
    input \duty_23__N_3516[14] ;
    output n29;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[18] ;
    output \FRAME_MATCHER.state[3] ;
    output tx_active;
    output \FRAME_MATCHER.state[2] ;
    output rx_data_ready;
    input n16911;
    output [7:0]\data_in_frame[21] ;
    input n16910;
    input n16909;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[7] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[8] ;
    output n4218;
    input n16908;
    input n16907;
    output [7:0]\data_in_frame[9] ;
    output \data_in_frame[9][5] ;
    output \data_in_frame[9][4] ;
    output \data_in_frame[9][3] ;
    output \data_in_frame[9][2] ;
    output \data_in_frame[9][1] ;
    output \data_in_frame[9][0] ;
    input n16906;
    output n78;
    input n16905;
    input n16904;
    input n16903;
    output [7:0]control_mode;
    input n16902;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[5] ;
    input n16901;
    output [7:0]\data_in_frame[15] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[14] ;
    input n16900;
    input n16899;
    output n12944;
    output \data_in_frame[10][1] ;
    output n2;
    output DE_c;
    output n8868;
    input n16898;
    input n16897;
    input n16896;
    input n16894;
    input n16893;
    input n16892;
    input n16891;
    input n16890;
    input n16889;
    input n16888;
    input n16887;
    input n16886;
    input n16885;
    input n16884;
    input n16882;
    input n16881;
    input n16880;
    input n16879;
    input n16878;
    input n16877;
    input n16876;
    input n16875;
    input n16874;
    input n35073;
    input n28937;
    input n16867;
    input VCC_net;
    input n17373;
    output [23:0]IntegralLimit;
    input n17372;
    input n17371;
    input n17370;
    input n17369;
    input n17368;
    input n17367;
    input n17335;
    input n17334;
    input n17333;
    input n17332;
    input n17331;
    input n17330;
    input n17329;
    input n17328;
    input n17327;
    input n17326;
    input n17325;
    input n17324;
    input n17323;
    input n17322;
    input n17321;
    input n17320;
    input n17314;
    input n17313;
    input n17312;
    input n17311;
    input n17310;
    input n17309;
    input n17308;
    input n17307;
    input n17306;
    input n17305;
    input n17304;
    input n17303;
    input n17302;
    input n17301;
    input n17300;
    input n17299;
    input n17298;
    input n17297;
    input n17296;
    input n17295;
    input n17294;
    input n17293;
    input n17292;
    input n17291;
    input n17290;
    input n17289;
    input n17288;
    input n17287;
    input n17286;
    input n17285;
    input n17284;
    input n17283;
    output \Kp[1] ;
    input n17282;
    output \Kp[2] ;
    input n17281;
    output \Kp[3] ;
    input n17280;
    output \Kp[4] ;
    input n17279;
    output \Kp[5] ;
    input n17278;
    output \Kp[6] ;
    input n17277;
    output \Kp[7] ;
    input n17276;
    output \Kp[8] ;
    input n17275;
    output \Kp[9] ;
    input n17274;
    output \Kp[10] ;
    input n17273;
    output \Kp[11] ;
    input n17272;
    output \Kp[12] ;
    input n17271;
    output \Kp[13] ;
    input n17270;
    output \Kp[14] ;
    input n17269;
    output \Kp[15] ;
    input n17268;
    output \Ki[1] ;
    input n17267;
    output \Ki[2] ;
    input n17266;
    output \Ki[3] ;
    input n17265;
    output \Ki[4] ;
    input n17264;
    output \Ki[5] ;
    input n17263;
    output \Ki[6] ;
    input n17262;
    output \Ki[7] ;
    input n17261;
    output \Ki[8] ;
    input n17260;
    output \Ki[9] ;
    input n17259;
    output \Ki[10] ;
    input n17258;
    output \Ki[11] ;
    input n17257;
    output \Ki[12] ;
    input n17256;
    output \Ki[13] ;
    input n17255;
    output \Ki[14] ;
    input n17254;
    output \Ki[15] ;
    input n17253;
    input n17252;
    input n17251;
    input n17250;
    input n17249;
    input n17248;
    input n17247;
    input n17246;
    input n17245;
    input n17244;
    input n17243;
    input n17242;
    input n17241;
    input n17240;
    input n17239;
    input n17238;
    input n17237;
    input n17236;
    input n17235;
    input n17234;
    input n17233;
    input n17232;
    output n4216;
    output n122;
    output n5;
    output n35368;
    input n17231;
    input n17230;
    input n17229;
    input n17228;
    input n17227;
    input n17226;
    input n17225;
    input n17224;
    input n17223;
    input n17222;
    input n17221;
    input n17220;
    input n17219;
    input n17218;
    input n17217;
    input n17216;
    input n17215;
    input n17214;
    input n17213;
    input n17212;
    input n17211;
    input n17210;
    input n17209;
    input n17208;
    input n17207;
    input n17206;
    input n17205;
    input n17204;
    input n17203;
    input n17202;
    input n17201;
    input n17200;
    input n17199;
    input n17198;
    input n17197;
    input n17196;
    input n17195;
    input n17194;
    input n17193;
    input n17192;
    input n17191;
    input n17190;
    input n17189;
    input n17188;
    input n17187;
    input n17186;
    input n17185;
    input n17184;
    input n17183;
    input n17182;
    input n17181;
    input n17180;
    input n17179;
    input n17178;
    input n17177;
    input n17176;
    input n17175;
    input n17174;
    input n17173;
    input n17172;
    input n17171;
    input n17170;
    input n17169;
    input n17168;
    input n17167;
    input n17166;
    input n17165;
    input n17164;
    input n17163;
    input n17162;
    input n17161;
    input n17160;
    input n17159;
    input n17158;
    input n17157;
    input n17156;
    input n17155;
    input n17154;
    input n17153;
    input n17152;
    input n17151;
    input n17150;
    input n17149;
    input n17148;
    input n17147;
    input n17146;
    input n17145;
    input n17144;
    input n17143;
    input n17142;
    input n17141;
    input n17140;
    input n17139;
    input n17138;
    input n17137;
    input n17136;
    input n17135;
    input n17134;
    input n17133;
    input n17132;
    input n17131;
    input n17130;
    input n17129;
    input n17128;
    input n17127;
    input n17126;
    input n17125;
    input n17124;
    input n17123;
    input n17122;
    input n17121;
    input n17120;
    input n17119;
    input n17118;
    input n17117;
    input n17116;
    output n29535;
    input n17115;
    input n17114;
    input n17113;
    input n17112;
    input n17111;
    output LED_c;
    input n17110;
    output n29532;
    input n17109;
    input n17108;
    input n17107;
    input n17106;
    input n17105;
    input n17104;
    input n17103;
    input n17102;
    input n17101;
    output [23:0]neopxl_color;
    input n17100;
    input n17099;
    input n17098;
    input n17097;
    input n17096;
    input n17095;
    input n17094;
    input n17093;
    input n17092;
    input n17091;
    input n17090;
    input n17089;
    input n17088;
    input n17087;
    input n17086;
    input n17085;
    input n17084;
    input n17083;
    input n17082;
    input n17081;
    input n17080;
    input n17079;
    input n16865;
    input n16864;
    output \Ki[0] ;
    input n16863;
    output \Kp[0] ;
    input n16862;
    input n16853;
    input n17031;
    input n17030;
    input n17029;
    input n17028;
    input n17027;
    input n17026;
    input n17025;
    input n17024;
    input n17023;
    input n17022;
    input n17021;
    input n17020;
    input n17019;
    input n17018;
    input n17017;
    input n17016;
    input n16967;
    input n16966;
    input n16965;
    input n16964;
    input n16963;
    input n16962;
    input n16961;
    input n16960;
    input n16959;
    input n16958;
    input n16957;
    input n16956;
    input n16955;
    input n16954;
    input n16953;
    input n16952;
    input n16935;
    input n16934;
    input n16933;
    input n16932;
    input n16931;
    input n16930;
    input n16929;
    input n16928;
    output n18701;
    output n29541;
    output n29542;
    output n29538;
    output n29539;
    output n6;
    output \r_SM_Main[1] ;
    output tx_o;
    output n4;
    input n16871;
    output n8947;
    output tx_enable;
    output n16710;
    output n16802;
    output n21215;
    output n4_adj_4;
    output r_Rx_Data;
    output n4_adj_5;
    output \r_Bit_Index[0] ;
    output n15595;
    input RX_N_2;
    output n15590;
    output n4_adj_6;
    input n17376;
    input n17380;
    input n16861;
    input n16860;
    input n16859;
    input n16858;
    input n16857;
    input n16856;
    input n16855;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n27980, n27954, n29800, n29864, n15666, n29939, n15726, 
        n2206, n18, n27912, n13916, n16, n27019, n30142, n20, 
        n29949, n28013, n31916, n30124, n29974, n29841, n10, n29913, 
        n15291, n31868, n29654, n30020, n16396, n29669, n6_c, 
        n29851, n29952, n31438, n24886;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n24887, n4016, n16631, n30164, n30002, n30240, n6_adj_3606, 
        n30057, n15266, n29584, n2_c, n3, n16920;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n15853, n16500, n12, n29854, n28046, n30149, n30150, 
        n15990, n29999, n1179, n14, n29627, n10_adj_3607, n30252, 
        n27956, n27076, n30014, n16034, n27239, n30641, n31430, 
        n29993, n14_adj_3608, n29996, n15, n29965, n29942, n15979, 
        n16919;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n27952, n30136, n6_adj_3609, n27664, n10_adj_3610, n16054, 
        n29892, n31034;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n19, n4017, n30060, n27972, n14_adj_3611, n29751, n15791, 
        n13, n29857, n2112, n29816, n27982, n15785, n4018, n6_adj_3612, 
        n29777, n30075, n29639, n12_adj_3613, n30170, n29642;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n33458, n26741, n30005, n29774, n1383, n27108, n27479, 
        n5_c, n33045, n7, n16426, n4019, n30026, n29684, n12_adj_3614, 
        n29867, n34660, n34804, n14_adj_3615, n34768, n33188, n30118, 
        n10_adj_3616, n29822, n6_adj_3617, n6_adj_3618, n5_adj_3619, 
        n1260, n15751, n30078, n29962, n7_adj_3620, n4020, n6_adj_3621, 
        n15366, n14_adj_3622, n15_adj_3623, n34702, n34618, n14_adj_3624, 
        n34774, n33195, n30204, n30099, n6_adj_3625, n42, n46, 
        n44, n36, n45, n16250, n29644, n43, n29793, n15633, 
        n48, n52, n26989, n27063, n47, n30198, n22, n15_adj_3626, 
        n20_adj_3627, n16592, n24, n16161, n29572, n16_adj_3628, 
        n30189, n17, n6_adj_3629, n2125, n29839, n6_adj_3630, n31807, 
        n6_adj_3631, n5_adj_3632, n6_adj_3633, n27938, n7_adj_3634, 
        n34708, n34696, n14_adj_3635, n34726, n33148, n27652, n10_adj_3636, 
        n12_adj_3637, n27053, n30139, n6_adj_3638, n30133, n30222, 
        n6_adj_3639, n33484, n30207, n29601, n12_adj_3640, n29681, 
        n1516, n5_adj_3641, n7_adj_3642, n4021, n34594, n34684, 
        n14_adj_3643, n34732, n33151, n14_adj_3644, n10_adj_3645, 
        n27050, n16461, n30105, n16_adj_3646, n29980, n17_adj_3647, 
        n29624, n16_adj_3648, n30087, n30045, n22_adj_3649, n30234, 
        n20_adj_3650, n30161, n24_adj_3651, n29729, n10_adj_3652, 
        n29589, n1380, n6_adj_3653, n16479, n6_adj_3654, n16146, 
        n8, n1519, n12_adj_3655, n29946, n6_adj_3656, n6_adj_3657, 
        n2128, n29675, n29921, n27930, n16070, n16918;
    wire [31:0]n33;
    wire [31:0]\FRAME_MATCHER.state_31__N_2404 ;
    
    wire n9017, \FRAME_MATCHER.i_31__N_2368 , n3303, n5_adj_3658, n5_adj_3660, 
        n34932;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n32236, n32270, n29447, n29504, n18_adj_3661, n30, n28, 
        n32272, n27;
    wire [31:0]\FRAME_MATCHER.state_31__N_2468 ;
    
    wire n7_adj_3662, n31275, n29199, n5_adj_3663, n29015, n4_c, 
        n29109, n29013, n29111, n29011, n29113, n29009, n29115, 
        n29007, n29117, n29005, n29119, n29003, n29121, n29001, 
        n29123, n28999, n29125, n7_adj_3664, n7_adj_3665, n28997, 
        n29127, n28995, n29129, n29017, n29107, n28993, n29131, 
        n28991, n29133, n28989, n29135, n28987, n29137, n28985, 
        n29139, n28983, n29141, n28981, n29143, n28979, n29145, 
        n28977, n4022, n29147, n28975, n29149, n28949, n29151, 
        n28973, n29153, n28971, n29155, n15542, n15459, n5_adj_3666, 
        n14_adj_3667, n10_adj_3668, n8_adj_3669, n67, n117, n16_adj_3670, 
        n6_adj_3671, n33102, n1733, n89, n115, n4_adj_3672, tx_transmit_N_3257, 
        n44_adj_3673, n42_adj_3674, n43_adj_3675, n41, n40, n39, 
        n50, n45_adj_3676, n6_adj_3677, n8_adj_3678, n14_adj_3679, 
        n15610, n15_adj_3680, n15462, n16_adj_3681, n17_adj_3682, 
        n15539, n31109, n10_adj_3683, n10_adj_3684, n14_adj_3685, 
        n15583, n18_adj_3686, n20_adj_3687, n15_adj_3688, n63_adj_3689, 
        n16_adj_3690, n17_adj_3691, n63_adj_3692, n20_adj_3693, n19_adj_3694, 
        n32264, n2_adj_3695, n884, \FRAME_MATCHER.i_31__N_2367 , n29019, 
        n29105, n16917, n16_adj_3696, n17_adj_3697, n4023, n23888, 
        n16916, n16915, n16914, n2_adj_3698, n24885, n10_adj_3699, 
        n29543, n16968, n4024, n30352;
    wire [2:0]r_SM_Main_2__N_3360;
    
    wire n21130, n29513, n114, n4_adj_3700, n22109, n31265, n10_adj_3701, 
        n16695;
    wire [0:0]n2863;
    
    wire n16913, n33187, n33186, n4025, n4026, n4027, n4028, n16912, 
        n21855, \FRAME_MATCHER.rx_data_ready_prev , n2_adj_3702, n24884;
    wire [7:0]n8825;
    
    wire n16652, n16773, n16_adj_3703, n4029, n29726, Kp_23__N_764, 
        n10_adj_3704, n17_adj_3705, n16245, n12_adj_3706, n22_adj_3707, 
        n16604, n29905, n16107, n16329, n24_adj_3708, n30011, n12_adj_3709, 
        n23, n30173, n15905, n27783, n29635, n25, n15856, n23828, 
        n1, n4030, n4031;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n4032, n16_adj_3710, n17_adj_3711, n4033, n4034, n4035, 
        n33170, n33169, n4036, n4037, n4038, n16969, n16_adj_3712, 
        n17_adj_3713, n4039, n29555, n17000;
    wire [7:0]\data_in_frame[9]_c ;   // verilog/coms.v(96[12:25])
    
    wire n17001, n17002, n8_adj_3714, n8_adj_3715, n28941, n28947, 
        n17003, n2_adj_3716, n24883, n92, n32156, n2_adj_3717, n24882, 
        n17004, n17005;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n32159, n31247, n17006, n17007, n2_adj_3718, n24881, n10_adj_3719, 
        n2_adj_3720, n24880, n2_adj_3721, n24879, n30501, n31011;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n31372, n29835, n31099, n16060, n31955, n30676, n30802, 
        n2_adj_3722, n3_adj_3723, n2_adj_3724, n24878, n2_adj_3725, 
        n3_adj_3726, n2_adj_3727, n3_adj_3728, n2_adj_3729, n3_adj_3730, 
        n2_adj_3731, n3_adj_3732, n2_adj_3733, n3_adj_3734, n2_adj_3735, 
        n3_adj_3736, n2_adj_3737, n3_adj_3738, n2_adj_3739, n3_adj_3740, 
        n3_adj_3741, n3_adj_3742, n3_adj_3743, n3_adj_3744, n3_adj_3745, 
        n3_adj_3746, n3_adj_3747, n3_adj_3748, n2_adj_3749, n3_adj_3750, 
        n2_adj_3751, n3_adj_3752, n2_adj_3753, n3_adj_3754, n2_adj_3755, 
        n3_adj_3756, n2_adj_3757, n3_adj_3758, n2_adj_3759, n3_adj_3760, 
        n2_adj_3761, n3_adj_3762, n2_adj_3763, n3_adj_3764, n2_adj_3765, 
        n3_adj_3766, n2_adj_3767, n3_adj_3768, n2_adj_3769, n3_adj_3770, 
        n2_adj_3771, n3_adj_3772, n2_adj_3773, n3_adj_3774, n2_adj_3775, 
        n3_adj_3776, n18487, n6_adj_3777, n33167, n33166, n161, 
        n21151, n29530, n18751, n24877, n24876, n15811, n16220, 
        n29971, n10_adj_3778, n29552, n16992, n16993, n16994, n24875, 
        n16493, n16094, n16995, n27936, n29609, n6_adj_3779, n29984, 
        n27918, n30231, n16445, n29767, n29797, n18_adj_3780, n29771, 
        n29884, n20_adj_3781, n29930, Kp_23__N_1261;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n30246, n30039, n30067, n42_adj_3782, n29604, n60, n58, 
        n68, n64, n29870, n62, n63_adj_3783, n30192, n30255, n30051, 
        n61, n30090, n29666, n29711, n15714, n66;
    wire [7:0]\data_in_frame[10]_c ;   // verilog/coms.v(96[12:25])
    
    wire n34034, n72, n30201, n15951, n29672, n65, n73, n31528, 
        n30249, n16_adj_3784, n30130, n27106, n19_adj_3785, n29927, 
        n22_adj_3786, n17_adj_3787, n27633, n30807, n30530, n30258, 
        n10_adj_3788, n30195, n27550, n29707, n15768, n30179, n27986, 
        Kp_23__N_1054, Kp_23__N_1026, n15918, n30023, n10_adj_3789, 
        Kp_23__N_1035, n9, n29848, n15777, n29717, n26977, Kp_23__N_1050, 
        n30111, n14_adj_3790, n15947, n15643, n13_adj_3791, n14_adj_3792, 
        n30114, n15_adj_3793, n30213, n6_adj_3794, n16011, n27061, 
        n30084, n30145, n12_adj_3795, n27008, n30219, n11, n16353, 
        n10_adj_3796, n16204, n28008, n14_adj_3797, n9_adj_3798, n29698, 
        n16333, n12_adj_3799, n8_adj_3800, n29928, n27683, n27944, 
        n29959, n29813, n16996, n29754, n15866, n29744, n6_adj_3801, 
        n31643, n7_adj_3802, n24_adj_3803, n22_adj_3804, n23_adj_3805, 
        n29787, n30081, n21, n29790, n30228, n6_adj_3806, n26998, 
        n27940, n16098, Kp_23__N_605, n29881, n10_adj_3807, n27402, 
        n29878, n8_adj_3808, n29764, n30186, n29825, n29910, n34, 
        n12_adj_3809, n30036, n29915, n16368, n4_adj_3810, n30216, 
        n28034, n29736, n30183, n14041, n10_adj_3812, n16267, n16280, 
        n29598, n8_adj_3813, n29546, n24_adj_3814, n38, n29834, 
        n29723, n36_adj_3815, n14048, n15941, n30070, n6_adj_3816, 
        n6_adj_3817, n29784, n10_adj_3818, n8_adj_3819, n29549, n8_adj_3820, 
        n29924, n14_adj_3821, n29663, n5_adj_3822, n28040, n22_adj_3823, 
        n37, n15914, n27996, n16192, n20_adj_3824, n18_adj_3825, 
        n22_adj_3826, n29875, n10_adj_3827, n30210, n14_adj_3828, 
        n10_adj_3829, n28001, n27959, n8_adj_3830, n31862, n29714, 
        n10_adj_3831, n9_adj_3832, n20_adj_3833, n16336, n19_adj_3834, 
        n21_adj_3835, n29902, n35, n6_adj_3836, n29632, n12_adj_3837, 
        n10_adj_3838, n29918, n31198, n29861, n6_adj_3839, n31486, 
        n7_adj_3840, n6_adj_3841, n31772, n31071, n27961, n31237, 
        n31201, n30612, n6_adj_3842, n6_adj_3843, n30590, n29733, 
        n30048, n10_adj_3844, n27992, n27093, n4_adj_3845, n13173, 
        n30_adj_3846, n30127, n28003, n10_adj_3847, n6_adj_3848, n32224, 
        n8_adj_3849, n22_adj_3850, n32226, n31240, n21_adj_3851, n6_adj_3852, 
        n31935, n32230, n26, n30_adj_3853, n17_adj_3854, n16997, 
        n16944, n16945, n16946, n29700, n24874, n27977, n6_adj_3855, 
        n16998, n16947, n16999, n30093, Kp_23__N_912, n15823, n30029, 
        n34801, n34534, n34795;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n31856, n6_adj_3856, n16948, n29898, n16949, n16950, n30017, 
        n30176, n10_adj_3857, n29621, n19_adj_3858, n15890, n34540, 
        n34789, n10_adj_3859, n34783, n34786, n34777, n34780, Kp_23__N_958, 
        n6_adj_3860, n34771, n27067, n2143, n29595, n14_adj_3861, 
        n34765, n13_adj_3862, n16951, n34759, n16936, n30096, n16937, 
        n16970, n30108, n29660, n16938, n16939, n14_adj_3863, n10_adj_3864, 
        n34762, n34753, n34756, n34747, n34750, n12_adj_3865, n34741, 
        n34744, n29647, n34735, n34738, n3_adj_3866, n34729, n16940, 
        n16941, n16942, n16943, n29689, n34723, n29692, n34705, 
        n34699, n30243, n15720, n34693, n10_adj_3867, n29558, n17072, 
        n34687, n34690, n34681, n17073, n10_adj_3868, n20_adj_3869, 
        n34669, n34672, n17074, n17075, Kp_23__N_737, n32, n17076, 
        n30_adj_3870, n17077, n17078, n16866, n31, n29_adj_3871, 
        n17388, n29934, n34657, n34546, n34651, n29810, n34552, 
        n34645, n29968, n29831, n34558, n33171, n34639, n14_adj_3872, 
        n7_adj_3873, n34564, n33168, n34633, n14_adj_3874, n7_adj_3875, 
        n34570, n33165, n34627, n14_adj_3876, n7_adj_3877, n34576, 
        n33159, n34621, n14_adj_3878, n7_adj_3879, n24873, n34615, 
        n29740, n10_adj_3880, n24872, n34591, n34585, n34588, n34579, 
        n34582, n24871, n24870, n10_adj_3881, n29837, n24869, n24901, 
        n16_adj_3882, n24868, n24900, n24899, n17_adj_3883, n24867, 
        n24898, n24866, n24897, n24896, n24865, n16971, n24895, 
        n24864, n24894, n24893, n24892, n33160, n33161, n34573, 
        n24891, n24890, n16895, n16883, n16868, n16972, n30102, 
        n16984, n16985, n16986, n34567, n16987, n16921, n16922, 
        n16923, n16924, n16925, n16926, n16927, n16988, n16989, 
        n59, n30439, n12_adj_3885, n16990, n24889, n34561, n24888, 
        n28050, n17071, n34555, n17070, n17069, n17068, n17067, 
        n17066, n17065, n17064, n17063, n17062, n17061, n17060, 
        n17059, n17058, n17057, n17056, n17055, n17054, n17053, 
        n17052, n17051, n17050, n17049, n17048, n17047, n17046, 
        n17045, n17044, n17043, n17042, n17041, n17040, n17039, 
        n17038, n17037, n17036, n17035, n17034, n17033, n17032, 
        n17015, n17014, n17013, n17012, n17011, n17010, n17009, 
        n17008, n16991, n16983, n16982, n16981, n16980, n31783, 
        n16979, n16978, n16977, n16976, n16975, n16974, n16973, 
        n28_adj_3886, n33193, n33194, n34549, n17_adj_3887, n16_adj_3888, 
        n26_adj_3889, n33196, n33197, n34543, n27_adj_3890, n17_adj_3891, 
        n16_adj_3892, n25_adj_3893, n33149, n33150, n34537, n17_adj_3894, 
        n16_adj_3895, n33152, n33153, n34531, n17_adj_3896, n16_adj_3897, 
        n10_adj_3898, n12_adj_3899, n13_adj_3900, n34519, n34522, 
        n33478, n5_adj_3901, n6_adj_3902, n5_adj_3903, n6_adj_3904, 
        n5_adj_3905, n6_adj_3906, n5_adj_3907;
    
    SB_LUT4 i3_4_lut (.I0(n27980), .I1(n27954), .I2(\data_out_frame[23] [7]), 
            .I3(n29800), .O(n29864));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[24] [5]), .I1(n15666), .I2(GND_net), 
            .I3(GND_net), .O(n29939));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_838 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15726));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_838.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut (.I0(n15726), .I1(n2206), .I2(n29939), .I3(\data_out_frame[24] [0]), 
            .O(n18));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(n27912), .I1(n13916), .I2(GND_net), .I3(GND_net), 
            .O(n16));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut (.I0(n27019), .I1(n18), .I2(n29864), .I3(n30142), 
            .O(n20));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n29949), .I1(n20), .I2(n16), .I3(n28013), 
            .O(n31916));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_839 (.I0(n31916), .I1(\data_out_frame[25] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30124));
    defparam i1_2_lut_adj_839.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut (.I0(n29974), .I1(n29841), .I2(\data_out_frame[25] [4]), 
            .I3(n30124), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n29913), .I1(n10), .I2(n15291), .I3(GND_net), 
            .O(n31868));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[20] [2]), .I1(n29654), .I2(\data_out_frame[18] [0]), 
            .I3(GND_net), .O(n30020));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_840 (.I0(\data_out_frame[17] [6]), .I1(n16396), 
            .I2(n29669), .I3(n6_c), .O(n15666));
    defparam i4_4_lut_adj_840.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_841 (.I0(n15666), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [6]), .I3(GND_net), .O(n29851));
    defparam i2_3_lut_adj_841.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_842 (.I0(\data_out_frame[25] [1]), .I1(n29952), 
            .I2(n29851), .I3(\data_out_frame[23] [0]), .O(n31438));
    defparam i3_4_lut_adj_842.LUT_INIT = 16'h6996;
    SB_CARRY add_43_25 (.CI(n24886), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n24887));
    SB_LUT4 i1_2_lut_adj_843 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n29669));
    defparam i1_2_lut_adj_843.LUT_INIT = 16'h6666;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n16631), .D(n4016));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_844 (.I0(n30164), .I1(n30002), .I2(n30240), .I3(n6_adj_3606), 
            .O(n30057));
    defparam i4_4_lut_adj_844.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_845 (.I0(n15266), .I1(\data_out_frame[24] [7]), 
            .I2(\data_out_frame[23] [0]), .I3(GND_net), .O(n29584));
    defparam i2_3_lut_adj_845.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_c), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n16920));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_846 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n15853));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[18] [2]), .I1(n30057), .I2(n16500), 
            .I3(n29669), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[17] [7]), .I1(n12), .I2(\data_out_frame[20] [3]), 
            .I3(n29854), .O(n28046));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_847 (.I0(n29974), .I1(n30149), .I2(GND_net), 
            .I3(GND_net), .O(n30150));
    defparam i1_2_lut_adj_847.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_848 (.I0(n15990), .I1(n29999), .I2(n1179), .I3(\data_out_frame[5] [0]), 
            .O(n14));
    defparam i6_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_849 (.I0(n29627), .I1(n14), .I2(n10_adj_3607), 
            .I3(n30252), .O(n29654));
    defparam i7_4_lut_adj_849.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_850 (.I0(n27956), .I1(\data_out_frame[23] [1]), 
            .I2(\data_out_frame[23] [0]), .I3(GND_net), .O(n30149));
    defparam i2_3_lut_adj_850.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_851 (.I0(\data_out_frame[25] [3]), .I1(n30149), 
            .I2(n27076), .I3(GND_net), .O(n29841));
    defparam i2_3_lut_adj_851.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_852 (.I0(\data_out_frame[20] [4]), .I1(n30014), 
            .I2(n29654), .I3(n16034), .O(n27239));
    defparam i3_4_lut_adj_852.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_853 (.I0(n27239), .I1(n29841), .I2(n30641), .I3(\data_out_frame[25] [2]), 
            .O(n31430));
    defparam i3_4_lut_adj_853.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_854 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n30164));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_854.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_855 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[16] [1]), 
            .I2(n29993), .I3(GND_net), .O(n14_adj_3608));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_855.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_856 (.I0(n30164), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[5] [1]), .I3(n29996), .O(n15));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_856.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n29965), .I2(n14_adj_3608), .I3(\data_out_frame[5] [3]), 
            .O(n16500));   // verilog/coms.v(85[17:28])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_857 (.I0(\data_out_frame[16] [4]), .I1(n29942), 
            .I2(\data_out_frame[18] [4]), .I3(n15979), .O(n27912));
    defparam i3_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n16919));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_858 (.I0(n27952), .I1(\data_out_frame[19] [0]), 
            .I2(n30136), .I3(n6_adj_3609), .O(n30641));
    defparam i4_4_lut_adj_858.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_859 (.I0(n27912), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29952));
    defparam i1_2_lut_adj_859.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_860 (.I0(\data_out_frame[16] [3]), .I1(n16500), 
            .I2(\data_out_frame[20] [5]), .I3(n27664), .O(n10_adj_3610));
    defparam i4_4_lut_adj_860.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_861 (.I0(\data_out_frame[18] [3]), .I1(n10_adj_3610), 
            .I2(\data_out_frame[18] [4]), .I3(GND_net), .O(n27956));
    defparam i5_3_lut_adj_861.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_862 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16054));
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_863 (.I0(n27956), .I1(n29952), .I2(n30641), .I3(GND_net), 
            .O(n15266));
    defparam i2_3_lut_adj_863.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29892));
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_865 (.I0(n27076), .I1(n29892), .I2(n15291), .I3(GND_net), 
            .O(n31034));
    defparam i2_3_lut_adj_865.LUT_INIT = 16'h6969;
    SB_LUT4 mux_987_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n4017));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_866 (.I0(n30060), .I1(n27972), .I2(\data_out_frame[18] [4]), 
            .I3(\data_out_frame[18] [5]), .O(n14_adj_3611));
    defparam i6_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_867 (.I0(\data_out_frame[18] [7]), .I1(n29751), 
            .I2(\data_out_frame[18] [6]), .I3(n15791), .O(n13));
    defparam i5_4_lut_adj_867.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(\data_out_frame[17] [5]), .I1(n13), .I2(n14_adj_3611), 
            .I3(GND_net), .O(n29857));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_868 (.I0(n2112), .I1(n29857), .I2(GND_net), .I3(GND_net), 
            .O(n30136));
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_869 (.I0(n27980), .I1(n29816), .I2(GND_net), 
            .I3(GND_net), .O(n27982));
    defparam i1_2_lut_adj_869.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_870 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n15785));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_870.LUT_INIT = 16'h6666;
    SB_LUT4 mux_987_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19] [2]), .O(n4018));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_871 (.I0(\data_out_frame[19] [6]), .I1(n15785), 
            .I2(\data_out_frame[19] [4]), .I3(n6_adj_3612), .O(n2112));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_872 (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15791));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_872.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_873 (.I0(n29777), .I1(n30075), .I2(\data_out_frame[11] [7]), 
            .I3(n29639), .O(n12_adj_3613));
    defparam i5_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_874 (.I0(\data_out_frame[5] [0]), .I1(n12_adj_3613), 
            .I2(n30170), .I3(\data_out_frame[11] [6]), .O(n15979));
    defparam i6_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_875 (.I0(n15979), .I1(n15791), .I2(GND_net), 
            .I3(GND_net), .O(n30014));
    defparam i1_2_lut_adj_875.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_876 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[14] [5]), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n29642));
    defparam i2_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_877 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[14] [0]), 
            .I2(\data_out_frame[14] [1]), .I3(GND_net), .O(n30075));
    defparam i2_3_lut_adj_877.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_878 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n30252));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_878.LUT_INIT = 16'h9696;
    SB_LUT4 i27784_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33458));   // verilog/coms.v(106[34:55])
    defparam i27784_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_4_lut_adj_879 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [2]), 
            .I2(n26741), .I3(\data_out_frame[15] [3]), .O(n30005));
    defparam i3_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_880 (.I0(\data_out_frame[13] [1]), .I1(n29774), 
            .I2(n1383), .I3(n27108), .O(n27479));
    defparam i3_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_4_lut (.I0(n5_c), .I1(n33458), 
            .I2(n33045), .I3(byte_transmit_counter[0]), .O(n7));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1_2_lut_adj_881 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16426));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_881.LUT_INIT = 16'h6666;
    SB_LUT4 mux_987_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n4019));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_4_lut_adj_882 (.I0(\data_out_frame[6] [5]), .I1(n16426), 
            .I2(n30026), .I3(n29684), .O(n12_adj_3614));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_883 (.I0(\data_out_frame[6] [3]), .I1(n12_adj_3614), 
            .I2(n29867), .I3(\data_out_frame[10] [5]), .O(n27108));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i1816161_i1_3_lut (.I0(n34660), .I1(n34804), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3615));
    defparam i1816161_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_884 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n30240));
    defparam i2_3_lut_adj_884.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_885 (.I0(\data_out_frame[9] [1]), .I1(n30240), 
            .I2(\data_out_frame[9] [5]), .I3(\data_out_frame[13] [7]), .O(n29965));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_885.LUT_INIT = 16'h6996;
    SB_LUT4 i27790_2_lut (.I0(n34768), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33188));
    defparam i27790_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_886 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n29867));
    defparam i1_2_lut_adj_886.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_887 (.I0(n29867), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[13] [2]), .I3(n30118), .O(n10_adj_3616));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_888 (.I0(\data_out_frame[13] [3]), .I1(n16396), 
            .I2(GND_net), .I3(GND_net), .O(n29822));
    defparam i1_2_lut_adj_888.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_889 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[6] [6]), .I3(n6_adj_3617), .O(n29639));
    defparam i4_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3618));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'ha300;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3619));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i472_2_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1260));   // verilog/coms.v(85[17:28])
    defparam i472_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_890 (.I0(\data_out_frame[9] [3]), .I1(n29777), 
            .I2(n1260), .I3(n15751), .O(n15990));
    defparam i3_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_891 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30078));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_892 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n29962));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_893 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30026));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut (.I0(n5_adj_3619), 
            .I1(n6_adj_3618), .I2(n33045), .I3(GND_net), .O(n7_adj_3620));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_987_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19] [4]), .O(n4020));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[8] [7]), .O(n30118));   // verilog/coms.v(85[17:28])
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_894 (.I0(\data_out_frame[7] [0]), .I1(n30118), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n6_adj_3621));   // verilog/coms.v(85[17:28])
    defparam i1_3_lut_adj_894.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_895 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[6] [7]), 
            .I2(n30078), .I3(n6_adj_3621), .O(n15366));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_896 (.I0(\data_out_frame[13] [3]), .I1(n15366), 
            .I2(GND_net), .I3(GND_net), .O(n29854));
    defparam i1_2_lut_adj_896.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_897 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n14_adj_3622));   // verilog/coms.v(85[17:70])
    defparam i5_3_lut_adj_897.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_898 (.I0(n30026), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[5] [0]), .I3(n29962), .O(n15_adj_3623));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_899 (.I0(n15_adj_3623), .I1(\data_out_frame[7] [1]), 
            .I2(n14_adj_3622), .I3(\data_out_frame[9] [0]), .O(n16034));   // verilog/coms.v(85[17:70])
    defparam i8_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i1817970_i1_3_lut (.I0(n34702), .I1(n34618), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3624));
    defparam i1817970_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27786_2_lut (.I0(n34774), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33195));
    defparam i27786_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30204));
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\data_out_frame[17] [2]), .I1(n30099), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3625));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_902 (.I0(n30204), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[17] [1]), .I3(n6_adj_3625), .O(n30060));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i1418_2_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2206));   // verilog/coms.v(78[16:27])
    defparam i1418_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(n30078), .I3(\data_out_frame[6] [4]), .O(n42));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n15990), .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[10] [5]), 
            .I3(\data_out_frame[10] [0]), .O(n46));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[10] [3]), .I3(\data_out_frame[13] [4]), 
            .O(n44));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(\data_out_frame[6] [0]), .I1(n36), .I2(n29822), 
            .I3(\data_out_frame[5] [4]), .O(n45));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n16250), .I1(n29644), .I2(n29965), .I3(\data_out_frame[5] [5]), 
            .O(n43));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n27479), .I1(n42), .I2(n29793), .I3(n15633), 
            .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n27108), .I1(\data_out_frame[12] [2]), .I2(n26989), 
            .I3(n27063), .O(n47));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_903 (.I0(\data_out_frame[16] [5]), .I1(n30005), 
            .I2(n30198), .I3(\data_out_frame[14] [2]), .O(n22));
    defparam i9_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(n47), .I1(n30252), .I2(n52), .I3(n48), .O(n15_adj_3626));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i7_3_lut (.I0(\data_out_frame[16] [1]), .I1(n30075), .I2(\data_out_frame[16] [6]), 
            .I3(GND_net), .O(n20_adj_3627));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut (.I0(n15_adj_3626), .I1(n22), .I2(n29642), .I3(n16592), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[14] [7]), .I1(n24), .I2(n20_adj_3627), 
            .I3(n16161), .O(n27972));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_904 (.I0(n27972), .I1(n2206), .I2(n30060), .I3(n29572), 
            .O(n16_adj_3628));
    defparam i6_4_lut_adj_904.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_905 (.I0(\data_out_frame[18] [0]), .I1(n30014), 
            .I2(n30189), .I3(\data_out_frame[17] [7]), .O(n17));
    defparam i7_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_906 (.I0(n17), .I1(\data_out_frame[17] [5]), .I2(n16_adj_3628), 
            .I3(n2112), .O(n27952));
    defparam i9_4_lut_adj_906.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_907 (.I0(n26989), .I1(n27982), .I2(n30136), .I3(n6_adj_3629), 
            .O(n13916));
    defparam i4_4_lut_adj_907.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_908 (.I0(n27019), .I1(n2125), .I2(GND_net), .I3(GND_net), 
            .O(n29839));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_909 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [5]), 
            .I2(n29839), .I3(n6_adj_3630), .O(n31807));
    defparam i4_4_lut_adj_909.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_910 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n29684));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_910.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_911 (.I0(n29684), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[8] [5]), .O(n29774));   // verilog/coms.v(75[16:27])
    defparam i2_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i6_3_lut (.I0(\data_out_frame[5] [7]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n6_adj_3631));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3632));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_912 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[10] [6]), 
            .I2(n29774), .I3(n6_adj_3633), .O(n27063));
    defparam i4_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\data_out_frame[17] [2]), .I1(n27063), 
            .I2(GND_net), .I3(GND_net), .O(n27938));
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut (.I0(n5_adj_3632), 
            .I1(n6_adj_3631), .I2(n33045), .I3(GND_net), .O(n7_adj_3634));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1812543_i1_3_lut (.I0(n34708), .I1(n34696), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3635));
    defparam i1812543_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27717_2_lut (.I0(n34726), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33148));
    defparam i27717_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_914 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16161));
    defparam i1_2_lut_adj_914.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_915 (.I0(\data_out_frame[18] [5]), .I1(n27652), 
            .I2(GND_net), .I3(GND_net), .O(n29942));
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_916 (.I0(\data_out_frame[5] [3]), .I1(n10_adj_3636), 
            .I2(\data_out_frame[14] [1]), .I3(\data_out_frame[7] [2]), .O(n12_adj_3637));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_917 (.I0(n27053), .I1(n12_adj_3637), .I2(n29993), 
            .I3(\data_out_frame[13] [7]), .O(n27664));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_918 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15633));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_919 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[14] [5]), 
            .I2(n30139), .I3(n6_adj_3638), .O(n30133));
    defparam i4_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_920 (.I0(n27664), .I1(n29942), .I2(n16161), .I3(GND_net), 
            .O(n30222));
    defparam i2_3_lut_adj_920.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_921 (.I0(n27053), .I1(n26989), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3639));
    defparam i1_2_lut_adj_921.LUT_INIT = 16'h6666;
    SB_LUT4 i27361_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n33045));   // verilog/coms.v(106[34:55])
    defparam i27361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_922 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[16] [5]), .I3(n6_adj_3639), .O(n30189));
    defparam i4_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i27809_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33484));   // verilog/coms.v(106[34:55])
    defparam i27809_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30207));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_924 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[10] [2]), .I3(n29601), .O(n12_adj_3640));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_924.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_925 (.I0(\data_out_frame[6] [1]), .I1(n12_adj_3640), 
            .I2(n29681), .I3(\data_out_frame[7] [6]), .O(n1516));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3641));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_4_lut (.I0(n5_adj_3641), 
            .I1(n33484), .I2(n33045), .I3(byte_transmit_counter[0]), .O(n7_adj_3642));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 mux_987_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19] [5]), .O(n4021));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i389_2_lut (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1179));   // verilog/coms.v(73[16:27])
    defparam i389_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n29999));
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i1813146_i1_3_lut (.I0(n34594), .I1(n34684), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3643));
    defparam i1813146_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27815_2_lut (.I0(n34732), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33151));
    defparam i27815_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_927 (.I0(n30170), .I1(n15751), .I2(n29644), .I3(\data_out_frame[14] [2]), 
            .O(n14_adj_3644));
    defparam i6_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_928 (.I0(\data_out_frame[14] [3]), .I1(n14_adj_3644), 
            .I2(n10_adj_3645), .I3(n1179), .O(n27652));
    defparam i7_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_929 (.I0(\data_out_frame[17] [0]), .I1(n27050), 
            .I2(\data_out_frame[16] [7]), .I3(n16461), .O(n30105));
    defparam i3_4_lut_adj_929.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_930 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[12] [4]), 
            .I2(n30105), .I3(n27652), .O(n16_adj_3646));
    defparam i6_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_931 (.I0(\data_out_frame[16] [4]), .I1(n29980), 
            .I2(n30207), .I3(n16592), .O(n17_adj_3647));
    defparam i7_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_932 (.I0(n17_adj_3647), .I1(n1516), .I2(n16_adj_3646), 
            .I3(\data_out_frame[19] [0]), .O(n27019));
    defparam i9_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29996));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29627));
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_935 (.I0(n29627), .I1(n29996), .I2(\data_out_frame[9] [5]), 
            .I3(GND_net), .O(n29624));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_935.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3648));   // verilog/coms.v(76[16:27])
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_936 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [1]), 
            .I2(n30087), .I3(n30045), .O(n22_adj_3649));   // verilog/coms.v(76[16:27])
    defparam i9_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_adj_937 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[12] [1]), 
            .I2(n30234), .I3(GND_net), .O(n20_adj_3650));   // verilog/coms.v(76[16:27])
    defparam i7_3_lut_adj_937.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_938 (.I0(n30002), .I1(n22_adj_3649), .I2(n16_adj_3648), 
            .I3(n30161), .O(n24_adj_3651));   // verilog/coms.v(76[16:27])
    defparam i11_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_939 (.I0(\data_out_frame[5] [5]), .I1(n24_adj_3651), 
            .I2(n20_adj_3650), .I3(n29624), .O(n27053));   // verilog/coms.v(76[16:27])
    defparam i12_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_out_frame[16] [5]), .I1(n27053), 
            .I2(GND_net), .I3(GND_net), .O(n29980));
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_941 (.I0(\data_out_frame[9] [7]), .I1(n30234), 
            .I2(GND_net), .I3(GND_net), .O(n30045));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_942 (.I0(\data_out_frame[12] [3]), .I1(n30045), 
            .I2(\data_out_frame[6] [0]), .I3(n29729), .O(n10_adj_3652));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_943 (.I0(\data_out_frame[5] [7]), .I1(n10_adj_3652), 
            .I2(\data_out_frame[8] [1]), .I3(GND_net), .O(n26989));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_943.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30198));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_945 (.I0(n29589), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[8] [4]), .O(n1383));   // verilog/coms.v(73[16:34])
    defparam i2_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_946 (.I0(\data_out_frame[10] [4]), .I1(n1380), 
            .I2(\data_out_frame[10] [5]), .I3(GND_net), .O(n6_adj_3653));   // verilog/coms.v(85[17:28])
    defparam i1_3_lut_adj_946.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_947 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(n1383), .I3(n6_adj_3653), .O(n16479));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_948 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n29793));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_949 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n29681));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_950 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [3]), .I3(n6_adj_3654), .O(n1380));   // verilog/coms.v(73[16:34])
    defparam i4_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29601));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_952 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n29589));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_out_frame[10] [4]), .I1(n1380), 
            .I2(GND_net), .I3(GND_net), .O(n16146));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_954 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[8] [2]), .I3(n29601), .O(n8));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_955 (.I0(n16146), .I1(n8), .I2(\data_out_frame[5] [6]), 
            .I3(n29589), .O(n1519));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30161));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n29729));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29572));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_959 (.I0(\data_out_frame[12] [5]), .I1(n1519), 
            .I2(GND_net), .I3(GND_net), .O(n16250));
    defparam i1_2_lut_adj_959.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16461));
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_961 (.I0(\data_out_frame[10] [1]), .I1(n30087), 
            .I2(\data_out_frame[5] [6]), .I3(n29729), .O(n12_adj_3655));   // verilog/coms.v(75[16:43])
    defparam i5_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_962 (.I0(\data_out_frame[7] [5]), .I1(n12_adj_3655), 
            .I2(\data_out_frame[12] [2]), .I3(n29793), .O(n27050));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_963 (.I0(n29946), .I1(\data_out_frame[16] [7]), 
            .I2(n30139), .I3(n6_adj_3656), .O(n2125));
    defparam i4_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_964 (.I0(\data_out_frame[19] [2]), .I1(n27938), 
            .I2(n30105), .I3(n6_adj_3657), .O(n2128));
    defparam i4_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_965 (.I0(n2128), .I1(n2125), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n29675));
    defparam i2_3_lut_adj_965.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_966 (.I0(n27019), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29921));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_967 (.I0(n30189), .I1(n30222), .I2(n30133), .I3(GND_net), 
            .O(n27930));
    defparam i2_3_lut_adj_967.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16070));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_969 (.I0(n16070), .I1(n27930), .I2(n29921), .I3(n29675), 
            .O(n29913));
    defparam i3_4_lut_adj_969.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n16918));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i17142_2_lut (.I0(n33[1]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2404 [1]));   // verilog/coms.v(142[4] 144[7])
    defparam i17142_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4989_2_lut (.I0(n63), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n9017));   // verilog/coms.v(157[6] 159[9])
    defparam i4989_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_323_Select_1_i5_4_lut (.I0(n63), .I1(\FRAME_MATCHER.i_31__N_2368 ), 
            .I2(n3303), .I3(n33[1]), .O(n5_adj_3658));
    defparam select_323_Select_1_i5_4_lut.LUT_INIT = 16'hccc4;
    SB_LUT4 i1_4_lut_adj_970 (.I0(n63_adj_3), .I1(n33[1]), .I2(\FRAME_MATCHER.i_31__N_2364 ), 
            .I3(n9017), .O(n5_adj_3660));
    defparam i1_4_lut_adj_970.LUT_INIT = 16'hd5f5;
    SB_LUT4 i3_4_lut_adj_971 (.I0(n5_adj_3660), .I1(\FRAME_MATCHER.state_31__N_2404 [1]), 
            .I2(n5_adj_3658), .I3(n29497), .O(n34932));
    defparam i3_4_lut_adj_971.LUT_INIT = 16'hfefa;
    SB_LUT4 i26563_2_lut (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32236));
    defparam i26563_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26596_4_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[0] [1]), .O(n32270));
    defparam i26596_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_972 (.I0(\data_in_frame[0] [7]), .I1(n32270), .I2(n32236), 
            .I3(\data_in_frame[0] [3]), .O(n29447));
    defparam i7_4_lut_adj_972.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_adj_973 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n29504));
    defparam i1_2_lut_adj_973.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_974 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3661));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(n18_adj_3661), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i11_4_lut_adj_975 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[1] [7]), .O(n28));
    defparam i11_4_lut_adj_975.LUT_INIT = 16'h0080;
    SB_LUT4 i26598_4_lut (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[2] [1]), .O(n32272));
    defparam i26598_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_976 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [6]), .I3(n29447), .O(n27));
    defparam i10_4_lut_adj_976.LUT_INIT = 16'h4000;
    SB_LUT4 i16_4_lut_adj_977 (.I0(n27), .I1(n32272), .I2(n28), .I3(n30), 
            .O(\FRAME_MATCHER.state_31__N_2468 [3]));
    defparam i16_4_lut_adj_977.LUT_INIT = 16'h2000;
    SB_LUT4 i1_4_lut_adj_978 (.I0(\FRAME_MATCHER.state_31__N_2468 [3]), .I1(n7_adj_3662), 
            .I2(n31275), .I3(n29504), .O(n29199));   // verilog/coms.v(112[11:16])
    defparam i1_4_lut_adj_978.LUT_INIT = 16'hcecc;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\FRAME_MATCHER.state [4]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29015));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_980 (.I0(\FRAME_MATCHER.state [4]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29109));
    defparam i1_2_lut_adj_980.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\FRAME_MATCHER.state [5]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29013));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_982 (.I0(\FRAME_MATCHER.state [5]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29111));
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_983 (.I0(\FRAME_MATCHER.state [6]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29011));
    defparam i1_2_lut_adj_983.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\FRAME_MATCHER.state [6]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29113));
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\FRAME_MATCHER.state [7]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29009));
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_986 (.I0(\FRAME_MATCHER.state [7]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29115));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_987 (.I0(\FRAME_MATCHER.state [8]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29007));
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\FRAME_MATCHER.state [8]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29117));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_989 (.I0(\FRAME_MATCHER.state [9]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29005));
    defparam i1_2_lut_adj_989.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_990 (.I0(\FRAME_MATCHER.state [9]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29119));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_991 (.I0(\FRAME_MATCHER.state [10]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29003));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_992 (.I0(\FRAME_MATCHER.state [10]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29121));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\FRAME_MATCHER.state [11]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29001));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_994 (.I0(\FRAME_MATCHER.state [11]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29123));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\FRAME_MATCHER.state [12]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28999));
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_996 (.I0(\FRAME_MATCHER.state [12]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29125));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_997 (.I0(\FRAME_MATCHER.state [13]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3664));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_998 (.I0(\FRAME_MATCHER.state [14]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3665));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_999 (.I0(\FRAME_MATCHER.state [15]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28997));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1000 (.I0(\FRAME_MATCHER.state [15]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29127));
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\FRAME_MATCHER.state [16]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28995));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1002 (.I0(\FRAME_MATCHER.state [16]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29129));
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1003 (.I0(\FRAME_MATCHER.state [17]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29017));
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(\FRAME_MATCHER.state [17]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29107));
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\FRAME_MATCHER.state [18]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28993));
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(\FRAME_MATCHER.state [18]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29131));
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\FRAME_MATCHER.state [19]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28991));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(\FRAME_MATCHER.state [19]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29133));
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(\FRAME_MATCHER.state [20]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28989));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(\FRAME_MATCHER.state [20]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29135));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(\FRAME_MATCHER.state [21]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28987));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(\FRAME_MATCHER.state [21]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29137));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\FRAME_MATCHER.state [22]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28985));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(\FRAME_MATCHER.state [22]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29139));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\FRAME_MATCHER.state [23]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28983));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(\FRAME_MATCHER.state [23]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29141));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(\FRAME_MATCHER.state [24]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28981));
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\FRAME_MATCHER.state [24]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29143));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(\FRAME_MATCHER.state [25]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28979));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(\FRAME_MATCHER.state [25]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29145));
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(\FRAME_MATCHER.state [26]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28977));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h8888;
    SB_LUT4 mux_987_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19] [6]), .O(n4022));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(\FRAME_MATCHER.state [26]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29147));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\FRAME_MATCHER.state [27]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28975));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(\FRAME_MATCHER.state [27]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29149));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\FRAME_MATCHER.state [28]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28949));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\FRAME_MATCHER.state [28]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29151));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\FRAME_MATCHER.state [29]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28973));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\FRAME_MATCHER.state [29]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29153));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\FRAME_MATCHER.state [30]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n28971));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\FRAME_MATCHER.state [30]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29155));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\FRAME_MATCHER.i [4]), .I1(n15542), .I2(GND_net), 
            .I3(GND_net), .O(n15459));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'heeee;
    SB_LUT4 i17139_4_lut (.I0(n5_adj_3666), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i17139_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i7_4_lut_adj_1032 (.I0(n29584), .I1(n14_adj_3667), .I2(n10_adj_3668), 
            .I3(\data_out_frame[23] [4]), .O(n30142));
    defparam i7_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i17147_4_lut (.I0(n8_adj_3669), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n15459), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i17147_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_3_lut_adj_1033 (.I0(\FRAME_MATCHER.i_31__N_2364 ), .I1(n771), 
            .I2(n12869), .I3(GND_net), .O(n67));
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'h2020;
    SB_LUT4 i123_3_lut (.I0(\FRAME_MATCHER.i_31__N_2368 ), .I1(n3303), .I2(n12869), 
            .I3(GND_net), .O(n117));   // verilog/coms.v(115[11:12])
    defparam i123_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i27531_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n16_adj_3670), 
            .I2(n6_adj_3671), .I3(GND_net), .O(n33102));   // verilog/coms.v(112[11:16])
    defparam i27531_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n1733), .I1(n33102), .I2(n89), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n2329));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h0544;
    SB_LUT4 i121_2_lut (.I0(n12869), .I1(n2329), .I2(GND_net), .I3(GND_net), 
            .O(n115));
    defparam i121_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28532_2_lut (.I0(byte_transmit_counter[7]), .I1(n4_adj_3672), 
            .I2(GND_net), .I3(GND_net), .O(tx_transmit_N_3257));
    defparam i28532_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i18_4_lut_adj_1035 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_3673));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut_adj_1035.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1036 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_3674));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut_adj_1036.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1037 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_3675));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut_adj_1037.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1038 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43_adj_3675), .I2(n42_adj_3674), 
            .I3(n44_adj_3673), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1039 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45_adj_3676));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1040 (.I0(n45_adj_3676), .I1(n50), .I2(n39), 
            .I3(n40), .O(n15542));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i2820_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3677));
    defparam i2820_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17149_4_lut (.I0(n8_adj_3678), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n15542), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i17149_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i5_3_lut_adj_1041 (.I0(\data_in[0] [3]), .I1(\data_in[2] [4]), 
            .I2(\data_in[3] [0]), .I3(GND_net), .O(n14_adj_3679));
    defparam i5_3_lut_adj_1041.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1042 (.I0(\data_in[1] [4]), .I1(\data_in[0] [6]), 
            .I2(n15610), .I3(\data_in[1] [5]), .O(n15_adj_3680));
    defparam i6_4_lut_adj_1042.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1043 (.I0(n15_adj_3680), .I1(\data_in[1] [0]), 
            .I2(n14_adj_3679), .I3(\data_in[2] [2]), .O(n15462));
    defparam i8_4_lut_adj_1043.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1044 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_3681));
    defparam i6_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1045 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_3682));
    defparam i7_4_lut_adj_1045.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1046 (.I0(n17_adj_3682), .I1(\data_in[1] [6]), 
            .I2(n16_adj_3681), .I3(\data_in[3] [7]), .O(n15539));
    defparam i9_4_lut_adj_1046.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_adj_1047 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n31109));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1047.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1048 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3683));
    defparam i4_4_lut_adj_1048.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1049 (.I0(\data_in[3] [4]), .I1(n10_adj_3683), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n15610));
    defparam i5_3_lut_adj_1049.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3684));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1050 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3685));
    defparam i6_4_lut_adj_1050.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1051 (.I0(\data_in[3] [6]), .I1(n14_adj_3685), 
            .I2(n10_adj_3684), .I3(\data_in[2] [1]), .O(n15583));
    defparam i7_4_lut_adj_1051.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1052 (.I0(\data_in[2] [4]), .I1(n15583), .I2(\data_in[1] [5]), 
            .I3(n15610), .O(n18_adj_3686));
    defparam i7_4_lut_adj_1052.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1053 (.I0(\data_in[0] [6]), .I1(n18_adj_3686), 
            .I2(\data_in[3] [0]), .I3(n15539), .O(n20_adj_3687));
    defparam i9_4_lut_adj_1053.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3688));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1054 (.I0(n15_adj_3688), .I1(n20_adj_3687), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_3689));
    defparam i10_4_lut_adj_1054.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1055 (.I0(n15462), .I1(\data_in[0] [7]), .I2(\data_in[2] [1]), 
            .I3(\data_in[3] [6]), .O(n16_adj_3690));
    defparam i6_4_lut_adj_1055.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1056 (.I0(n15539), .I1(\data_in[0] [2]), .I2(\data_in[3] [3]), 
            .I3(\data_in[3] [1]), .O(n17_adj_3691));
    defparam i7_4_lut_adj_1056.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1057 (.I0(n17_adj_3691), .I1(\data_in[2] [3]), 
            .I2(n16_adj_3690), .I3(\data_in[3] [5]), .O(n63_adj_3692));
    defparam i9_4_lut_adj_1057.LUT_INIT = 16'hfbff;
    SB_LUT4 i8_4_lut_adj_1058 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n15583), .I3(\data_in[0] [1]), .O(n20_adj_3693));
    defparam i8_4_lut_adj_1058.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1059 (.I0(n15462), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_3694));
    defparam i7_4_lut_adj_1059.LUT_INIT = 16'hfeff;
    SB_LUT4 i26590_4_lut (.I0(\data_in[1] [3]), .I1(\data_in[0] [5]), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [2]), .O(n32264));
    defparam i26590_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n32264), .I1(n19_adj_3694), .I2(n20_adj_3693), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_3_lut_adj_1060 (.I0(\FRAME_MATCHER.i_31__N_2370 ), .I1(n4452), 
            .I2(n12869), .I3(GND_net), .O(n2_adj_3695));
    defparam i1_3_lut_adj_1060.LUT_INIT = 16'h2020;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(n884), .I1(n2_adj_3695), .I2(\FRAME_MATCHER.i_31__N_2367 ), 
            .I3(n12869), .O(n4_c));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\FRAME_MATCHER.state [31]), .I1(n5_adj_3663), 
            .I2(GND_net), .I3(GND_net), .O(n29019));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(\FRAME_MATCHER.state [31]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n29105));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n16917));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3696));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3697));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_987_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19] [7]), .O(n4023));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(\FRAME_MATCHER.state[0] ), .I1(n23888), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2367 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n16916));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n16915));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i17_2_lut (.I0(PWMLimit[14]), .I1(\duty_23__N_3516[14] ), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(4[26:30])
    defparam i17_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n16914));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_24_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n24885), .O(n2_adj_3698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n24885), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n24886));
    SB_LUT4 i12859_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n16968));
    defparam i12859_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_987_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n4024));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i24688_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n30352));
    defparam i24688_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i17033_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3360[0]), .I2(GND_net), 
            .I3(GND_net), .O(n21130));
    defparam i17033_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n29513));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n114));   // verilog/coms.v(112[11:16])
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1067 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_3700));
    defparam i1_4_lut_adj_1067.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_1068 (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[3]), 
            .I2(byte_transmit_counter[6]), .I3(n4_adj_3700), .O(n4_adj_3672));
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'hfefa;
    SB_LUT4 i2_4_lut_adj_1069 (.I0(\FRAME_MATCHER.state[0] ), .I1(n22109), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(n114), .O(n31265));
    defparam i2_4_lut_adj_1069.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut_adj_1070 (.I0(n29513), .I1(n21130), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(byte_transmit_counter[7]), .O(n10_adj_3701));
    defparam i4_4_lut_adj_1070.LUT_INIT = 16'h0020;
    SB_LUT4 i1_3_lut_adj_1071 (.I0(n4_adj_3672), .I1(n16695), .I2(n10_adj_3701), 
            .I3(GND_net), .O(n2863[0]));
    defparam i1_3_lut_adj_1071.LUT_INIT = 16'hdcdc;
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n16913));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i27789_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33187));
    defparam i27789_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27813_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33186));
    defparam i27813_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_987_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n4025));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n4026));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n4027));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n4028));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n16912));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3360[0]), .C(clk32MHz), 
            .D(n2863[0]), .R(n31265));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1072 (.I0(\FRAME_MATCHER.state [6]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n21855));
    defparam i3_4_lut_adj_1072.LUT_INIT = 16'hfffe;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n16911));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_23_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n24884), .O(n2_adj_3702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n16652), .D(n8825[7]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n16910));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1073 (.I0(\FRAME_MATCHER.state [24]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [17]), .I3(\FRAME_MATCHER.state [22]), 
            .O(n16_adj_3703));   // verilog/coms.v(127[12] 300[6])
    defparam i6_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n16909));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_987_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n4029));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1074 (.I0(n31109), .I1(n29726), .I2(Kp_23__N_764), 
            .I3(\data_in_frame[4] [5]), .O(n10_adj_3704));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1075 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [18]), 
            .I2(\FRAME_MATCHER.state [25]), .I3(\FRAME_MATCHER.state [20]), 
            .O(n17_adj_3705));   // verilog/coms.v(127[12] 300[6])
    defparam i7_4_lut_adj_1075.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1076 (.I0(n16245), .I1(\data_in_frame[2] [6]), 
            .I2(\data_in_frame[7] [2]), .I3(\data_in_frame[4] [6]), .O(n12_adj_3706));
    defparam i5_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1077 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [31]), 
            .I2(\FRAME_MATCHER.state [13]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n22_adj_3707));
    defparam i8_4_lut_adj_1077.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1078 (.I0(n16604), .I1(n12_adj_3706), .I2(n29905), 
            .I3(n16107), .O(n16329));
    defparam i6_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1079 (.I0(\FRAME_MATCHER.state [28]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(\FRAME_MATCHER.state [14]), .I3(\FRAME_MATCHER.state [9]), 
            .O(n24_adj_3708));
    defparam i10_4_lut_adj_1079.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1080 (.I0(\data_in_frame[1] [7]), .I1(n30011), 
            .I2(\data_in_frame[6] [1]), .I3(\data_in_frame[2] [0]), .O(n12_adj_3709));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1081 (.I0(\FRAME_MATCHER.state [11]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(\FRAME_MATCHER.state [10]), .I3(\FRAME_MATCHER.state [29]), 
            .O(n23));
    defparam i9_4_lut_adj_1081.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1082 (.I0(\data_in_frame[8] [3]), .I1(n12_adj_3709), 
            .I2(n30173), .I3(\data_in_frame[6] [2]), .O(n15905));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1083 (.I0(n17_adj_3705), .I1(\FRAME_MATCHER.state [19]), 
            .I2(n16_adj_3703), .I3(\FRAME_MATCHER.state [26]), .O(n27783));   // verilog/coms.v(127[12] 300[6])
    defparam i9_4_lut_adj_1083.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n29635));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h6666;
    SB_LUT4 i11_3_lut_adj_1085 (.I0(\FRAME_MATCHER.state [23]), .I1(n22_adj_3707), 
            .I2(\FRAME_MATCHER.state [12]), .I3(GND_net), .O(n25));
    defparam i11_3_lut_adj_1085.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n15856));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1087 (.I0(n25), .I1(n27783), .I2(n23), .I3(n24_adj_3708), 
            .O(n23828));
    defparam i1_4_lut_adj_1087.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1088 (.I0(n1), .I1(n23888), .I2(n29447), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n4218));
    defparam i3_4_lut_adj_1088.LUT_INIT = 16'h0040;
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n16908));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_987_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n4030));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n16907));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_987_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n4031));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[17] [0]), .O(n4032));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n16652), .D(n8825[6]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3710));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3711));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_987_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[17] [1]), .O(n4033));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[17] [2]), .O(n4034));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[17] [3]), .O(n4035));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i27794_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33170));
    defparam i27794_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27796_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33169));
    defparam i27796_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_987_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n4036));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17] [5]), .O(n4037));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[17] [6]), .O(n4038));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12860_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n16969));
    defparam i12860_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3712));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3713));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_987_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17] [7]), .O(n4039));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_987_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n4016));   // verilog/coms.v(127[12] 300[6])
    defparam mux_987_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12891_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n17000));
    defparam i12891_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12892_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[6]), 
            .I3(\data_in_frame[9]_c [6]), .O(n17001));
    defparam i12892_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12893_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[5]), 
            .I3(\data_in_frame[9][5] ), .O(n17002));
    defparam i12893_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n29105), .S(n29019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n29155), .S(n28971));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n29153), .S(n28973));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n29151), .S(n28949));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n29149), .S(n28975));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n29147), .S(n28977));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n29145), .S(n28979));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n29143), .S(n28981));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n29141), .S(n28983));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n29139), .S(n28985));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n29137), .S(n28987));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n29135), .S(n28989));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n29133), .S(n28991));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n29131), .S(n28993));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n29107), .S(n29017));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n29129), .S(n28995));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n29127), .S(n28997));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n7_adj_3665), .S(n8_adj_3714));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n7_adj_3664), .S(n8_adj_3715));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n29125), .S(n28999));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n29123), .S(n29001));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n29121), .S(n29003));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n29119), .S(n29005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n29117), .S(n29007));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n29115), .S(n29009));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n29113), .S(n29011));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n29111), .S(n29013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n29109), .S(n29015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n28941), .S(n29199));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n28947), .S(n34932));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n16652), .D(n8825[5]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_23 (.CI(n24884), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n24885));
    SB_LUT4 i12894_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[4]), 
            .I3(\data_in_frame[9][4] ), .O(n17003));
    defparam i12894_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_22_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n24883), .O(n2_adj_3716)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1089 (.I0(\FRAME_MATCHER.state_31__N_2468 [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n92), .I3(\FRAME_MATCHER.state[2] ), .O(n32156));
    defparam i3_4_lut_adj_1089.LUT_INIT = 16'h0040;
    SB_CARRY add_43_22 (.CI(n24883), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n24884));
    SB_LUT4 add_43_21_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n24882), .O(n2_adj_3717)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12895_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[3]), 
            .I3(\data_in_frame[9][3] ), .O(n17004));
    defparam i12895_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12896_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[2]), 
            .I3(\data_in_frame[9][2] ), .O(n17005));
    defparam i12896_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n16652), .D(n8825[4]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n16652), .D(n8825[3]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n16652), .D(n8825[2]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n16652), .D(n8825[1]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n16695), .D(n29913));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28645_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n32156), .I2(n32159), 
            .I3(n6_adj_3671), .O(n31247));
    defparam i28645_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i12897_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[1]), 
            .I3(\data_in_frame[9][1] ), .O(n17006));
    defparam i12897_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12898_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29555), .I2(rx_data[0]), 
            .I3(\data_in_frame[9][0] ), .O(n17007));
    defparam i12898_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[19] [3]), .I3(GND_net), .O(n6_adj_3612));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1090 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[19] [2]), 
            .I2(n16479), .I3(GND_net), .O(n6_adj_3656));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1090.LUT_INIT = 16'h9696;
    SB_CARRY add_43_21 (.CI(n24882), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n24883));
    SB_LUT4 add_43_20_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n24881), .O(n2_adj_3718)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n24881), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n24882));
    SB_LUT4 i5_3_lut_4_lut (.I0(n26989), .I1(\data_out_frame[19] [3]), .I2(\data_out_frame[17] [1]), 
            .I3(n10_adj_3719), .O(n27954));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_19_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n24880), .O(n2_adj_3720)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_19 (.CI(n24880), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n24881));
    SB_LUT4 add_43_18_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n24879), .O(n2_adj_3721)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[10] [1]), .I3(\data_out_frame[10] [2]), 
            .O(n30234));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n16695), .D(n31807));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n16695), .D(n31034));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n16695), .D(n31430));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n16695), .D(n30150));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n16695), .D(n31438));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n16695), .D(n31868));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n16695), .D(n30501));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n16695), .D(n31011));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n16695), .D(n31372));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n16695), .D(n29835));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n16695), .D(n31099));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n16695), .D(n16060));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n16695), .D(n31955));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n16695), .D(n30676));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n16695), .D(n30802));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3722), .S(n3_adj_3723));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_18 (.CI(n24879), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n24880));
    SB_LUT4 add_43_17_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n24878), .O(n2_adj_3724)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3725), .S(n3_adj_3726));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3727), .S(n3_adj_3728));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3729), .S(n3_adj_3730));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3731), .S(n3_adj_3732));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3733), .S(n3_adj_3734));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3735), .S(n3_adj_3736));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3737), .S(n3_adj_3738));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3739), .S(n3_adj_3740));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3698), .S(n3_adj_3741));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3702), .S(n3_adj_3742));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3716), .S(n3_adj_3743));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3717), .S(n3_adj_3744));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3718), .S(n3_adj_3745));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3720), .S(n3_adj_3746));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3721), .S(n3_adj_3747));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3724), .S(n3_adj_3748));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3749), .S(n3_adj_3750));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3751), .S(n3_adj_3752));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3753), .S(n3_adj_3754));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3755), .S(n3_adj_3756));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3757), .S(n3_adj_3758));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3759), .S(n3_adj_3760));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3761), .S(n3_adj_3762));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3763), .S(n3_adj_3764));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3765), .S(n3_adj_3766));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3767), .S(n3_adj_3768));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3769), .S(n3_adj_3770));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3771), .S(n3_adj_3772));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3773), .S(n3_adj_3774));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3775), .S(n3_adj_3776));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n16631), 
            .D(n4039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n16906));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1091 (.I0(n18487), .I1(n23828), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3777));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h2222;
    SB_LUT4 i27798_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33167));
    defparam i27798_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27800_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33166));
    defparam i27800_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1092 (.I0(\FRAME_MATCHER.state[2] ), .I1(n21855), 
            .I2(n30352), .I3(n6_adj_3777), .O(n16631));
    defparam i4_4_lut_adj_1092.LUT_INIT = 16'h0200;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1093 (.I0(n21151), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n29530));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1093.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(n23828), .I1(n21855), .I2(GND_net), 
            .I3(GND_net), .O(n22109));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\FRAME_MATCHER.state[3] ), .I1(n78), 
            .I2(GND_net), .I3(GND_net), .O(n18751));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1096 (.I0(\FRAME_MATCHER.i_31__N_2368 ), .I1(n31275), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n1733));
    defparam i2_3_lut_adj_1096.LUT_INIT = 16'hbaba;
    SB_LUT4 i2_3_lut_4_lut_adj_1097 (.I0(\data_out_frame[18] [7]), .I1(n29980), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[17] [1]), 
            .O(n29946));
    defparam i2_3_lut_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1098 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[12] [0]), 
            .I2(\data_out_frame[11] [5]), .I3(GND_net), .O(n6_adj_3617));
    defparam i1_2_lut_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[12] [0]), 
            .I2(n27050), .I3(GND_net), .O(n10_adj_3645));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n16631), 
            .D(n4038));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_17 (.CI(n24878), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n24879));
    SB_LUT4 add_43_16_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n24877), .O(n2_adj_3749)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1099 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n15751));
    defparam i1_2_lut_3_lut_adj_1099.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1100 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n6_adj_3606));
    defparam i1_2_lut_3_lut_adj_1100.LUT_INIT = 16'h9696;
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n16631), 
            .D(n4037));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n16631), 
            .D(n4036));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n16631), 
            .D(n4035));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n16631), 
            .D(n4034));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n16631), 
            .D(n4033));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n16631), 
            .D(n4032));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n16631), 
            .D(n4031));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n16631), 
            .D(n4030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n16905));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n16631), 
            .D(n4029));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n16631), 
            .D(n4028));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n16631), 
            .D(n4027));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n16631), 
            .D(n4026));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n16631), .D(n4025));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n16631), .D(n4024));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n16631), .D(n4023));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n16631), .D(n4022));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n16631), .D(n4021));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n16631), .D(n4020));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n16631), .D(n4019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n16631), .D(n4018));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n16631), .D(n4017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n16904));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_16 (.CI(n24877), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n24878));
    SB_LUT4 add_43_15_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n24876), .O(n2_adj_3751)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n16903));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n16902));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1101 (.I0(n15811), .I1(n16220), .I2(\data_in_frame[7] [5]), 
            .I3(n29971), .O(n10_adj_3778));
    defparam i4_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1102 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[13] [6]), .I3(GND_net), .O(n10_adj_3607));
    defparam i2_2_lut_3_lut_adj_1102.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1103 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[11] [6]), .I3(GND_net), .O(n29993));
    defparam i1_2_lut_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i12883_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n16992));
    defparam i12883_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_15 (.CI(n24876), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n24877));
    SB_LUT4 i12884_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n16993));
    defparam i12884_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12885_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n16994));
    defparam i12885_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_14_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n24875), .O(n2_adj_3753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_3_lut_adj_1104 (.I0(n16493), .I1(n10_adj_3778), .I2(\data_in_frame[5] [4]), 
            .I3(GND_net), .O(n16094));
    defparam i5_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i12886_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n16995));
    defparam i12886_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n16901));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1105 (.I0(\data_in_frame[15] [6]), .I1(n27936), 
            .I2(n29609), .I3(n6_adj_3779), .O(n29984));
    defparam i4_4_lut_adj_1105.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(n27918), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30231));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1107 (.I0(n16445), .I1(n29767), .I2(n29609), 
            .I3(n29797), .O(n18_adj_3780));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1108 (.I0(n29771), .I1(n18_adj_3780), .I2(\data_in_frame[18] [3]), 
            .I3(n29884), .O(n20_adj_3781));   // verilog/coms.v(74[16:43])
    defparam i9_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1109 (.I0(\data_in_frame[13] [7]), .I1(n20_adj_3781), 
            .I2(n16445), .I3(\data_in_frame[15] [7]), .O(n29930));   // verilog/coms.v(74[16:43])
    defparam i10_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_15__7__I_0_3897_2_lut (.I0(\data_in_frame[15] [7]), 
            .I1(\data_in_frame[15] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1261));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_15__7__I_0_3897_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30246));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n29771));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30039));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i4_2_lut_adj_1113 (.I0(\data_in_frame[16] [4]), .I1(n30067), 
            .I2(GND_net), .I3(GND_net), .O(n42_adj_3782));   // verilog/coms.v(74[16:43])
    defparam i4_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_LUT4 i22_4_lut (.I0(n29604), .I1(\data_in_frame[12] [0]), .I2(\data_in_frame[16] [5]), 
            .I3(\data_in_frame[14] [7]), .O(n60));   // verilog/coms.v(74[16:43])
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1114 (.I0(n30039), .I1(n29771), .I2(n27918), 
            .I3(n30246), .O(n58));   // verilog/coms.v(74[16:43])
    defparam i20_4_lut_adj_1114.LUT_INIT = 16'h9669;
    SB_LUT4 i30_4_lut (.I0(\data_in_frame[14] [1]), .I1(n60), .I2(n42_adj_3782), 
            .I3(\data_in_frame[14] [3]), .O(n68));   // verilog/coms.v(74[16:43])
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[15] [4]), .I3(\data_in_frame[10] [6]), .O(n64));   // verilog/coms.v(74[16:43])
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1115 (.I0(n29870), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[16] [2]), .I3(\data_in_frame[16] [6]), .O(n62));   // verilog/coms.v(74[16:43])
    defparam i24_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1116 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[14] [2]), .I3(Kp_23__N_1261), .O(n63_adj_3783));   // verilog/coms.v(74[16:43])
    defparam i25_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(\data_in_frame[16] [3]), .I1(n30192), .I2(n30255), 
            .I3(n30051), .O(n61));   // verilog/coms.v(74[16:43])
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n30090), .I1(n29666), .I2(n29711), .I3(n15714), 
            .O(n66));   // verilog/coms.v(74[16:43])
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34_4_lut (.I0(\data_in_frame[10]_c [2]), .I1(n68), .I2(n58), 
            .I3(n34034), .O(n72));   // verilog/coms.v(74[16:43])
    defparam i34_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i27_4_lut (.I0(n30201), .I1(n15951), .I2(n29672), .I3(\data_in_frame[11] [5]), 
            .O(n65));   // verilog/coms.v(74[16:43])
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35_4_lut (.I0(n61), .I1(n63_adj_3783), .I2(n62), .I3(n64), 
            .O(n73));   // verilog/coms.v(74[16:43])
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i37_4_lut (.I0(n73), .I1(n65), .I2(n72), .I3(n66), .O(n31528));   // verilog/coms.v(74[16:43])
    defparam i37_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut (.I0(n30249), .I1(\data_in_frame[18] [2]), .I2(n29930), 
            .I3(GND_net), .O(n16_adj_3784));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1117 (.I0(n30130), .I1(n27106), .I2(\data_in_frame[17] [7]), 
            .I3(n30231), .O(n19_adj_3785));
    defparam i7_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1118 (.I0(n19_adj_3785), .I1(n29927), .I2(n16_adj_3784), 
            .I3(n31528), .O(n22_adj_3786));
    defparam i10_4_lut_adj_1118.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1119 (.I0(n17_adj_3787), .I1(n22_adj_3786), .I2(\data_in_frame[18] [1]), 
            .I3(n27633), .O(n30807));
    defparam i11_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1120 (.I0(n30249), .I1(n30530), .I2(\data_in_frame[19] [0]), 
            .I3(n30258), .O(n10_adj_3788));
    defparam i4_4_lut_adj_1120.LUT_INIT = 16'h9669;
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n16900));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_adj_1121 (.I0(n30195), .I1(n10_adj_3788), .I2(\data_in_frame[18] [7]), 
            .I3(GND_net), .O(n27550));
    defparam i5_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1122 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n29707));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1123 (.I0(n15768), .I1(n30179), .I2(n27986), 
            .I3(Kp_23__N_1054), .O(n29672));
    defparam i3_4_lut_adj_1123.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1124 (.I0(Kp_23__N_1026), .I1(n15918), .I2(n30023), 
            .I3(n29672), .O(n10_adj_3789));
    defparam i4_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_adj_1125 (.I0(Kp_23__N_1035), .I1(n16094), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i3_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1126 (.I0(\data_in_frame[11] [1]), .I1(n9), .I2(\data_in_frame[10] [7]), 
            .I3(n10_adj_3789), .O(n29848));
    defparam i2_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1127 (.I0(n15777), .I1(\data_in_frame[9][2] ), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n29717));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1128 (.I0(n26977), .I1(Kp_23__N_1050), .I2(n30111), 
            .I3(n15777), .O(n14_adj_3790));
    defparam i6_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1129 (.I0(\data_in_frame[13] [3]), .I1(n29848), 
            .I2(n15947), .I3(n15643), .O(n13_adj_3791));
    defparam i5_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n16899));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_adj_1130 (.I0(\data_in_frame[15] [5]), .I1(n13_adj_3791), 
            .I2(n14_adj_3790), .I3(GND_net), .O(n27918));
    defparam i1_3_lut_adj_1130.LUT_INIT = 16'h6969;
    SB_LUT4 i5_3_lut_adj_1131 (.I0(\data_in_frame[17] [7]), .I1(n27918), 
            .I2(n29717), .I3(GND_net), .O(n14_adj_3792));
    defparam i5_3_lut_adj_1131.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1132 (.I0(n30114), .I1(\data_in_frame[16] [1]), 
            .I2(n26977), .I3(n29797), .O(n15_adj_3793));
    defparam i6_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1133 (.I0(n15_adj_3793), .I1(n29707), .I2(n14_adj_3792), 
            .I3(n16445), .O(n30213));
    defparam i8_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1134 (.I0(\FRAME_MATCHER.state_31__N_2468 [3]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n22109), .I3(n6_adj_3794), .O(n12944));
    defparam i4_4_lut_adj_1134.LUT_INIT = 16'h0200;
    SB_LUT4 i2_3_lut_adj_1135 (.I0(n16011), .I1(\data_in_frame[9][5] ), 
            .I2(n15918), .I3(GND_net), .O(n27061));
    defparam i2_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1136 (.I0(\data_in_frame[14] [0]), .I1(n29767), 
            .I2(\data_in_frame[11] [6]), .I3(n27061), .O(n27936));
    defparam i1_4_lut_adj_1136.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1137 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30084));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[11] [5]), .I1(n27936), 
            .I2(GND_net), .I3(GND_net), .O(n29797));
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1139 (.I0(n29971), .I1(n30145), .I2(\data_in_frame[5] [2]), 
            .I3(n29726), .O(n12_adj_3795));
    defparam i5_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut_adj_1140 (.I0(n27008), .I1(n30219), .I2(n29666), 
            .I3(GND_net), .O(n11));
    defparam i4_3_lut_adj_1140.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1141 (.I0(Kp_23__N_1035), .I1(n11), .I2(n16353), 
            .I3(n12_adj_3795), .O(n10_adj_3796));
    defparam i2_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1142 (.I0(n16204), .I1(n28008), .I2(\data_in_frame[11] [7]), 
            .I3(\data_in_frame[9] [7]), .O(n14_adj_3797));
    defparam i6_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1143 (.I0(\data_in_frame[14] [2]), .I1(n9_adj_3798), 
            .I2(n14_adj_3797), .I3(n10_adj_3796), .O(n29698));
    defparam i1_4_lut_adj_1143.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1144 (.I0(n29797), .I1(n30084), .I2(n16333), 
            .I3(\data_in_frame[9][3] ), .O(n12_adj_3799));
    defparam i5_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1145 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[14] [1]), 
            .I2(n12_adj_3799), .I3(n8_adj_3800), .O(n29884));
    defparam i1_4_lut_adj_1145.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1146 (.I0(n29928), .I1(n27683), .I2(GND_net), 
            .I3(GND_net), .O(n27944));
    defparam i1_2_lut_adj_1146.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_in_frame[9][1] ), .I1(\data_in_frame[9][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n15714));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_in_frame[9][3] ), .I1(\data_in_frame[9][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n15643));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1149 (.I0(n27986), .I1(n30179), .I2(n30023), 
            .I3(n29959), .O(n28008));
    defparam i3_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1150 (.I0(n16204), .I1(Kp_23__N_1050), .I2(\data_in_frame[9][5] ), 
            .I3(GND_net), .O(n29813));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1150.LUT_INIT = 16'h9696;
    SB_LUT4 i12887_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n16996));
    defparam i12887_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[9][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n29754));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1152 (.I0(n16094), .I1(n29813), .I2(n28008), 
            .I3(GND_net), .O(Kp_23__N_1035));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1152.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1153 (.I0(\data_in_frame[8] [0]), .I1(n15866), 
            .I2(n29744), .I3(n6_adj_3801), .O(n31643));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1154 (.I0(n7_adj_3802), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[6] [3]), .I3(\data_in_frame[9]_c [6]), .O(n24_adj_3803));
    defparam i10_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1155 (.I0(\data_in_frame[9][0] ), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[4] [2]), .I3(Kp_23__N_1035), .O(n22_adj_3804));
    defparam i8_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1156 (.I0(n16353), .I1(\data_in_frame[8] [4]), 
            .I2(n29754), .I3(\data_in_frame[8] [2]), .O(n23_adj_3805));
    defparam i9_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1157 (.I0(\data_in_frame[7] [7]), .I1(n31643), 
            .I2(n29787), .I3(n30081), .O(n21));
    defparam i7_4_lut_adj_1157.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1158 (.I0(n21), .I1(n23_adj_3805), .I2(n22_adj_3804), 
            .I3(n24_adj_3803), .O(n30145));
    defparam i13_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[9][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n29790));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1160 (.I0(n29790), .I1(\data_in_frame[13] [7]), 
            .I2(n30228), .I3(n6_adj_3806), .O(n26998));
    defparam i4_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1161 (.I0(n29884), .I1(n26998), .I2(\data_in_frame[16] [3]), 
            .I3(n29698), .O(n27940));
    defparam i3_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1162 (.I0(n16098), .I1(Kp_23__N_605), .I2(n27944), 
            .I3(n29881), .O(n10_adj_3807));
    defparam i4_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1163 (.I0(n27940), .I1(n10_adj_3807), .I2(n27402), 
            .I3(GND_net), .O(n29878));
    defparam i5_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1164 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[19] [3]), .O(n8_adj_3808));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1165 (.I0(\data_in_frame[19] [4]), .I1(n8_adj_3808), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[19] [5]), .O(Kp_23__N_605));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_in_frame[9][5] ), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n29764));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(\data_in_frame[12] [1]), .I1(n16011), 
            .I2(GND_net), .I3(GND_net), .O(n30186));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1168 (.I0(\data_out_frame[25] [6]), .I1(n29825), 
            .I2(\data_out_frame[23] [4]), .I3(n2128), .O(n30802));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1169 (.I0(\data_out_frame[23] [6]), .I1(n27954), 
            .I2(\data_out_frame[25] [7]), .I3(n29839), .O(n29825));
    defparam i3_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1170 (.I0(n30020), .I1(n29825), .I2(n29910), 
            .I3(\data_out_frame[24] [5]), .O(n34));
    defparam i13_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1171 (.I0(\data_in_frame[12] [2]), .I1(n30186), 
            .I2(\data_in_frame[10][1] ), .I3(n29764), .O(n12_adj_3809));
    defparam i5_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1172 (.I0(\data_in_frame[9]_c [6]), .I1(n12_adj_3809), 
            .I2(\data_in_frame[14] [3]), .I3(n30036), .O(n29915));
    defparam i6_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1173 (.I0(\data_in_frame[18] [7]), .I1(n16368), 
            .I2(\data_in_frame[16] [6]), .I3(n4_adj_3810), .O(n30130));
    defparam i2_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1174 (.I0(\data_in_frame[16] [5]), .I1(n30216), 
            .I2(n30130), .I3(n29915), .O(n28034));
    defparam i3_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9]_c [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1050));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n2329), .I1(n2), .I2(n33[1]), .I3(n63), 
            .O(n28947));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'he0ee;
    SB_LUT4 i28358_2_lut (.I0(n16353), .I1(\data_in_frame[10]_c [0]), .I2(GND_net), 
            .I3(GND_net), .O(n34034));   // verilog/coms.v(96[12:25])
    defparam i28358_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1175 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[12] [2]), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n30051));   // verilog/coms.v(96[12:25])
    defparam i2_3_lut_adj_1175.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1176 (.I0(n29736), .I1(n30051), .I2(n34034), 
            .I3(GND_net), .O(n27106));   // verilog/coms.v(96[12:25])
    defparam i2_3_lut_adj_1176.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1177 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[9] [7]), 
            .I2(n30183), .I3(n14041), .O(n10_adj_3812));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1178 (.I0(n31275), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n4452), .O(n29497));
    defparam i1_2_lut_3_lut_4_lut_adj_1178.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(n16094), .I1(\data_in_frame[10][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n29711));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n29870));
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1181 (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n78), .I3(n63_adj_3), .O(n16_adj_3670));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1181.LUT_INIT = 16'hfd00;
    SB_LUT4 i1_2_lut_adj_1182 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16267));
    defparam i1_2_lut_adj_1182.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1183 (.I0(n16280), .I1(n29598), .I2(\data_in_frame[6] [0]), 
            .I3(\data_in_frame[7] [7]), .O(n14041));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1184 (.I0(n1733), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n8_adj_3813), .O(n29546));
    defparam i1_2_lut_3_lut_4_lut_adj_1184.LUT_INIT = 16'hfff7;
    SB_LUT4 i17_4_lut_adj_1185 (.I0(\data_out_frame[23] [5]), .I1(n34), 
            .I2(n24_adj_3814), .I3(n29952), .O(n38));
    defparam i17_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1186 (.I0(n29946), .I1(n29834), .I2(n29857), 
            .I3(n29723), .O(n36_adj_3815));
    defparam i15_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1187 (.I0(n117), .I1(n67), .I2(n12869), 
            .I3(n2329), .O(n5_adj_3663));
    defparam i1_2_lut_3_lut_4_lut_adj_1187.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(\data_in_frame[10] [3]), .I1(n14048), 
            .I2(GND_net), .I3(GND_net), .O(n15941));
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1189 (.I0(n30070), .I1(n29736), .I2(n15941), 
            .I3(n6_adj_3816), .O(n30195));
    defparam i4_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[16] [6]), .I1(n30195), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3817));
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1191 (.I0(\data_in_frame[16] [7]), .I1(n27106), 
            .I2(n29784), .I3(n6_adj_3817), .O(n30530));
    defparam i4_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(n30530), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30216));
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1193 (.I0(\data_in_frame[17] [1]), .I1(n30258), 
            .I2(n16267), .I3(n30067), .O(n10_adj_3818));
    defparam i4_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1194 (.I0(n1733), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n8_adj_3819), .O(n29549));
    defparam i1_2_lut_3_lut_4_lut_adj_1194.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1195 (.I0(n1733), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n8_adj_3820), .O(n29555));
    defparam i1_2_lut_3_lut_4_lut_adj_1195.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[19] [1]), .I1(n28034), 
            .I2(GND_net), .I3(GND_net), .O(n29924));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h9999;
    SB_LUT4 i2_2_lut_adj_1197 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3821));
    defparam i2_2_lut_adj_1197.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(n15905), .I1(n15951), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1026));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1199 (.I0(\data_in_frame[15] [2]), .I1(n29663), 
            .I2(\data_in_frame[15] [3]), .I3(\data_in_frame[13] [2]), .O(n29604));
    defparam i3_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1200 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[10] [4]), .I3(GND_net), .O(n30090));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1201 (.I0(\data_in_frame[17] [4]), .I1(n30090), 
            .I2(n29959), .I3(n29604), .O(n27683));
    defparam i3_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30070));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_in_frame[7] [7]), .I1(n27986), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3822));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i16_4_lut_adj_1204 (.I0(\data_out_frame[17] [0]), .I1(n28046), 
            .I2(n28040), .I3(n22_adj_3823), .O(n37));
    defparam i16_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1205 (.I0(\data_in_frame[10]_c [2]), .I1(n5_adj_3822), 
            .I2(n15914), .I3(n27996), .O(n29736));
    defparam i1_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1206 (.I0(\data_in_frame[15] [1]), .I1(n16267), 
            .I2(n14048), .I3(n16192), .O(n20_adj_3824));
    defparam i8_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i6_2_lut (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3825));
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1207 (.I0(\data_in_frame[15] [2]), .I1(n20_adj_3824), 
            .I2(n14_adj_3821), .I3(n15768), .O(n22_adj_3826));
    defparam i10_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1208 (.I0(\data_in_frame[17] [3]), .I1(n22_adj_3826), 
            .I2(n18_adj_3825), .I3(\data_in_frame[10] [3]), .O(n29875));
    defparam i11_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1209 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[13] [6]), 
            .I2(n10_adj_3827), .I3(n26977), .O(n30210));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1210 (.I0(n30192), .I1(n15768), .I2(n29736), 
            .I3(\data_in_frame[10] [6]), .O(n14_adj_3828));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1211 (.I0(\data_in_frame[17] [2]), .I1(n14_adj_3828), 
            .I2(n10_adj_3829), .I3(n29663), .O(n27633));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(n27633), .I1(n29875), .I2(GND_net), 
            .I3(GND_net), .O(n28001));
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(n27683), .I1(n29875), .I2(GND_net), 
            .I3(GND_net), .O(n27959));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1214 (.I0(n15918), .I1(n29848), .I2(n29813), 
            .I3(n8_adj_3830), .O(n31862));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1215 (.I0(n29714), .I1(n15768), .I2(n31862), 
            .I3(n30039), .O(n10_adj_3831));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_adj_1216 (.I0(\data_in_frame[12] [7]), .I1(n15905), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3832));   // verilog/coms.v(75[16:43])
    defparam i3_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1217 (.I0(\data_in_frame[17] [5]), .I1(n9_adj_3832), 
            .I2(\data_in_frame[15] [3]), .I3(n10_adj_3831), .O(n29927));
    defparam i2_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1218 (.I0(n30111), .I1(n16192), .I2(n15918), 
            .I3(n30179), .O(n20_adj_3833));
    defparam i8_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1219 (.I0(\data_in_frame[15] [4]), .I1(n30201), 
            .I2(n29714), .I3(n16336), .O(n19_adj_3834));
    defparam i7_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1220 (.I0(n7_adj_3802), .I1(\data_in_frame[9][1] ), 
            .I2(\data_in_frame[9][5] ), .I3(\data_in_frame[13] [3]), .O(n21_adj_3835));
    defparam i9_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1221 (.I0(n30210), .I1(Kp_23__N_1261), .I2(n30807), 
            .I3(n29984), .O(n29902));
    defparam i3_4_lut_adj_1221.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut_adj_1222 (.I0(n31916), .I1(n30142), .I2(n30207), 
            .I3(n30005), .O(n35));
    defparam i14_4_lut_adj_1222.LUT_INIT = 16'h9669;
    SB_LUT4 i20_4_lut_adj_1223 (.I0(n35), .I1(n37), .I2(n36_adj_3815), 
            .I3(n38), .O(n30676));
    defparam i20_4_lut_adj_1223.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1224 (.I0(n29949), .I1(\data_out_frame[23] [7]), 
            .I2(n2128), .I3(n6_adj_3836), .O(n31955));
    defparam i4_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1225 (.I0(\data_in_frame[4] [2]), .I1(n29632), 
            .I2(\data_in_frame[8] [4]), .I3(\data_in_frame[1] [4]), .O(n12_adj_3837));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1226 (.I0(n29928), .I1(n29902), .I2(GND_net), 
            .I3(GND_net), .O(n29881));
    defparam i1_2_lut_adj_1226.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1227 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[10] [3]), 
            .I2(n14048), .I3(\data_in_frame[14] [5]), .O(n4_adj_3810));
    defparam i1_2_lut_3_lut_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30114));
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1229 (.I0(n27940), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[19] [0]), .I3(n29902), .O(n10_adj_3838));
    defparam i4_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1230 (.I0(\data_in_frame[21] [5]), .I1(n29918), 
            .I2(\data_in_frame[19] [4]), .I3(\data_in_frame[19] [3]), .O(n31198));
    defparam i3_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1231 (.I0(\data_in_frame[18] [1]), .I1(n30114), 
            .I2(n29861), .I3(n6_adj_3839), .O(n31486));
    defparam i4_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1232 (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3840));   // verilog/coms.v(268[9:85])
    defparam i2_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1233 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[20] [6]), 
            .I2(\data_in_frame[18] [4]), .I3(GND_net), .O(n6_adj_3841));
    defparam i2_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1234 (.I0(n7_adj_3840), .I1(n27959), .I2(\data_in_frame[21] [6]), 
            .I3(n28001), .O(n31772));   // verilog/coms.v(268[9:85])
    defparam i4_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1235 (.I0(\data_in_frame[18] [5]), .I1(n10_adj_3838), 
            .I2(Kp_23__N_605), .I3(GND_net), .O(n31071));
    defparam i5_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1236 (.I0(\data_in_frame[19] [2]), .I1(n29924), 
            .I2(\data_in_frame[21] [3]), .I3(n27961), .O(n31237));
    defparam i3_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1237 (.I0(\data_in_frame[21] [1]), .I1(n29918), 
            .I2(n29878), .I3(n28034), .O(n31201));
    defparam i3_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1238 (.I0(\data_in_frame[18] [1]), .I1(n30213), 
            .I2(\data_in_frame[18] [2]), .I3(\data_in_frame[20] [3]), .O(n30612));
    defparam i3_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1239 (.I0(\data_in_frame[19] [6]), .I1(n29861), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3842));
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1240 (.I0(\data_in_frame[19] [2]), .I1(n27961), 
            .I2(\data_in_frame[19] [3]), .I3(GND_net), .O(n6_adj_3843));   // verilog/coms.v(268[9:85])
    defparam i2_3_lut_adj_1240.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1241 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[20] [0]), 
            .I2(n27683), .I3(n6_adj_3842), .O(n30590));
    defparam i4_4_lut_adj_1241.LUT_INIT = 16'h9669;
    SB_CARRY add_43_14 (.CI(n24875), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n24876));
    SB_LUT4 i6_4_lut_adj_1242 (.I0(n15856), .I1(n12_adj_3837), .I2(n29635), 
            .I3(\data_in_frame[0] [0]), .O(n16336));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1243 (.I0(n29733), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[7] [0]), .I3(n30048), .O(n10_adj_3844));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1244 (.I0(n29723), .I1(\data_out_frame[24] [2]), 
            .I2(n27992), .I3(GND_net), .O(n27093));
    defparam i2_3_lut_adj_1244.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[5] [1]), .I3(n15811), .O(n29905));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1245 (.I0(n27093), .I1(n4_adj_3845), .I2(n28040), 
            .I3(\data_out_frame[24] [3]), .O(n31099));
    defparam i3_4_lut_adj_1245.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1246 (.I0(n15914), .I1(n15918), .I2(\data_in_frame[9] [7]), 
            .I3(\data_in_frame[9]_c [6]), .O(n16353));
    defparam i1_2_lut_3_lut_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_LUT4 i14379_3_lut_4_lut_4_lut (.I0(n13173), .I1(n30_adj_3846), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n1), .O(n18487));   // verilog/coms.v(238[12:32])
    defparam i14379_3_lut_4_lut_4_lut.LUT_INIT = 16'h0454;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1247 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[5] [2]), .I3(\data_in_frame[2] [6]), .O(n30127));
    defparam i1_2_lut_3_lut_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1248 (.I0(n28034), .I1(n28003), .I2(\data_in_frame[21] [0]), 
            .I3(n29878), .O(n10_adj_3847));
    defparam i4_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i26551_4_lut (.I0(\data_in_frame[21] [7]), .I1(n31198), .I2(n6_adj_3848), 
            .I3(n27944), .O(n32224));
    defparam i26551_4_lut.LUT_INIT = 16'hdeed;
    SB_LUT4 i6_4_lut_adj_1249 (.I0(n30213), .I1(n31486), .I2(n8_adj_3849), 
            .I3(n30807), .O(n22_adj_3850));
    defparam i6_4_lut_adj_1249.LUT_INIT = 16'h1221;
    SB_LUT4 i26553_4_lut (.I0(\data_in_frame[21] [4]), .I1(n30590), .I2(n6_adj_3843), 
            .I3(n28003), .O(n32226));
    defparam i26553_4_lut.LUT_INIT = 16'hdeed;
    SB_LUT4 i5_4_lut_adj_1250 (.I0(n31240), .I1(n28001), .I2(n10_adj_3847), 
            .I3(n27550), .O(n21_adj_3851));
    defparam i5_4_lut_adj_1250.LUT_INIT = 16'h1441;
    SB_LUT4 i2_2_lut_adj_1251 (.I0(n29930), .I1(n27940), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3852));
    defparam i2_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1252 (.I0(n29984), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[20] [4]), .I3(n29930), .O(n31935));   // verilog/coms.v(85[17:63])
    defparam i2_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i26557_4_lut (.I0(n27402), .I1(n31772), .I2(n6_adj_3841), 
            .I3(n27940), .O(n32230));
    defparam i26557_4_lut.LUT_INIT = 16'hdeed;
    SB_LUT4 i10_4_lut_adj_1253 (.I0(n30612), .I1(n31201), .I2(n31237), 
            .I3(n31071), .O(n26));
    defparam i10_4_lut_adj_1253.LUT_INIT = 16'h0400;
    SB_LUT4 i14_4_lut_adj_1254 (.I0(n21_adj_3851), .I1(n32226), .I2(n22_adj_3850), 
            .I3(n32224), .O(n30_adj_3853));
    defparam i14_4_lut_adj_1254.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_1255 (.I0(\data_in_frame[18] [4]), .I1(n31935), 
            .I2(n6_adj_3852), .I3(\data_in_frame[20] [5]), .O(n17_adj_3854));
    defparam i1_4_lut_adj_1255.LUT_INIT = 16'h8448;
    SB_LUT4 i15_4_lut_adj_1256 (.I0(n17_adj_3854), .I1(n30_adj_3853), .I2(n26), 
            .I3(n32230), .O(n30_adj_3846));
    defparam i15_4_lut_adj_1256.LUT_INIT = 16'h0080;
    SB_LUT4 i12888_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[2]), 
            .I3(\data_in_frame[10]_c [2]), .O(n16997));
    defparam i12888_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12835_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n16944));
    defparam i12835_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12836_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n16945));
    defparam i12836_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12837_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n16946));
    defparam i12837_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1257 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[5] [6]), .O(n29700));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_13_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n24874), .O(n2_adj_3755)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_13 (.CI(n24874), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n24875));
    SB_LUT4 i1_2_lut_adj_1258 (.I0(n27977), .I1(n30099), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3855));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1259 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n29816), .I3(n6_adj_3855), .O(n27992));
    defparam i4_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i12889_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[1]), 
            .I3(\data_in_frame[10][1] ), .O(n16998));
    defparam i12889_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12838_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n16947));
    defparam i12838_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12890_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29552), .I2(rx_data[0]), 
            .I3(\data_in_frame[10]_c [0]), .O(n16999));
    defparam i12890_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1260 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[5] [0]), .O(n16107));
    defparam i1_2_lut_3_lut_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1261 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[6] [1]), 
            .I2(n30093), .I3(\data_in_frame[6] [7]), .O(Kp_23__N_912));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1262 (.I0(n15823), .I1(n16245), .I2(\data_in_frame[4] [5]), 
            .I3(n27008), .O(n30029));
    defparam i1_2_lut_4_lut_adj_1262.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1263 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[6] [7]), 
            .I2(n16107), .I3(\data_in_frame[7] [1]), .O(n29726));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29744));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n34801));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n34801_bdd_4_lut (.I0(n34801), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n34804));
    defparam n34801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1265 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[4] [6]), .O(n30048));
    defparam i1_2_lut_3_lut_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n34534), .I2(n33151), .I3(byte_transmit_counter[4]), .O(n34795));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n34795_bdd_4_lut (.I0(n34795), .I1(n14_adj_3643), .I2(n7_adj_3642), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n34795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[20] [0]), .I1(n27992), 
            .I2(GND_net), .I3(GND_net), .O(n28040));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1267 (.I0(n28013), .I1(n29939), .I2(n28040), 
            .I3(\data_out_frame[24] [4]), .O(n31372));
    defparam i3_4_lut_adj_1267.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1268 (.I0(n31856), .I1(\data_out_frame[24] [5]), 
            .I2(n28013), .I3(\data_out_frame[25] [0]), .O(n31011));
    defparam i3_4_lut_adj_1268.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1269 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n15823));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1269.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1270 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n29632));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1270.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1271 (.I0(n16070), .I1(n15853), .I2(n29892), 
            .I3(n6_adj_3856), .O(n31856));
    defparam i4_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i12839_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n16948));
    defparam i12839_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1272 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n15866));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1272.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(\data_in_frame[7] [4]), .I1(n29898), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n30219));
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1274 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n29787));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1274.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1275 (.I0(n27239), .I1(n29851), .I2(n31856), 
            .I3(GND_net), .O(n30501));
    defparam i2_3_lut_adj_1275.LUT_INIT = 16'h6969;
    SB_LUT4 i12840_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n16949));
    defparam i12840_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12841_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n16950));
    defparam i12841_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(n30017), .I1(n27977), .I2(\data_out_frame[19] [5]), 
            .I3(n30176), .O(n10_adj_3857));
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1277 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(n29621), .I3(\data_in_frame[4] [6]), .O(n19_adj_3858));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n15890));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29071 (.I0(byte_transmit_counter[3]), 
            .I1(n34540), .I2(n33148), .I3(byte_transmit_counter[4]), .O(n34789));
    defparam byte_transmit_counter_3__bdd_4_lut_29071.LUT_INIT = 16'he4aa;
    SB_LUT4 n34789_bdd_4_lut (.I0(n34789), .I1(n14_adj_3635), .I2(n7_adj_3634), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n34789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1279 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [5]), 
            .I2(n15890), .I3(n29787), .O(n10_adj_3859));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29076 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n34783));
    defparam byte_transmit_counter_0__bdd_4_lut_29076.LUT_INIT = 16'he4aa;
    SB_LUT4 n34783_bdd_4_lut (.I0(n34783), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n34786));
    defparam n34783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29061 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n34777));
    defparam byte_transmit_counter_0__bdd_4_lut_29061.LUT_INIT = 16'he4aa;
    SB_LUT4 n34777_bdd_4_lut (.I0(n34777), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n34780));
    defparam n34777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 equal_1123_i8_2_lut (.I0(Kp_23__N_958), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3830));   // verilog/coms.v(236[9:81])
    defparam equal_1123_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(n16034), .I1(n30057), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3860));
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29056 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n34771));
    defparam byte_transmit_counter_0__bdd_4_lut_29056.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1281 (.I0(n27067), .I1(\data_out_frame[19] [7]), 
            .I2(n29751), .I3(n6_adj_3860), .O(n2143));
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 n34771_bdd_4_lut (.I0(n34771), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n34774));
    defparam n34771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1282 (.I0(n29595), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[6] [5]), .O(n14_adj_3861));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29051 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n34765));
    defparam byte_transmit_counter_0__bdd_4_lut_29051.LUT_INIT = 16'he4aa;
    SB_LUT4 n34765_bdd_4_lut (.I0(n34765), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n34768));
    defparam n34765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1283 (.I0(\data_out_frame[20] [1]), .I1(n2143), 
            .I2(n28046), .I3(GND_net), .O(n28013));
    defparam i2_3_lut_adj_1283.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1284 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[2] [3]), .O(n13_adj_3862));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i12842_3_lut_4_lut (.I0(n8_adj_3669), .I1(n29530), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n16951));
    defparam i12842_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29046 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n34759));
    defparam byte_transmit_counter_0__bdd_4_lut_29046.LUT_INIT = 16'he4aa;
    SB_LUT4 i12827_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n16936));
    defparam i12827_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1285 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(GND_net), .O(n30096));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1285.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1286 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n30176));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i12828_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n16937));
    defparam i12828_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12861_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n16970));
    defparam i12861_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(n1516), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30108));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1288 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[17] [3]), 
            .I2(n27479), .I3(\data_out_frame[15] [1]), .O(n29660));
    defparam i2_4_lut_adj_1288.LUT_INIT = 16'h9669;
    SB_LUT4 i12829_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n16938));
    defparam i12829_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12830_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n16939));
    defparam i12830_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1289 (.I0(n30017), .I1(\data_out_frame[17] [6]), 
            .I2(n16479), .I3(n27067), .O(n14_adj_3863));
    defparam i6_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1290 (.I0(n27977), .I1(n14_adj_3863), .I2(n10_adj_3864), 
            .I3(\data_out_frame[20] [0]), .O(n29800));
    defparam i7_4_lut_adj_1290.LUT_INIT = 16'h9669;
    SB_LUT4 n34759_bdd_4_lut (.I0(n34759), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n34762));
    defparam n34759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 equal_1123_i7_3_lut (.I0(n13_adj_3862), .I1(\data_in_frame[8] [6]), 
            .I2(n14_adj_3861), .I3(GND_net), .O(n7_adj_3802));   // verilog/coms.v(236[9:81])
    defparam equal_1123_i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29041 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n34753));
    defparam byte_transmit_counter_0__bdd_4_lut_29041.LUT_INIT = 16'he4aa;
    SB_LUT4 n34753_bdd_4_lut (.I0(n34753), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n34756));
    defparam n34753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1291 (.I0(n30108), .I1(n29660), .I2(n29642), 
            .I3(n30176), .O(n10_adj_3719));
    defparam i4_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1292 (.I0(n30127), .I1(n30219), .I2(\data_in_frame[0] [4]), 
            .I3(GND_net), .O(n15918));
    defparam i2_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29036 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n34747));
    defparam byte_transmit_counter_0__bdd_4_lut_29036.LUT_INIT = 16'he4aa;
    SB_LUT4 n34747_bdd_4_lut (.I0(n34747), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n34750));
    defparam n34747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1293 (.I0(n15866), .I1(n29632), .I2(\data_in_frame[6] [4]), 
            .I3(\data_in_frame[4] [3]), .O(n12_adj_3865));   // verilog/coms.v(166[9:87])
    defparam i5_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29031 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n34741));
    defparam byte_transmit_counter_0__bdd_4_lut_29031.LUT_INIT = 16'he4aa;
    SB_LUT4 n34741_bdd_4_lut (.I0(n34741), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n34744));
    defparam n34741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1294 (.I0(\data_in_frame[8] [5]), .I1(n12_adj_3865), 
            .I2(n29647), .I3(\data_in_frame[6] [3]), .O(n15768));   // verilog/coms.v(166[9:87])
    defparam i6_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29026 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n34735));
    defparam byte_transmit_counter_0__bdd_4_lut_29026.LUT_INIT = 16'he4aa;
    SB_LUT4 n34735_bdd_4_lut (.I0(n34735), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n34738));
    defparam n34735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1295 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n3_adj_3866));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29021 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n34729));
    defparam byte_transmit_counter_0__bdd_4_lut_29021.LUT_INIT = 16'he4aa;
    SB_LUT4 n34729_bdd_4_lut (.I0(n34729), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n34732));
    defparam n34729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1296 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(\data_in_frame[0] [2]), .O(n29733));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i12831_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n16940));
    defparam i12831_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12832_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n16941));
    defparam i12832_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_in_frame[1] [5]), .I1(n30011), 
            .I2(GND_net), .I3(GND_net), .O(n29598));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i12833_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n16942));
    defparam i12833_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12834_3_lut_4_lut (.I0(n8_adj_3820), .I1(n29530), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n16943));
    defparam i12834_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1298 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[15] [0]), 
            .I2(n15905), .I3(n16336), .O(n30067));
    defparam i2_3_lut_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n29689));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_adj_1300 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [5]), 
            .I2(n29660), .I3(GND_net), .O(n10_adj_3864));
    defparam i2_2_lut_3_lut_adj_1300.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29016 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n34723));
    defparam byte_transmit_counter_0__bdd_4_lut_29016.LUT_INIT = 16'he4aa;
    SB_LUT4 n34723_bdd_4_lut (.I0(n34723), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n34726));
    defparam n34723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1301 (.I0(\data_out_frame[12] [5]), .I1(n1519), 
            .I2(\data_out_frame[17] [4]), .I3(GND_net), .O(n30017));
    defparam i1_2_lut_3_lut_adj_1301.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n29692));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1303 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n29647));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1303.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29011 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n34705));
    defparam byte_transmit_counter_0__bdd_4_lut_29011.LUT_INIT = 16'he4aa;
    SB_LUT4 n34705_bdd_4_lut (.I0(n34705), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n34708));
    defparam n34705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1304 (.I0(\data_out_frame[15] [1]), .I1(n1516), 
            .I2(\data_out_frame[19] [4]), .I3(GND_net), .O(n29910));
    defparam i1_2_lut_3_lut_adj_1304.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28996 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n34699));
    defparam byte_transmit_counter_0__bdd_4_lut_28996.LUT_INIT = 16'he4aa;
    SB_LUT4 n34699_bdd_4_lut (.I0(n34699), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n34702));
    defparam n34699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1305 (.I0(\data_in_frame[0] [6]), .I1(n15811), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n16604));
    defparam i2_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1306 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[15] [0]), 
            .I2(n16336), .I3(GND_net), .O(n10_adj_3829));
    defparam i2_2_lut_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1307 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n29595));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1307.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1308 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n29898));
    defparam i2_3_lut_adj_1308.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1309 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[5] [1]), 
            .I2(n15811), .I3(GND_net), .O(n30243));
    defparam i2_3_lut_adj_1309.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30173));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1311 (.I0(\data_in_frame[5] [5]), .I1(n29898), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[5] [4]), .O(n15720));
    defparam i3_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28991 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n34693));
    defparam byte_transmit_counter_0__bdd_4_lut_28991.LUT_INIT = 16'he4aa;
    SB_LUT4 n34693_bdd_4_lut (.I0(n34693), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n34696));
    defparam n34693_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12963_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n17072));
    defparam i12963_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1312 (.I0(n2128), .I1(n2125), .I2(\data_out_frame[23] [5]), 
            .I3(n30124), .O(n6_adj_3856));
    defparam i1_2_lut_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28986 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n34687));
    defparam byte_transmit_counter_0__bdd_4_lut_28986.LUT_INIT = 16'he4aa;
    SB_LUT4 n34687_bdd_4_lut (.I0(n34687), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n34690));
    defparam n34687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1313 (.I0(\data_in_frame[4] [5]), .I1(n27008), 
            .I2(n30081), .I3(Kp_23__N_764), .O(n27996));
    defparam i2_3_lut_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28981 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n34681));
    defparam byte_transmit_counter_0__bdd_4_lut_28981.LUT_INIT = 16'he4aa;
    SB_LUT4 i12964_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n17073));
    defparam i12964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n34681_bdd_4_lut (.I0(n34681), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n34684));
    defparam n34681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1314 (.I0(\data_in_frame[2] [1]), .I1(n29692), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [7]), .O(n10_adj_3868));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1315 (.I0(n30183), .I1(n29621), .I2(n10_adj_3868), 
            .I3(\data_in_frame[0] [5]), .O(n20_adj_3869));   // verilog/coms.v(78[16:27])
    defparam i2_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28976 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n34669));
    defparam byte_transmit_counter_0__bdd_4_lut_28976.LUT_INIT = 16'he4aa;
    SB_LUT4 n34669_bdd_4_lut (.I0(n34669), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n34672));
    defparam n34669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12965_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n17074));
    defparam i12965_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12966_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n17075));
    defparam i12966_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1316 (.I0(Kp_23__N_737), .I1(n19_adj_3858), .I2(\data_in_frame[4] [7]), 
            .I3(n20_adj_3869), .O(n32));   // verilog/coms.v(78[16:27])
    defparam i14_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i12967_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n17076));
    defparam i12967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1317 (.I0(n15720), .I1(n30173), .I2(n30243), 
            .I3(n30096), .O(n30_adj_3870));   // verilog/coms.v(78[16:27])
    defparam i12_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i12968_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n17077));
    defparam i12968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12969_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n17078));
    defparam i12969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12757_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29558), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n16866));
    defparam i12757_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_76_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_3699));   // verilog/coms.v(154[7:23])
    defparam equal_76_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_84_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_3867));   // verilog/coms.v(154[7:23])
    defparam equal_84_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13_4_lut_adj_1318 (.I0(n29595), .I1(\data_in_frame[3] [1]), 
            .I2(n3_adj_3866), .I3(n16604), .O(n31));   // verilog/coms.v(78[16:27])
    defparam i13_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1319 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[3] [3]), 
            .I2(n30127), .I3(\data_in_frame[5] [7]), .O(n29_adj_3871));   // verilog/coms.v(78[16:27])
    defparam i11_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i19794_3_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n92), 
            .I2(DE_c), .I3(\FRAME_MATCHER.state[0] ), .O(n17388));   // verilog/coms.v(112[11:16])
    defparam i19794_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i17_4_lut_adj_1320 (.I0(n29_adj_3871), .I1(n31), .I2(n30_adj_3870), 
            .I3(n32), .O(n27008));   // verilog/coms.v(78[16:27])
    defparam i17_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1321 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(n29700), .I3(GND_net), .O(n30183));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1321.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(\data_in_frame[4] [5]), .I1(n27008), 
            .I2(GND_net), .I3(GND_net), .O(n29934));
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28966 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n34657));
    defparam byte_transmit_counter_0__bdd_4_lut_28966.LUT_INIT = 16'he4aa;
    SB_LUT4 n34657_bdd_4_lut (.I0(n34657), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n34660));
    defparam n34657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(n15823), .I1(n16245), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_764));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29066 (.I0(byte_transmit_counter[3]), 
            .I1(n34546), .I2(n33195), .I3(byte_transmit_counter[4]), .O(n34651));
    defparam byte_transmit_counter_3__bdd_4_lut_29066.LUT_INIT = 16'he4aa;
    SB_LUT4 n34651_bdd_4_lut (.I0(n34651), .I1(n14_adj_3624), .I2(n7_adj_3620), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n34651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n29810));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_28951 (.I0(byte_transmit_counter[3]), 
            .I1(n34552), .I2(n33188), .I3(byte_transmit_counter[4]), .O(n34645));
    defparam byte_transmit_counter_3__bdd_4_lut_28951.LUT_INIT = 16'he4aa;
    SB_LUT4 n34645_bdd_4_lut (.I0(n34645), .I1(n14_adj_3615), .I2(n7), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n34645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1325 (.I0(n29810), .I1(n30093), .I2(\data_in_frame[6] [7]), 
            .I3(n16280), .O(n30081));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1326 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(Kp_23__N_737), .O(n29968));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1327 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n29831));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1327.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1328 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(n29968), .O(n15811));   // verilog/coms.v(73[16:34])
    defparam i2_3_lut_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_28946 (.I0(byte_transmit_counter[3]), 
            .I1(n34558), .I2(n33171), .I3(byte_transmit_counter[4]), .O(n34639));
    defparam byte_transmit_counter_3__bdd_4_lut_28946.LUT_INIT = 16'he4aa;
    SB_LUT4 n34639_bdd_4_lut (.I0(n34639), .I1(n14_adj_3872), .I2(n7_adj_3873), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n34639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_28941 (.I0(byte_transmit_counter[3]), 
            .I1(n34564), .I2(n33168), .I3(byte_transmit_counter[4]), .O(n34633));
    defparam byte_transmit_counter_3__bdd_4_lut_28941.LUT_INIT = 16'he4aa;
    SB_LUT4 n34633_bdd_4_lut (.I0(n34633), .I1(n14_adj_3874), .I2(n7_adj_3875), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n34633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_28936 (.I0(byte_transmit_counter[3]), 
            .I1(n34570), .I2(n33165), .I3(byte_transmit_counter[4]), .O(n34627));
    defparam byte_transmit_counter_3__bdd_4_lut_28936.LUT_INIT = 16'he4aa;
    SB_LUT4 n34627_bdd_4_lut (.I0(n34627), .I1(n14_adj_3876), .I2(n7_adj_3877), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n34627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1329 (.I0(n15666), .I1(\data_out_frame[24] [3]), 
            .I2(\data_out_frame[24] [4]), .I3(n4_adj_3845), .O(n29835));
    defparam i1_2_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_28931 (.I0(byte_transmit_counter[3]), 
            .I1(n34576), .I2(n33159), .I3(byte_transmit_counter[4]), .O(n34621));
    defparam byte_transmit_counter_3__bdd_4_lut_28931.LUT_INIT = 16'he4aa;
    SB_LUT4 n34621_bdd_4_lut (.I0(n34621), .I1(n14_adj_3878), .I2(n7_adj_3879), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n34621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1330 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29621));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1330.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_12_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n24873), .O(n2_adj_3757)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28956 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n34615));
    defparam byte_transmit_counter_0__bdd_4_lut_28956.LUT_INIT = 16'he4aa;
    SB_LUT4 n34615_bdd_4_lut (.I0(n34615), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n34618));
    defparam n34615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [4]), 
            .I2(n4_adj_3845), .I3(GND_net), .O(n29834));
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29740));
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1333 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[19] [1]), 
            .I2(n28034), .I3(n27550), .O(n31240));
    defparam i2_3_lut_4_lut_adj_1333.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1334 (.I0(\data_in_frame[2] [5]), .I1(n29621), 
            .I2(n10_adj_3880), .I3(n29740), .O(n16011));
    defparam i5_3_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_CARRY add_43_12 (.CI(n24873), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n24874));
    SB_LUT4 i2_3_lut_4_lut_adj_1335 (.I0(\data_in_frame[1] [3]), .I1(n29689), 
            .I2(\data_in_frame[7] [6]), .I3(n15720), .O(n15914));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_11_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n24872), .O(n2_adj_3759)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_11 (.CI(n24872), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n24873));
    SB_LUT4 i3_3_lut_4_lut (.I0(n29928), .I1(n29902), .I2(\data_in_frame[20] [1]), 
            .I3(\data_in_frame[19] [7]), .O(n8_adj_3849));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28922 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n34591));
    defparam byte_transmit_counter_0__bdd_4_lut_28922.LUT_INIT = 16'he4aa;
    SB_LUT4 n34591_bdd_4_lut (.I0(n34591), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n34594));
    defparam n34591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_737));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28903 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n34585));
    defparam byte_transmit_counter_0__bdd_4_lut_28903.LUT_INIT = 16'he4aa;
    SB_LUT4 n34585_bdd_4_lut (.I0(n34585), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n34588));
    defparam n34585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1336 (.I0(\data_in_frame[20] [2]), .I1(n30084), 
            .I2(n10_adj_3827), .I3(n26977), .O(n6_adj_3839));
    defparam i1_2_lut_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28898 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n34579));
    defparam byte_transmit_counter_0__bdd_4_lut_28898.LUT_INIT = 16'he4aa;
    SB_LUT4 n34579_bdd_4_lut (.I0(n34579), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n34582));
    defparam n34579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1337 (.I0(\data_in_frame[1] [3]), .I1(n29689), 
            .I2(\data_in_frame[5] [5]), .I3(n16220), .O(n16280));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_10_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n24871), .O(n2_adj_3761)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n24871), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n24872));
    SB_LUT4 add_43_9_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n24870), .O(n2_adj_3763)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n29971));
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1339 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(n10_adj_3881), .I3(\data_in_frame[1] [4]), .O(n29837));   // verilog/coms.v(78[16:27])
    defparam i5_3_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_CARRY add_43_9 (.CI(n24870), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n24871));
    SB_LUT4 add_43_8_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n24869), .O(n2_adj_3765)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n24901), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3882));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1340 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[3] [6]), .O(n30011));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_CARRY add_43_8 (.CI(n24869), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n24870));
    SB_LUT4 add_43_7_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n24868), .O(n2_adj_3767)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n24900), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_8 (.CI(n24900), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n24901));
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n24899), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_7 (.CI(n24868), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n24869));
    SB_LUT4 i5_3_lut_4_lut_adj_1341 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[5] [7]), 
            .I2(n10_adj_3812), .I3(\data_in_frame[6] [0]), .O(n30036));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3883));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_6_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n24867), .O(n2_adj_3769)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3971_7 (.CI(n24899), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n24900));
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n24898), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1342 (.I0(\data_in_frame[19] [6]), .I1(n27683), 
            .I2(n29875), .I3(\data_in_frame[19] [5]), .O(n6_adj_3848));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1342.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[14] [6]), .I3(GND_net), .O(n30192));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_CARRY add_3971_6 (.CI(n24898), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n24899));
    SB_CARRY add_43_6 (.CI(n24867), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n24868));
    SB_LUT4 add_43_5_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n24866), .O(n2_adj_3771)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n24897), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_5 (.CI(n24866), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n24867));
    SB_CARRY add_3971_5 (.CI(n24897), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n24898));
    SB_LUT4 i1_2_lut_4_lut_adj_1344 (.I0(n29910), .I1(n10_adj_3857), .I2(n27938), 
            .I3(\data_out_frame[23] [6]), .O(n29949));
    defparam i1_2_lut_4_lut_adj_1344.LUT_INIT = 16'h9669;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n24896), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1345 (.I0(n29910), .I1(n10_adj_3857), .I2(n27938), 
            .I3(\data_out_frame[20] [0]), .O(n29723));
    defparam i1_2_lut_4_lut_adj_1345.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_4_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n24865), .O(n2_adj_3773)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_3_lut_4_lut_adj_1346 (.I0(n3_adj_3866), .I1(n16245), .I2(n10_adj_3844), 
            .I3(\data_in_frame[4] [4]), .O(n16333));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1347 (.I0(n3_adj_3866), .I1(n16245), .I2(n10_adj_3859), 
            .I3(n15823), .O(Kp_23__N_958));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i12862_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n16971));
    defparam i12862_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1348 (.I0(n13173), .I1(n30_adj_3846), 
            .I2(n18751), .I3(\FRAME_MATCHER.state[2] ), .O(n8868));   // verilog/coms.v(238[12:32])
    defparam i1_2_lut_3_lut_4_lut_adj_1348.LUT_INIT = 16'h0400;
    SB_LUT4 i2_4_lut_4_lut (.I0(n29800), .I1(\data_out_frame[20] [1]), .I2(n2143), 
            .I3(n27980), .O(n4_adj_3845));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1349 (.I0(n29864), .I1(\data_out_frame[24] [1]), 
            .I2(n28040), .I3(\data_out_frame[24] [0]), .O(n6_adj_3836));
    defparam i1_2_lut_4_lut_adj_1349.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1350 (.I0(n29864), .I1(\data_out_frame[24] [1]), 
            .I2(n28040), .I3(n27093), .O(n16060));
    defparam i1_2_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_4 (.CI(n24896), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n24897));
    SB_CARRY add_43_4 (.CI(n24865), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n24866));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n24895), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1351 (.I0(n21_adj_3835), .I1(n19_adj_3834), 
            .I2(n20_adj_3833), .I3(n29927), .O(n29928));
    defparam i1_2_lut_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n16652), .D(n8825[0]), .R(n16773));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1352 (.I0(n21_adj_3835), .I1(n19_adj_3834), 
            .I2(n20_adj_3833), .I3(n30231), .O(n29861));
    defparam i1_2_lut_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_3 (.CI(n24895), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n24896));
    SB_LUT4 add_43_3_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n24864), .O(n2_adj_3775)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1353 (.I0(\data_in_frame[12] [6]), .I1(n10_adj_3818), 
            .I2(\data_in_frame[10] [5]), .I3(n27633), .O(n28003));
    defparam i1_2_lut_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1354 (.I0(\data_in_frame[12] [6]), .I1(n10_adj_3818), 
            .I2(\data_in_frame[10] [5]), .I3(n29875), .O(n29918));
    defparam i1_2_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1355 (.I0(\data_in_frame[12] [6]), .I1(n10_adj_3818), 
            .I2(\data_in_frame[10] [5]), .I3(n30216), .O(n27961));
    defparam i1_2_lut_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3257), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_3 (.CI(n24864), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n24865));
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3257), 
            .CO(n24895));
    SB_LUT4 add_43_33_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n24894), .O(n2_adj_3722)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_2_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_c)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n24864));
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(\data_in_frame[8] [1]), .I1(n14041), 
            .I2(n29837), .I3(GND_net), .O(n27986));
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(\data_in_frame[8] [1]), .I1(n14041), 
            .I2(n15951), .I3(GND_net), .O(n14048));
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_32_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n24893), .O(n2_adj_3725)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n24893), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n24894));
    SB_LUT4 i2_3_lut_adj_1358 (.I0(n29831), .I1(n29968), .I2(\data_in_frame[3] [1]), 
            .I3(GND_net), .O(n16493));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1358.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_31_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n24892), .O(n2_adj_3727)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(n15914), .I1(n15918), .I2(n16336), 
            .I3(GND_net), .O(n30023));
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_CARRY add_43_31 (.CI(n24892), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n24893));
    SB_LUT4 i2_3_lut_4_lut_adj_1360 (.I0(\data_in_frame[16] [4]), .I1(n29915), 
            .I2(\data_in_frame[18] [6]), .I3(n29698), .O(n30249));
    defparam i2_3_lut_4_lut_adj_1360.LUT_INIT = 16'h9669;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n16898));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1361 (.I0(\data_in_frame[16] [4]), .I1(n29915), 
            .I2(n26998), .I3(\data_in_frame[16] [3]), .O(n27402));
    defparam i2_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(n16011), .I1(n16329), .I2(\data_in_frame[14] [1]), 
            .I3(GND_net), .O(n6_adj_3806));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n33160), .I2(n33161), .I3(byte_transmit_counter[2]), .O(n34573));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1363 (.I0(n16011), .I1(n16329), .I2(n16333), 
            .I3(n10_adj_3704), .O(n30179));
    defparam i1_2_lut_3_lut_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(n16011), .I1(n16329), .I2(\data_in_frame[9][4] ), 
            .I3(GND_net), .O(n29767));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_30_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n24891), .O(n2_adj_3729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(n10_adj_3704), .I1(n16333), .I2(n29767), 
            .I3(GND_net), .O(n26977));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1366 (.I0(n15905), .I1(n15951), .I2(Kp_23__N_1054), 
            .I3(\data_in_frame[9][0] ), .O(n29959));
    defparam i2_3_lut_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_CARRY add_43_30 (.CI(n24891), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n24892));
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(n10_adj_3704), .I1(n16333), .I2(\data_in_frame[13] [4]), 
            .I3(n29717), .O(n15947));   // verilog/coms.v(72[16:41])
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_29_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n24890), .O(n2_adj_3731)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(n10_adj_3704), .I1(n16329), .I2(\data_in_frame[9][3] ), 
            .I3(GND_net), .O(n16445));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(n10_adj_3704), .I1(n16329), .I2(n27061), 
            .I3(GND_net), .O(n30111));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1370 (.I0(\data_in_frame[9][0] ), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[10] [7]), .I3(GND_net), .O(n30201));
    defparam i1_2_lut_3_lut_adj_1370.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(\data_in_frame[9][0] ), .I1(\data_in_frame[11] [2]), 
            .I2(Kp_23__N_1054), .I3(GND_net), .O(n15777));
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1372 (.I0(n16333), .I1(Kp_23__N_958), .I2(n30246), 
            .I3(n29754), .O(n29609));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n16897));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(n16333), .I1(Kp_23__N_958), .I2(\data_in_frame[8] [1]), 
            .I3(GND_net), .O(n6_adj_3801));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(Kp_23__N_958), .I1(\data_in_frame[8] [7]), 
            .I2(n7_adj_3802), .I3(GND_net), .O(Kp_23__N_1054));
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n16896));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n16895));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n16894));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n16893));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n16892));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n16891));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n16890));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n16889));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n16888));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n16887));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n16886));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n16885));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n16884));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n16883));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n16882));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n16881));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n16880));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n16879));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n16878));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n16877));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n16876));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n16875));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n16874));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state[2] ), .C(clk32MHz), 
           .D(n35073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n28937));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n16868));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n16867));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n16866));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1375 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n29663));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1376 (.I0(\data_in_frame[10] [4]), .I1(n15905), 
            .I2(n15951), .I3(GND_net), .O(n6_adj_3816));
    defparam i1_2_lut_3_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1377 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[16] [7]), 
            .I2(n16368), .I3(GND_net), .O(n30258));
    defparam i1_2_lut_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_LUT4 select_295_Select_1_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_3776));
    defparam select_295_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_2_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_3774));
    defparam select_295_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_3_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_3772));
    defparam select_295_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_4_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_3770));
    defparam select_295_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_5_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_3768));
    defparam select_295_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_6_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_3766));
    defparam select_295_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_DFFE driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .E(VCC_net), .D(n17388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n17373));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_295_Select_7_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_3764));
    defparam select_295_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_8_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_3762));
    defparam select_295_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n17372));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n17371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n17370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n17369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n17368));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n17367));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n34573_bdd_4_lut (.I0(n34573), .I1(n17_adj_3883), .I2(n16_adj_3882), 
            .I3(byte_transmit_counter[2]), .O(n34576));
    defparam n34573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1378 (.I0(\data_in_frame[7] [3]), .I1(n29905), 
            .I2(n16493), .I3(\data_in_frame[4] [7]), .O(n10_adj_3880));
    defparam i4_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 select_295_Select_9_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_3760));
    defparam select_295_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_10_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_3758));
    defparam select_295_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_11_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_3756));
    defparam select_295_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i2_3_lut_4_lut_adj_1379 (.I0(n16094), .I1(\data_in_frame[10][1] ), 
            .I2(n30036), .I3(\data_in_frame[12] [3]), .O(n16368));
    defparam i2_3_lut_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 select_295_Select_12_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_3754));
    defparam select_295_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_3_lut_adj_1380 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[10] [3]), 
            .I2(n14048), .I3(GND_net), .O(n29784));
    defparam i1_2_lut_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n17335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n17334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n17333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n17332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n17331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n17330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n17329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n17328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n17327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n17326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n17325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n17324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n17323));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n17322));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n17321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n17320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n17314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n17313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n17312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n17311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n17310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n17309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n17308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n17307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n17306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n17305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n17304));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n17303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n17302));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n17301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n17300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n17299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n17298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n17297));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n17296));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n17295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n17294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n17293));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n17292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n17291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n17290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n17289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n17288));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n17287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n17286));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n17285));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n17284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n17283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n17282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n17281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n17280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n17279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n17278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n17277));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n17276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n17275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n17274));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n17273));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n17272));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n17271));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n17270));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n17269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n17268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n17267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n17266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n17265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n17264));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n17263));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n17262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n17261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n17260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n17259));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n17258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n17257));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n17256));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n17255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n17254));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n17253));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n17252));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n17251));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n17250));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n17249));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n17248));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n17247));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n17246));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n17245));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n17244));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n17243));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n17242));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n17241));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n17240));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n17239));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n17238));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n17237));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n17236));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n17235));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n17234));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n17233));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n17232));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_295_Select_13_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_3752));
    defparam select_295_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i4_4_lut_adj_1381 (.I0(\data_in_frame[8] [0]), .I1(n29700), 
            .I2(Kp_23__N_912), .I3(n30029), .O(n10_adj_3881));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1382 (.I0(Kp_23__N_764), .I1(n29934), .I2(n30145), 
            .I3(\data_in_frame[11] [7]), .O(n30228));
    defparam i2_3_lut_4_lut_adj_1382.LUT_INIT = 16'h9669;
    SB_LUT4 select_295_Select_14_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_3750));
    defparam select_295_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1383 (.I0(n21151), .I1(n8_adj_3669), .I2(GND_net), 
            .I3(GND_net), .O(n29558));
    defparam i1_2_lut_adj_1383.LUT_INIT = 16'hdddd;
    SB_LUT4 select_295_Select_15_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_3748));
    defparam select_295_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_4_lut_adj_1384 (.I0(\data_in_frame[9][3] ), .I1(\data_in_frame[9][2] ), 
            .I2(\data_in_frame[9][1] ), .I3(\data_in_frame[9][4] ), .O(n16204));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1385 (.I0(n27683), .I1(n29875), .I2(n27961), 
            .I3(GND_net), .O(n16098));
    defparam i1_2_lut_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 select_295_Select_16_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_3747));
    defparam select_295_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_4_lut_adj_1386 (.I0(n30029), .I1(n30145), .I2(\data_in_frame[11] [7]), 
            .I3(n16011), .O(n8_adj_3800));
    defparam i1_2_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i14583_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10]_c [0]), 
            .I2(n4216), .I3(GND_net), .O(n16868));
    defparam i14583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_in_frame[12] [1]), .I1(n16011), 
            .I2(\data_in_frame[10]_c [0]), .I3(GND_net), .O(n9_adj_3798));
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 select_295_Select_17_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_3746));
    defparam select_295_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i12863_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n16972));
    defparam i12863_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n6_adj_3794));
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'h0404;
    SB_LUT4 select_295_Select_18_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_3745));
    defparam select_295_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i17146_3_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n63_adj_3689), 
            .I2(n63_adj_3692), .I3(GND_net), .O(n122));   // verilog/coms.v(139[4] 141[7])
    defparam i17146_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_323_Select_2_i5_4_lut (.I0(n122), .I1(\FRAME_MATCHER.i_31__N_2368 ), 
            .I2(n3303), .I3(n63), .O(n5));
    defparam select_323_Select_2_i5_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i17140_rep_195_2_lut (.I0(n122), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n35368));   // verilog/coms.v(142[4] 144[7])
    defparam i17140_rep_195_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_295_Select_19_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_3744));
    defparam select_295_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n17231));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n17230));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n17229));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n17228));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n17227));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n17226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n17225));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n17224));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n17223));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n17222));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n17221));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n17220));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n17219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n17218));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n17217));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n17216));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n17215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n17214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n17213));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n17212));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n17211));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n17210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n17209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n17208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n17207));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n17206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n17205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n17204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n17203));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n17202));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n17201));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n17200));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n17199));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n17198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n17197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n17196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n17195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n17194));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n17193));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n17192));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n17191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n17190));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n17189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n17188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n17187));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n17186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n17185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n17184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n17183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n17182));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n17181));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n17180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n17179));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n17178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n17177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n17176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n17175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n17174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n17173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n17172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n17171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n17170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n17169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n17168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n17167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n17166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n17165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n17164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n17163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n17162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n17161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n17160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n17159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n17158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n17157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n17156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n17155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n17154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n17153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n17152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n17151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n17150));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n17149));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n17148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n17147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n17146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n17145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n17144));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n17143));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n17142));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n17141));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n17140));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n17139));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n17138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n17137));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n17136));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n17135));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n17134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n17133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n17132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n17131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n17130));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n17129));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n17128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n17127));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n17126));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n17125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n17124));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n17123));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n17122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n17121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n17120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n17119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n17118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n17117));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_295_Select_20_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_3743));
    defparam select_295_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i2_3_lut_4_lut_adj_1389 (.I0(n13916), .I1(n27952), .I2(n16054), 
            .I3(n15266), .O(n27076));
    defparam i2_3_lut_4_lut_adj_1389.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(n13916), .I1(n27952), .I2(\data_out_frame[23] [2]), 
            .I3(GND_net), .O(n30102));
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h6969;
    SB_LUT4 i12875_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n16984));
    defparam i12875_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12876_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n16985));
    defparam i12876_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_295_Select_21_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_3742));
    defparam select_295_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_22_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_3741));
    defparam select_295_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_23_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_3740));
    defparam select_295_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_24_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_3738));
    defparam select_295_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_25_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_3736));
    defparam select_295_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_26_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_3734));
    defparam select_295_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i12877_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n16986));
    defparam i12877_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_295_Select_27_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_3732));
    defparam select_295_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_28_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_3730));
    defparam select_295_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i5_3_lut_4_lut_adj_1391 (.I0(\data_in_frame[18] [5]), .I1(n27959), 
            .I2(n27961), .I3(\data_in_frame[18] [4]), .O(n17_adj_3787));
    defparam i5_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 select_295_Select_29_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_3728));
    defparam select_295_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_30_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_3726));
    defparam select_295_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_295_Select_31_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_3723));
    defparam select_295_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_28888 (.I0(byte_transmit_counter[1]), 
            .I1(n33166), .I2(n33167), .I3(byte_transmit_counter[2]), .O(n34567));
    defparam byte_transmit_counter_1__bdd_4_lut_28888.LUT_INIT = 16'he4aa;
    SB_LUT4 select_295_Select_0_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n1733), .I2(n18751), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_295_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1392 (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n6_adj_3671), .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(\FRAME_MATCHER.i_31__N_2368 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1392.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(\FRAME_MATCHER.state[2] ), .I1(n6_adj_3671), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n23888));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n31275), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2364 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'h0202;
    SB_LUT4 i2_3_lut_4_lut_adj_1395 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[16] [0]), .I3(\data_in_frame[13] [6]), .O(n30255));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i12878_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n16987));
    defparam i12878_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12812_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n16921));
    defparam i12812_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1396 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n16245));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1396.LUT_INIT = 16'h9696;
    SB_LUT4 i12813_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n16922));
    defparam i12813_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12814_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n16923));
    defparam i12814_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12815_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n16924));
    defparam i12815_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1397 (.I0(n15890), .I1(n15856), .I2(\data_in_frame[6] [4]), 
            .I3(GND_net), .O(n30093));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1397.LUT_INIT = 16'h9696;
    SB_LUT4 i12816_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n16925));
    defparam i12816_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n17116));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12817_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n16926));
    defparam i12817_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12818_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n16927));
    defparam i12818_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12879_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n16988));
    defparam i12879_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12811_3_lut_4_lut (.I0(n8_adj_3819), .I1(n29530), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n16920));
    defparam i12811_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1398 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n29530), .I3(\FRAME_MATCHER.i [0]), .O(n29535));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1398.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1399 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n21151), .I3(\FRAME_MATCHER.i [0]), .O(n29552));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1399.LUT_INIT = 16'hffdf;
    SB_LUT4 equal_72_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3819));   // verilog/coms.v(154[7:23])
    defparam equal_72_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n17115));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14584_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9]_c [6]), 
            .I2(n4216), .I3(GND_net), .O(n16883));
    defparam i14584_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n17114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n17113));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1400 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9][5] ), 
            .I2(\data_in_frame[11] [7]), .I3(n15643), .O(n29666));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n17112));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12880_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n16989));
    defparam i12880_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n17111));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n31247), .D(n59), 
            .R(n30439));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12803_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n16912));
    defparam i12803_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12804_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n16913));
    defparam i12804_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n17110));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12805_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n16914));
    defparam i12805_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12806_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n16915));
    defparam i12806_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n34567_bdd_4_lut (.I0(n34567), .I1(n17_adj_3713), .I2(n16_adj_3712), 
            .I3(byte_transmit_counter[2]), .O(n34570));
    defparam n34567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1401 (.I0(n29733), .I1(n29934), .I2(\data_in_frame[8] [1]), 
            .I3(n29598), .O(n12_adj_3885));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i12807_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n16916));
    defparam i12807_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12808_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n16917));
    defparam i12808_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_29 (.CI(n24890), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n24891));
    SB_LUT4 i12881_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n16990));
    defparam i12881_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_28_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n24889), .O(n2_adj_3733)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14578_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10]_c [2]), 
            .I2(n4216), .I3(GND_net), .O(n16895));
    defparam i14578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12809_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n16918));
    defparam i12809_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12810_3_lut_4_lut (.I0(n8_adj_3813), .I1(n29530), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n16919));
    defparam i12810_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_79_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3813));   // verilog/coms.v(154[7:23])
    defparam equal_79_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_CARRY add_43_28 (.CI(n24889), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n24890));
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_28883 (.I0(byte_transmit_counter[1]), 
            .I1(n33169), .I2(n33170), .I3(byte_transmit_counter[2]), .O(n34561));
    defparam byte_transmit_counter_1__bdd_4_lut_28883.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1402 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n29530), .I3(\FRAME_MATCHER.i [0]), .O(n29532));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1402.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n17109));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1403 (.I0(n15777), .I1(n29707), .I2(\data_in_frame[16] [0]), 
            .I3(\data_in_frame[13] [6]), .O(n6_adj_3779));
    defparam i1_2_lut_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_27_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n24888), .O(n2_adj_3735)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1404 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n21151), .I3(\FRAME_MATCHER.i [0]), .O(n29543));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1404.LUT_INIT = 16'hbfff;
    SB_LUT4 n34561_bdd_4_lut (.I0(n34561), .I1(n17_adj_3711), .I2(n16_adj_3710), 
            .I3(byte_transmit_counter[2]), .O(n34564));
    defparam n34561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n17108));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_27 (.CI(n24888), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n24889));
    SB_LUT4 i1_2_lut_adj_1405 (.I0(n27996), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28050));
    defparam i1_2_lut_adj_1405.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n17107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n17106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n17105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n17104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n17103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n17102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n17101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n17100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n17099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n17098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n17097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n17096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n17095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n17094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n17093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n17092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n17091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n17090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n17089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n17088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n17087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n17086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n17085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n17084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n17083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n17082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n17081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n17080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n17079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n17078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n16865));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n16864));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n16863));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n16862));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n17077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n17076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n17075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n17074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n17073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n17072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n17071));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1406 (.I0(\data_out_frame[24] [1]), .I1(n16054), 
            .I2(n27239), .I3(\data_out_frame[23] [3]), .O(n14_adj_3667));
    defparam i6_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_28878 (.I0(byte_transmit_counter[1]), 
            .I1(n33186), .I2(n33187), .I3(byte_transmit_counter[2]), .O(n34555));
    defparam byte_transmit_counter_1__bdd_4_lut_28878.LUT_INIT = 16'he4aa;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n16853));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n17070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n17069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n17068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n17067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n17066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n17065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n17064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n17063));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n17062));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n17061));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n17060));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n17059));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n17058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n17057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n17056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n17055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n17054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n17053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n17052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n17051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n17050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n17049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n17048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n17047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n17046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n17045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n17044));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n17043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n17042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n17041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n17040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n17039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n17038));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n17037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n17036));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n17035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n17034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n17033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n17032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n17031));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n34555_bdd_4_lut (.I0(n34555), .I1(n17_adj_3697), .I2(n16_adj_3696), 
            .I3(byte_transmit_counter[2]), .O(n34558));
    defparam n34555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n17030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n17029));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n17028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n17027));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n17026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n17025));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n17024));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n17023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n17022));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n17021));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n17020));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n17019));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n17018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n17017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n17016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n17015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n17014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n17013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n17012));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n17011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n17010));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n17009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n17008));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9][0] ), .C(clk32MHz), 
           .D(n17007));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9][1] ), .C(clk32MHz), 
           .D(n17006));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9][2] ), .C(clk32MHz), 
           .D(n17005));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9][3] ), .C(clk32MHz), 
           .D(n17004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9][4] ), .C(clk32MHz), 
           .D(n17003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9][5] ), .C(clk32MHz), 
           .D(n17002));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9]_c [6]), .C(clk32MHz), 
           .D(n17001));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n17000));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1407 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n1519), .I3(n1516), .O(n6_adj_3638));
    defparam i1_2_lut_3_lut_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10]_c [0]), .C(clk32MHz), 
           .D(n16999));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10][1] ), .C(clk32MHz), 
           .D(n16998));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12882_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29549), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n16991));
    defparam i12882_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10]_c [2]), .C(clk32MHz), 
           .D(n16997));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n16996));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n16995));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n16994));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n16993));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n16992));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n16991));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n16990));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n16989));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n16988));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n16987));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n16986));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n16985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n16984));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n16983));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n16982));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n16981));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n16980));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1408 (.I0(\data_in_frame[6] [1]), .I1(n12_adj_3885), 
            .I2(n30093), .I3(n16245), .O(n31783));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n16979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n16978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n16977));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n16976));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n16975));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n16974));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n16973));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n16972));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n16971));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n16970));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n16969));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n16968));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n16967));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n16966));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n16965));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n16964));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n16963));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n16962));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n16961));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n16960));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n16959));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n16958));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n16957));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n16956));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n16955));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_26_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n24887), .O(n2_adj_3737)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n16954));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n16953));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n16952));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_1409 (.I0(n29837), .I1(n31783), .I2(n16011), 
            .I3(n28050), .O(n28_adj_3886));
    defparam i12_4_lut_adj_1409.LUT_INIT = 16'hdfff;
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n16951));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n16950));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n16949));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1410 (.I0(n26741), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[17] [5]), .I3(GND_net), .O(n27067));
    defparam i1_2_lut_3_lut_adj_1410.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_28873 (.I0(byte_transmit_counter[1]), 
            .I1(n33193), .I2(n33194), .I3(byte_transmit_counter[2]), .O(n34549));
    defparam byte_transmit_counter_1__bdd_4_lut_28873.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n1519), .I3(n29572), .O(n24_adj_3814));
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 n34549_bdd_4_lut (.I0(n34549), .I1(n17_adj_3887), .I2(n16_adj_3888), 
            .I3(byte_transmit_counter[2]), .O(n34552));
    defparam n34549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10_4_lut_adj_1411 (.I0(n15768), .I1(n15918), .I2(n7_adj_3802), 
            .I3(n8_adj_3830), .O(n26_adj_3889));
    defparam i10_4_lut_adj_1411.LUT_INIT = 16'hfffb;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n16948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n16947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n16946));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n16945));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n16944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n16943));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_28868 (.I0(byte_transmit_counter[1]), 
            .I1(n33196), .I2(n33197), .I3(byte_transmit_counter[2]), .O(n34543));
    defparam byte_transmit_counter_1__bdd_4_lut_28868.LUT_INIT = 16'he4aa;
    SB_LUT4 i12955_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n17064));
    defparam i12955_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n16942));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n16941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n16940));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12956_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n17065));
    defparam i12956_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_26 (.CI(n24887), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n24888));
    SB_LUT4 i12957_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n17066));
    defparam i12957_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12958_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n17067));
    defparam i12958_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n16939));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n16938));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n16937));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11_4_lut_adj_1412 (.I0(n16333), .I1(n16336), .I2(n16094), 
            .I3(n15914), .O(n27_adj_3890));
    defparam i11_4_lut_adj_1412.LUT_INIT = 16'hfeff;
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n16936));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n16935));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n16934));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n34543_bdd_4_lut (.I0(n34543), .I1(n17_adj_3891), .I2(n16_adj_3892), 
            .I3(byte_transmit_counter[2]), .O(n34546));
    defparam n34543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12959_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n17068));
    defparam i12959_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12960_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n17069));
    defparam i12960_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1413 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[16] [5]), 
            .I2(n27053), .I3(n30133), .O(n6_adj_3629));
    defparam i1_2_lut_3_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1414 (.I0(n26741), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[17] [4]), .I3(\data_out_frame[17] [6]), 
            .O(n30099));
    defparam i2_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i12961_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n17070));
    defparam i12961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12962_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29555), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n17071));
    defparam i12962_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1415 (.I0(n15905), .I1(n16329), .I2(n10_adj_3704), 
            .I3(n15951), .O(n25_adj_3893));
    defparam i9_4_lut_adj_1415.LUT_INIT = 16'hfffe;
    SB_LUT4 i12867_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n16976));
    defparam i12867_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n16933));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n16932));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n16931));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12868_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n16977));
    defparam i12868_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12864_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n16973));
    defparam i12864_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i27803_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33161));
    defparam i27803_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27806_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33160));
    defparam i27806_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12947_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n17056));
    defparam i12947_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n16930));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n16929));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n16928));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n16927));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12948_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n17057));
    defparam i12948_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12949_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n17058));
    defparam i12949_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12950_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n17059));
    defparam i12950_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_25_lut (.I0(n1733), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n24886), .O(n2_adj_3739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n16926));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n16925));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n16924));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n16923));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n16922));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n16921));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12865_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n16974));
    defparam i12865_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12869_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n16978));
    defparam i12869_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12866_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29543), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n16975));
    defparam i12866_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12951_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n17060));
    defparam i12951_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12952_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n17061));
    defparam i12952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12953_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n17062));
    defparam i12953_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12870_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n16979));
    defparam i12870_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12954_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29552), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n17063));
    defparam i12954_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1416 (.I0(\FRAME_MATCHER.state[0] ), .I1(n92), 
            .I2(n18487), .I3(\FRAME_MATCHER.state[2] ), .O(n32159));
    defparam i2_3_lut_4_lut_adj_1416.LUT_INIT = 16'h0e00;
    SB_LUT4 i1_2_lut_3_lut_adj_1417 (.I0(\FRAME_MATCHER.state[0] ), .I1(n92), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(GND_net), .O(n16695));
    defparam i1_2_lut_3_lut_adj_1417.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1418 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n23828), .I3(n21855), .O(n78));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1418.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n23828), .I3(n21855), .O(n31275));
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'hfffe;
    SB_LUT4 i12939_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n17048));
    defparam i12939_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12940_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n17049));
    defparam i12940_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12941_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n17050));
    defparam i12941_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12942_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n17051));
    defparam i12942_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12943_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n17052));
    defparam i12943_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12944_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n17053));
    defparam i12944_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12945_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n17054));
    defparam i12945_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_28863 (.I0(byte_transmit_counter[1]), 
            .I1(n33149), .I2(n33150), .I3(byte_transmit_counter[2]), .O(n34537));
    defparam byte_transmit_counter_1__bdd_4_lut_28863.LUT_INIT = 16'he4aa;
    SB_LUT4 i12946_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29549), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n17055));
    defparam i12946_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n34537_bdd_4_lut (.I0(n34537), .I1(n17_adj_3894), .I2(n16_adj_3895), 
            .I3(byte_transmit_counter[2]), .O(n34540));
    defparam n34537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12931_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n17040));
    defparam i12931_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12932_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n17041));
    defparam i12932_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12933_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n17042));
    defparam i12933_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1420 (.I0(n25_adj_3893), .I1(n27_adj_3890), .I2(n26_adj_3889), 
            .I3(n28_adj_3886), .O(n1));
    defparam i15_4_lut_adj_1420.LUT_INIT = 16'hfffe;
    SB_LUT4 i12934_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n17043));
    defparam i12934_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12935_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n17044));
    defparam i12935_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12936_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n17045));
    defparam i12936_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_28858 (.I0(byte_transmit_counter[1]), 
            .I1(n33152), .I2(n33153), .I3(byte_transmit_counter[2]), .O(n34531));
    defparam byte_transmit_counter_1__bdd_4_lut_28858.LUT_INIT = 16'he4aa;
    SB_LUT4 i12937_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n17046));
    defparam i12937_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12938_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29546), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n17047));
    defparam i12938_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12871_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n16980));
    defparam i12871_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12872_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n16981));
    defparam i12872_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(n23828), .I1(n21855), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(GND_net), .O(n6_adj_3671));
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'hfefe;
    SB_LUT4 i17053_2_lut_3_lut (.I0(n1733), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n21151));
    defparam i17053_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i12873_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n16982));
    defparam i12873_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1422 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3668));
    defparam i2_2_lut_adj_1422.LUT_INIT = 16'h6666;
    SB_LUT4 n34531_bdd_4_lut (.I0(n34531), .I1(n17_adj_3896), .I2(n16_adj_3897), 
            .I3(byte_transmit_counter[2]), .O(n34534));
    defparam n34531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12923_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n17032));
    defparam i12923_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12924_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n17033));
    defparam i12924_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1423 (.I0(n29810), .I1(n29689), .I2(\data_in_frame[8] [2]), 
            .I3(n30096), .O(n10_adj_3898));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1424 (.I0(\data_in_frame[11] [0]), .I1(n7_adj_3802), 
            .I2(GND_net), .I3(GND_net), .O(n16192));
    defparam i1_2_lut_adj_1424.LUT_INIT = 16'h6666;
    SB_LUT4 i12925_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n17034));
    defparam i12925_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n29714));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1426 (.I0(\data_in_frame[16] [0]), .I1(n15947), 
            .I2(\data_in_frame[18] [0]), .I3(n29790), .O(n10_adj_3827));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i12926_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n17035));
    defparam i12926_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12927_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n17036));
    defparam i12927_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12874_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29546), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n16983));
    defparam i12874_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3897));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3896));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27808_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33153));
    defparam i27808_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12928_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n17037));
    defparam i12928_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i27812_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33152));
    defparam i27812_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14595_1_lut (.I0(PWMLimit[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18701));   // verilog/coms.v(127[12] 300[6])
    defparam i14595_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_2_lut_adj_1427 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_3899));   // verilog/coms.v(238[12:32])
    defparam i4_2_lut_adj_1427.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1428 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3900));   // verilog/coms.v(238[12:32])
    defparam i5_4_lut_adj_1428.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_28893 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n34519));
    defparam byte_transmit_counter_0__bdd_4_lut_28893.LUT_INIT = 16'he4aa;
    SB_LUT4 n34519_bdd_4_lut (.I0(n34519), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n34522));
    defparam n34519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1429 (.I0(n13_adj_3900), .I1(\data_in_frame[0] [7]), 
            .I2(n12_adj_3899), .I3(\data_in_frame[0] [5]), .O(n13173));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1429.LUT_INIT = 16'hfffb;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3895));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1430 (.I0(n26989), .I1(\data_out_frame[19] [3]), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[15] [1]), 
            .O(n6_adj_3657));
    defparam i1_2_lut_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i12929_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n17038));
    defparam i12929_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1431 (.I0(n13173), .I1(n1), .I2(GND_net), .I3(GND_net), 
            .O(n19));
    defparam i1_2_lut_adj_1431.LUT_INIT = 16'heeee;
    SB_LUT4 i12930_3_lut_4_lut (.I0(n10_adj_3867), .I1(n29543), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n17039));
    defparam i12930_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1432 (.I0(n16396), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [2]), .I3(n27063), .O(n27977));
    defparam i2_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3894));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27814_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33150));
    defparam i27814_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27816_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33149));
    defparam i27816_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1433 (.I0(n26989), .I1(\data_out_frame[19] [3]), 
            .I2(\data_out_frame[18] [1]), .I3(\data_out_frame[17] [3]), 
            .O(n22_adj_3823));
    defparam i1_2_lut_3_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1434 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(GND_net), .O(n59));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1434.LUT_INIT = 16'h5454;
    SB_LUT4 i28478_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n92), .I3(GND_net), .O(n30439));
    defparam i28478_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_4_lut_adj_1435 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[0] [7]), .O(n16220));
    defparam i1_2_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1436 (.I0(n6_adj_3677), .I1(n21151), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n10_adj_3699), .O(n29541));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_4_lut_adj_1436.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_4_lut_adj_1437 (.I0(n6_adj_3677), .I1(n21151), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n10_adj_3867), .O(n29542));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_4_lut_adj_1437.LUT_INIT = 16'hfff7;
    SB_LUT4 i2_2_lut_3_lut_adj_1438 (.I0(n63_adj_3692), .I1(n63_adj_3689), 
            .I2(n63), .I3(GND_net), .O(n12869));   // verilog/coms.v(139[4] 141[7])
    defparam i2_2_lut_3_lut_adj_1438.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1439 (.I0(n16396), .I1(\data_out_frame[15] [3]), 
            .I2(n27479), .I3(GND_net), .O(n27980));
    defparam i1_2_lut_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_LUT4 i17082_2_lut_3_lut (.I0(n63_adj_3692), .I1(n63_adj_3689), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n33[1]));   // verilog/coms.v(139[4] 141[7])
    defparam i17082_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1440 (.I0(n117), .I1(n67), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(GND_net), .O(n7_adj_3662));
    defparam i1_2_lut_3_lut_adj_1440.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3892));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3891));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1441 (.I0(n23828), .I1(n21855), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state[2] ), .O(n92));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1441.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1442 (.I0(n6_adj_3677), .I1(n21151), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n10_adj_3699), .O(n29538));
    defparam i1_2_lut_4_lut_adj_1442.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_4_lut_adj_1443 (.I0(n6_adj_3677), .I1(n21151), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n10_adj_3867), .O(n29539));
    defparam i1_2_lut_4_lut_adj_1443.LUT_INIT = 16'hff7f;
    SB_LUT4 i28536_3_lut_4_lut (.I0(n63_adj_3), .I1(tx_active), .I2(r_SM_Main_2__N_3360[0]), 
            .I3(\FRAME_MATCHER.i_31__N_2367 ), .O(n16652));
    defparam i28536_3_lut_4_lut.LUT_INIT = 16'h5755;
    SB_LUT4 i27674_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33197));
    defparam i27674_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27668_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33196));
    defparam i27668_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(\FRAME_MATCHER.state[2] ), .I1(n18751), 
            .I2(n29447), .I3(n30_adj_3846), .O(n4216));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'h2000;
    SB_LUT4 i28372_2_lut_3_lut (.I0(n16652), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n23888), .I3(GND_net), .O(n16773));
    defparam i28372_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i1_2_lut_4_lut_adj_1445 (.I0(tx_active), .I1(r_SM_Main_2__N_3360[0]), 
            .I2(byte_transmit_counter[7]), .I3(n4_adj_3672), .O(n884));
    defparam i1_2_lut_4_lut_adj_1445.LUT_INIT = 16'heeef;
    SB_LUT4 i1_2_lut_3_lut_adj_1446 (.I0(n31275), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2370 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1446.LUT_INIT = 16'h4040;
    SB_LUT4 i1543_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_3678));
    defparam i1543_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 equal_66_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3820));
    defparam equal_66_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_4_lut_adj_1447 (.I0(n23888), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n18751), .I3(n63_adj_3), .O(n89));   // verilog/coms.v(112[11:16])
    defparam i1_2_lut_4_lut_adj_1447.LUT_INIT = 16'haeff;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n15542), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_3666));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 equal_67_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3669));
    defparam equal_67_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_4_lut_adj_1448 (.I0(\FRAME_MATCHER.state[3] ), .I1(n12869), 
            .I2(n2329), .I3(n2_adj_3695), .O(n28941));
    defparam i1_3_lut_4_lut_adj_1448.LUT_INIT = 16'haa80;
    SB_LUT4 i12899_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n17008));
    defparam i12899_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1449 (.I0(\FRAME_MATCHER.state[0] ), .I1(n23888), 
            .I2(n21130), .I3(tx_transmit_N_3257), .O(n2));
    defparam i1_2_lut_4_lut_adj_1449.LUT_INIT = 16'h8880;
    SB_LUT4 i2_3_lut_4_lut_adj_1450 (.I0(n27050), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[16] [6]), .I3(n16592), .O(n30139));
    defparam i2_3_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i12900_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n17009));
    defparam i12900_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3888));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3887));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27783_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33194));
    defparam i27783_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12901_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n17010));
    defparam i12901_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12902_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n17011));
    defparam i12902_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i27532_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33193));
    defparam i27532_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1451 (.I0(\data_out_frame[12] [5]), .I1(n1519), 
            .I2(\data_out_frame[14] [4]), .I3(\data_out_frame[14] [3]), 
            .O(n16592));
    defparam i1_2_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1452 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n30087));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n33478));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3901));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12903_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n17012));
    defparam i12903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1453 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n6_adj_3654));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1453.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_4_lut (.I0(n5_adj_3901), 
            .I1(byte_transmit_counter[0]), .I2(n33045), .I3(n33478), .O(n7_adj_3879));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1813749_i1_3_lut (.I0(n34588), .I1(n34690), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3878));
    defparam i1813749_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1454 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n30002));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_LUT4 i27774_2_lut (.I0(n34738), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33159));
    defparam i27774_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12904_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n17013));
    defparam i12904_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3902));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3903));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut (.I0(n5_adj_3903), 
            .I1(n6_adj_3902), .I2(n33045), .I3(GND_net), .O(n7_adj_3877));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12905_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n17014));
    defparam i12905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12906_3_lut_4_lut (.I0(n10_adj_3699), .I1(n29558), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n17015));
    defparam i12906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1814352_i1_3_lut (.I0(n34582), .I1(n34762), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3876));
    defparam i1814352_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27771_2_lut (.I0(n34744), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33165));
    defparam i27771_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3904));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3905));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut (.I0(n5_adj_3905), 
            .I1(n6_adj_3904), .I2(n33045), .I3(GND_net), .O(n7_adj_3875));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1455 (.I0(n117), .I1(n67), .I2(n115), .I3(\FRAME_MATCHER.state [13]), 
            .O(n8_adj_3715));
    defparam i1_2_lut_4_lut_adj_1455.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1456 (.I0(n117), .I1(n67), .I2(n115), .I3(\FRAME_MATCHER.state [14]), 
            .O(n8_adj_3714));
    defparam i1_2_lut_4_lut_adj_1456.LUT_INIT = 16'hfe00;
    SB_LUT4 i1814955_i1_3_lut (.I0(n34522), .I1(n34780), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3874));
    defparam i1814955_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27799_2_lut (.I0(n34750), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33168));
    defparam i27799_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3906));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha003;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3907));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut (.I0(n5_adj_3907), 
            .I1(n6_adj_3906), .I2(n33045), .I3(GND_net), .O(n7_adj_3873));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1815558_i1_3_lut (.I0(n34672), .I1(n34786), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3872));
    defparam i1815558_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27795_2_lut (.I0(n34756), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33171));
    defparam i27795_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1457 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[9] [4]), .O(n29644));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_4_lut (.I0(n29627), .I1(n29996), .I2(\data_out_frame[9] [5]), 
            .I3(\data_out_frame[14] [2]), .O(n10_adj_3636));   // verilog/coms.v(71[16:27])
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1458 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[10] [4]), 
            .I2(n1380), .I3(GND_net), .O(n6_adj_3633));
    defparam i1_2_lut_3_lut_adj_1458.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1459 (.I0(n2329), .I1(n2), .I2(n3303), 
            .I3(\FRAME_MATCHER.i_31__N_2368 ), .O(n6));
    defparam i2_3_lut_4_lut_adj_1459.LUT_INIT = 16'hefee;
    SB_LUT4 i3_4_lut_3_lut_4_lut (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[5] [4]), .O(n30170));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_2_lut_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(n29639), .I3(GND_net), .O(n36));
    defparam i9_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(n16034), .I1(\data_out_frame[13] [3]), 
            .I2(n15366), .I3(GND_net), .O(n26741));
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1461 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n29777));
    defparam i1_2_lut_3_lut_adj_1461.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1462 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(n10_adj_3616), .I3(\data_out_frame[6] [6]), .O(n16396));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1463 (.I0(\data_out_frame[23] [4]), .I1(n13916), 
            .I2(n27952), .I3(\data_out_frame[23] [2]), .O(n6_adj_3630));
    defparam i1_2_lut_4_lut_adj_1463.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1464 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[18] [0]), 
            .I2(n27980), .I3(n29816), .O(n29751));
    defparam i1_3_lut_4_lut_adj_1464.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1465 (.I0(\data_out_frame[13] [3]), .I1(n16396), 
            .I2(\data_out_frame[15] [4]), .I3(n15366), .O(n29816));
    defparam i2_3_lut_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1466 (.I0(n27019), .I1(\data_out_frame[23] [3]), 
            .I2(n30102), .I3(n27930), .O(n15291));
    defparam i2_3_lut_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1467 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(n10_adj_3898), .I3(\data_in_frame[5] [6]), .O(n15951));   // verilog/coms.v(78[16:27])
    defparam i5_3_lut_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1468 (.I0(n27980), .I1(n29816), .I2(n30222), 
            .I3(GND_net), .O(n6_adj_3609));
    defparam i1_2_lut_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1469 (.I0(n28046), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[25] [2]), .I3(n29584), .O(n29974));
    defparam i2_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1470 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[20] [2]), 
            .I2(n29654), .I3(\data_out_frame[18] [0]), .O(n6_c));
    defparam i1_2_lut_4_lut_adj_1470.LUT_INIT = 16'h6996;
    uart_tx tx (.clk32MHz(clk32MHz), .\r_SM_Main_2__N_3360[0] (r_SM_Main_2__N_3360[0]), 
            .r_SM_Main({Open_10, \r_SM_Main[1] , Open_11}), .GND_net(GND_net), 
            .tx_o(tx_o), .tx_data({tx_data}), .VCC_net(VCC_net), .n4(n4), 
            .n16871(n16871), .tx_active(tx_active), .n8947(n8947), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.n16710(n16710), .clk32MHz(clk32MHz), .n16802(n16802), 
            .GND_net(GND_net), .n21215(n21215), .n4(n4_adj_4), .r_Rx_Data(r_Rx_Data), 
            .n4_adj_1(n4_adj_5), .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n15595(n15595), 
            .RX_N_2(RX_N_2), .VCC_net(VCC_net), .n15590(n15590), .n4_adj_2(n4_adj_6), 
            .n17376(n17376), .rx_data_ready(rx_data_ready), .n17380(n17380), 
            .rx_data({rx_data}), .n16861(n16861), .n16860(n16860), .n16859(n16859), 
            .n16858(n16858), .n16857(n16857), .n16856(n16856), .n16855(n16855)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, \r_SM_Main_2__N_3360[0] , r_SM_Main, GND_net, 
            tx_o, tx_data, VCC_net, n4, n16871, tx_active, n8947, 
            tx_enable) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    input \r_SM_Main_2__N_3360[0] ;
    output [2:0]r_SM_Main;
    input GND_net;
    output tx_o;
    input [7:0]tx_data;
    input VCC_net;
    output n4;
    input n16871;
    output tx_active;
    output n8947;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n307;
    
    wire n16716;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n24336;
    wire [8:0]n41;
    
    wire n4140;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n16785, n44, n24370, n22;
    wire [2:0]r_SM_Main_c;   // verilog/uart_tx.v(31[16:25])
    
    wire n10738, n34720, n34606, o_Tx_Serial_N_3388, n3, n12936;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n10, n31194, n25576, n25575, n25574, n25573, n25572, 
        n25571, n25570, n25569, n30755, n34717, n3_adj_3605, n34603, 
        n29251;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n16716), 
            .D(n307[2]), .R(n24336));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n16716), 
            .D(n307[1]), .R(n24336));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1130__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n4140), .D(n41[4]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1130__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n4140), .D(n41[3]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1130__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n4140), .D(n41[2]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1130__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n4140), .D(n41[1]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i24_4_lut (.I0(\r_SM_Main_2__N_3360[0] ), .I1(n44), .I2(r_SM_Main[1]), 
            .I3(n24370), .O(n22));   // verilog/uart_tx.v(31[16:25])
    defparam i24_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i25_3_lut (.I0(n22), .I1(n24370), .I2(r_SM_Main_c[0]), .I3(GND_net), 
            .O(n10738));   // verilog/uart_tx.v(31[16:25])
    defparam i25_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1816764_i1_3_lut (.I0(n34720), .I1(n34606), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3388));
    defparam i1816764_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main_c[0]), .I1(o_Tx_Serial_N_3388), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n4140), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n10738), 
            .R(r_SM_Main_c[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1130__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n4140), .D(n41[5]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1058_1_lut (.I0(r_SM_Main_c[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4140));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1058_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(33[16:27])
    defparam i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[4]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[5]), .I1(n10), .I2(r_Clock_Count[2]), 
            .I3(GND_net), .O(n31194));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[8]), 
            .I3(n31194), .O(n24370));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n44));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut (.I0(r_SM_Main[1]), .I1(n16716), .I2(n44), .I3(GND_net), 
            .O(n24336));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main_c[0]), .I1(r_SM_Main_c[2]), .I2(r_SM_Main[1]), 
            .I3(n24370), .O(n16716));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i20300_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(33[16:27])
    defparam i20300_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 r_Clock_Count_1130_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n25576), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1130_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n25575), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_9 (.CI(n25575), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n25576));
    SB_LUT4 r_Clock_Count_1130_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n25574), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_8 (.CI(n25574), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n25575));
    SB_LUT4 r_Clock_Count_1130_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n25573), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_7 (.CI(n25573), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n25574));
    SB_LUT4 r_Clock_Count_1130_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n25572), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_6 (.CI(n25572), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n25573));
    SB_LUT4 r_Clock_Count_1130_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n25571), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_5 (.CI(n25571), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n25572));
    SB_LUT4 r_Clock_Count_1130_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n25570), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_4 (.CI(n25570), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n25571));
    SB_LUT4 r_Clock_Count_1130_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n25569), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_3 (.CI(n25569), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n25570));
    SB_LUT4 r_Clock_Count_1130_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n25569));
    SB_DFFESR r_Clock_Count_1130__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n4140), .D(n41[0]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i3_3_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), 
            .I2(r_SM_Main_c[2]), .I3(\r_SM_Main_2__N_3360[0] ), .O(n12936));
    defparam i3_3_lut_4_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(r_SM_Main_c[0]), .I1(n24370), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_c[2]), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(r_SM_Main_c[0]), .I1(n24370), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_c[2]), .O(n30755));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n34717));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n34717_bdd_4_lut (.I0(n34717), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n34720));
    defparam n34717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i26_2_lut_3_lut (.I0(r_SM_Main_c[0]), .I1(n24370), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3_adj_3605));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i26_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_29006 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n34603));
    defparam r_Bit_Index_0__bdd_4_lut_29006.LUT_INIT = 16'he4aa;
    SB_LUT4 n34603_bdd_4_lut (.I0(n34603), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n34606));
    defparam n34603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR r_Clock_Count_1130__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n4140), .D(n41[6]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n12936), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3605), 
            .R(r_SM_Main_c[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n16871));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n29251));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i12_3_lut (.I0(n16716), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n29251));   // verilog/uart_tx.v(31[16:25])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 i4921_2_lut (.I0(\r_SM_Main_2__N_3360[0] ), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n8947));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i4921_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR r_Clock_Count_1130__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n4140), .D(n41[8]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1130__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n4140), .D(n41[7]), .R(n16785));   // verilog/uart_tx.v(118[34:51])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main_c[2]), .C(clk32MHz), .D(n30755));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i28407_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), 
            .I2(n24370), .I3(r_SM_Main_c[2]), .O(n16785));
    defparam i28407_3_lut_4_lut.LUT_INIT = 16'h00f1;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n16710, clk32MHz, n16802, GND_net, n21215, n4, r_Rx_Data, 
            n4_adj_1, \r_Bit_Index[0] , n15595, RX_N_2, VCC_net, n15590, 
            n4_adj_2, n17376, rx_data_ready, n17380, rx_data, n16861, 
            n16860, n16859, n16858, n16857, n16856, n16855) /* synthesis syn_module_defined=1 */ ;
    output n16710;
    input clk32MHz;
    output n16802;
    input GND_net;
    output n21215;
    output n4;
    output r_Rx_Data;
    output n4_adj_1;
    output \r_Bit_Index[0] ;
    output n15595;
    input RX_N_2;
    input VCC_net;
    output n15590;
    output n4_adj_2;
    input n17376;
    output rx_data_ready;
    input n17380;
    output [7:0]rx_data;
    input n16861;
    input n16860;
    input n16859;
    input n16858;
    input n16857;
    input n16856;
    input n16855;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [7:0]n37;
    
    wire n16700;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n16783;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n19135, n19143, n21803;
    wire [2:0]r_SM_Main_2__N_3286;
    
    wire n2, n19148, n19149, n29508, r_Rx_Data_R, n15441, n31, 
        n5, n8, n6, n25568, n25567, n25566, n25565, n25564, 
        n25563, n25562, n3, n29205, n16659, n21933;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n16710), 
            .D(n326[2]), .R(n16802));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n16710), 
            .D(n326[1]), .R(n16802));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1128__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n16700), .D(n37[7]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1128__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n16700), .D(n37[6]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1128__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n16700), .D(n37[5]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1128__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n16700), .D(n37[4]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1128__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n16700), .D(n37[3]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(n19135), .I2(GND_net), .I3(GND_net), 
            .O(n19143));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n21803), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main_2__N_3286[2]), .I3(GND_net), .O(n2));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'h2c2c;
    SB_LUT4 i15046_3_lut (.I0(n19148), .I1(n2), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n19149));   // verilog/uart_rx.v(36[17:26])
    defparam i15046_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_1128__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n16700), .D(n37[2]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1128__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n16700), .D(n37[1]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3286[2]), 
            .R(n29508));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i17117_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n21215));
    defparam i17117_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_94_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_94_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n19149), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 equal_97_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_97_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_833 (.I0(n15441), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n15595));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_833.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_2));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i3_4_lut (.I0(n31), .I1(r_Clock_Count[5]), .I2(r_Clock_Count[2]), 
            .I3(n5), .O(n19135));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i12674_3_lut (.I0(n16700), .I1(r_SM_Main[2]), .I2(n8), .I3(GND_net), 
            .O(n16783));   // verilog/uart_rx.v(120[34:51])
    defparam i12674_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_2_lut (.I0(n19135), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/uart_rx.v(36[17:26])
    defparam i2_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n6), .I3(r_Rx_Data), 
            .O(n16700));   // verilog/uart_rx.v(36[17:26])
    defparam i1_4_lut.LUT_INIT = 16'h3233;
    SB_LUT4 i1191_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1191_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_834 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(r_Clock_Count[4]), .I3(r_Clock_Count[3]), .O(n5));
    defparam i3_4_lut_adj_834.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_835 (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(120[34:51])
    defparam i1_2_lut_adj_835.LUT_INIT = 16'heeee;
    SB_LUT4 i17713_4_lut (.I0(r_Clock_Count[5]), .I1(n31), .I2(r_Clock_Count[2]), 
            .I3(n5), .O(r_SM_Main_2__N_3286[2]));
    defparam i17713_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n21803));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i12693_3_lut (.I0(n16710), .I1(n21803), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n16802));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12693_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3286[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n16710));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1198_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1198_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 r_Clock_Count_1128_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n25568), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1128_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n25567), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1128_add_4_8 (.CI(n25567), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n25568));
    SB_LUT4 r_Clock_Count_1128_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n25566), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1128_add_4_7 (.CI(n25566), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n25567));
    SB_LUT4 r_Clock_Count_1128_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n25565), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1128_add_4_6 (.CI(n25565), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n25566));
    SB_LUT4 r_Clock_Count_1128_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n25564), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1128_add_4_5 (.CI(n25564), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n25565));
    SB_LUT4 r_Clock_Count_1128_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n25563), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1128_add_4_4 (.CI(n25563), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n25564));
    SB_LUT4 r_Clock_Count_1128_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n25562), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1128_add_4_3 (.CI(n25562), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n25563));
    SB_LUT4 r_Clock_Count_1128_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1128_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1128_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n25562));
    SB_DFFESR r_Clock_Count_1128__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n16700), .D(n37[0]), .R(n16783));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i15045_3_lut_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n19135), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n19148));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15045_3_lut_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_4_lut_adj_836 (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3286[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n15441));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i2_4_lut_adj_836.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_adj_837 (.I0(\r_Bit_Index[0] ), .I1(n15441), .I2(GND_net), 
            .I3(GND_net), .O(n15590));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_837.LUT_INIT = 16'heeee;
    SB_LUT4 equal_98_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_98_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n17376));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n29205));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n17380));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n16861));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n16860));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n16859));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n16858));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n16857));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n16856));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n16855));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i19_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n19135), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3286[2]), .O(n8));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i19_3_lut_4_lut.LUT_INIT = 16'h08f8;
    SB_LUT4 i21_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3286[2]), 
            .I3(r_SM_Main[0]), .O(n16659));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i21_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n16659), 
            .I3(rx_data_ready), .O(n29205));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i28540_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n29508));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i28540_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i17832_2_lut (.I0(r_SM_Main_2__N_3286[2]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n21933));
    defparam i17832_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15042_4_lut (.I0(r_Rx_Data), .I1(n21933), .I2(r_SM_Main[1]), 
            .I3(n19143), .O(n3));   // verilog/uart_rx.v(36[17:26])
    defparam i15042_4_lut.LUT_INIT = 16'h3530;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n33856, VCC_net, INHA_c, clk32MHz, n15455, pwm_counter, 
            GND_net, n15453) /* synthesis syn_module_defined=1 */ ;
    input n33856;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n15455;
    output [31:0]pwm_counter;
    input GND_net;
    input n15453;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n31299, n18, n24, n22, n26, n21, pwm_counter_31__N_555;
    wire [31:0]n133;
    
    wire n25561, n25560, n25559, n25558, n25557, n25556, n25555, 
        n25554, n25553, n25552, n25551, n25550, n25549, n25548, 
        n25547, n25546, n25545, n25544, n25543, n25542, n25541, 
        n25540, n25539, n25538, n25537, n25536, n25535, n25534, 
        n25533, n25532, n25531;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n33856), 
            .R(n15455));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n31299));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n31299), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n18));
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[22]), .I2(pwm_counter[14]), 
            .I3(pwm_counter[18]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(pwm_counter[21]), .I1(n15453), .I2(pwm_counter[16]), 
            .I3(pwm_counter[12]), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(pwm_counter[15]), .I1(n24), .I2(n18), .I3(pwm_counter[19]), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_2_lut (.I0(pwm_counter[11]), .I1(pwm_counter[20]), .I2(GND_net), 
            .I3(GND_net), .O(n21));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i17129_4_lut (.I0(n21), .I1(pwm_counter[31]), .I2(n26), .I3(n22), 
            .O(pwm_counter_31__N_555));   // verilog/pwm.v(18[8:40])
    defparam i17129_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 pwm_counter_1126_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[31]), 
            .I3(n25561), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1126_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n25560), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_32 (.CI(n25560), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n25561));
    SB_LUT4 pwm_counter_1126_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n25559), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_31 (.CI(n25559), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n25560));
    SB_LUT4 pwm_counter_1126_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n25558), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_30 (.CI(n25558), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n25559));
    SB_LUT4 pwm_counter_1126_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n25557), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_29 (.CI(n25557), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n25558));
    SB_LUT4 pwm_counter_1126_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n25556), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_28 (.CI(n25556), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n25557));
    SB_LUT4 pwm_counter_1126_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n25555), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_27 (.CI(n25555), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n25556));
    SB_LUT4 pwm_counter_1126_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n25554), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_26 (.CI(n25554), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n25555));
    SB_LUT4 pwm_counter_1126_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n25553), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_25 (.CI(n25553), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n25554));
    SB_LUT4 pwm_counter_1126_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n25552), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_24 (.CI(n25552), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n25553));
    SB_LUT4 pwm_counter_1126_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n25551), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_23 (.CI(n25551), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n25552));
    SB_LUT4 pwm_counter_1126_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n25550), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_22 (.CI(n25550), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n25551));
    SB_LUT4 pwm_counter_1126_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n25549), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_21 (.CI(n25549), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n25550));
    SB_LUT4 pwm_counter_1126_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n25548), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_20 (.CI(n25548), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n25549));
    SB_LUT4 pwm_counter_1126_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n25547), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_19 (.CI(n25547), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n25548));
    SB_LUT4 pwm_counter_1126_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n25546), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_18 (.CI(n25546), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n25547));
    SB_LUT4 pwm_counter_1126_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n25545), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_17 (.CI(n25545), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n25546));
    SB_LUT4 pwm_counter_1126_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n25544), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_16 (.CI(n25544), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n25545));
    SB_LUT4 pwm_counter_1126_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n25543), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_15 (.CI(n25543), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n25544));
    SB_LUT4 pwm_counter_1126_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n25542), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_14 (.CI(n25542), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n25543));
    SB_LUT4 pwm_counter_1126_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n25541), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_13 (.CI(n25541), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n25542));
    SB_LUT4 pwm_counter_1126_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n25540), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_12 (.CI(n25540), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n25541));
    SB_LUT4 pwm_counter_1126_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n25539), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_11 (.CI(n25539), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n25540));
    SB_LUT4 pwm_counter_1126_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n25538), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_10 (.CI(n25538), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n25539));
    SB_LUT4 pwm_counter_1126_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n25537), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_9 (.CI(n25537), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n25538));
    SB_LUT4 pwm_counter_1126_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n25536), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_8 (.CI(n25536), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n25537));
    SB_LUT4 pwm_counter_1126_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n25535), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_7 (.CI(n25535), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n25536));
    SB_LUT4 pwm_counter_1126_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n25534), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_6 (.CI(n25534), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n25535));
    SB_LUT4 pwm_counter_1126_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n25533), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_5 (.CI(n25533), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n25534));
    SB_LUT4 pwm_counter_1126_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n25532), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_4 (.CI(n25532), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n25533));
    SB_LUT4 pwm_counter_1126_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n25531), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_3 (.CI(n25531), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n25532));
    SB_LUT4 pwm_counter_1126_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1126_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1126_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n25531));
    SB_DFFSR pwm_counter_1126__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n133[10]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n133[11]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n133[12]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n133[13]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n133[14]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n133[15]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n133[16]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n133[17]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n133[18]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n133[19]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n133[20]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n133[21]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n133[22]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1126__i31 (.Q(pwm_counter[31]), .C(clk32MHz), .D(n133[31]), 
            .R(pwm_counter_31__N_555));   // verilog/pwm.v(17[20:33])
    
endmodule
