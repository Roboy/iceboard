// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jan 29 2020 18:32:34

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    output USBPU;
    output TX;
    inout SDA;
    inout SCL;
    input RX;
    output NEOPXL;
    output LED;
    output INLC;
    output INLB;
    output INLA;
    output INHC;
    output INHB;
    output INHA;
    input HALL3;
    input HALL2;
    input HALL1;
    input FAULT_N;
    input ENCODER1_B;
    input ENCODER1_A;
    input ENCODER0_B;
    input ENCODER0_A;
    output DE;
    input CS_MISO;
    output CS_CLK;
    output CS;
    input CLK;

    wire N__30138;
    wire N__30137;
    wire N__30136;
    wire N__30129;
    wire N__30128;
    wire N__30127;
    wire N__30120;
    wire N__30119;
    wire N__30118;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30102;
    wire N__30101;
    wire N__30100;
    wire N__30093;
    wire N__30092;
    wire N__30091;
    wire N__30084;
    wire N__30083;
    wire N__30082;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30066;
    wire N__30065;
    wire N__30064;
    wire N__30057;
    wire N__30056;
    wire N__30055;
    wire N__30048;
    wire N__30047;
    wire N__30046;
    wire N__30039;
    wire N__30038;
    wire N__30037;
    wire N__30030;
    wire N__30029;
    wire N__30028;
    wire N__30021;
    wire N__30020;
    wire N__30019;
    wire N__30012;
    wire N__30011;
    wire N__30010;
    wire N__30003;
    wire N__30002;
    wire N__30001;
    wire N__29984;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29962;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29930;
    wire N__29927;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29915;
    wire N__29912;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29900;
    wire N__29897;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29867;
    wire N__29866;
    wire N__29865;
    wire N__29864;
    wire N__29863;
    wire N__29862;
    wire N__29861;
    wire N__29860;
    wire N__29859;
    wire N__29858;
    wire N__29857;
    wire N__29856;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29817;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29805;
    wire N__29798;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29786;
    wire N__29785;
    wire N__29782;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29764;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29716;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29695;
    wire N__29694;
    wire N__29693;
    wire N__29690;
    wire N__29689;
    wire N__29688;
    wire N__29687;
    wire N__29684;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29658;
    wire N__29657;
    wire N__29656;
    wire N__29651;
    wire N__29646;
    wire N__29641;
    wire N__29636;
    wire N__29633;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29625;
    wire N__29624;
    wire N__29619;
    wire N__29616;
    wire N__29611;
    wire N__29608;
    wire N__29603;
    wire N__29598;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29545;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29496;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29458;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29394;
    wire N__29391;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29304;
    wire N__29299;
    wire N__29296;
    wire N__29291;
    wire N__29288;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29276;
    wire N__29273;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29252;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29212;
    wire N__29211;
    wire N__29210;
    wire N__29209;
    wire N__29208;
    wire N__29207;
    wire N__29206;
    wire N__29205;
    wire N__29204;
    wire N__29203;
    wire N__29200;
    wire N__29199;
    wire N__29198;
    wire N__29187;
    wire N__29186;
    wire N__29185;
    wire N__29184;
    wire N__29181;
    wire N__29180;
    wire N__29179;
    wire N__29178;
    wire N__29177;
    wire N__29176;
    wire N__29175;
    wire N__29174;
    wire N__29173;
    wire N__29172;
    wire N__29171;
    wire N__29170;
    wire N__29169;
    wire N__29168;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29124;
    wire N__29117;
    wire N__29112;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29098;
    wire N__29097;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29091;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29061;
    wire N__29054;
    wire N__29049;
    wire N__29044;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29010;
    wire N__29001;
    wire N__28998;
    wire N__28985;
    wire N__28982;
    wire N__28981;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28967;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28933;
    wire N__28932;
    wire N__28931;
    wire N__28930;
    wire N__28929;
    wire N__28928;
    wire N__28927;
    wire N__28926;
    wire N__28925;
    wire N__28924;
    wire N__28923;
    wire N__28922;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28916;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28908;
    wire N__28905;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28897;
    wire N__28896;
    wire N__28893;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28884;
    wire N__28883;
    wire N__28882;
    wire N__28879;
    wire N__28878;
    wire N__28877;
    wire N__28876;
    wire N__28875;
    wire N__28874;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28845;
    wire N__28844;
    wire N__28843;
    wire N__28842;
    wire N__28841;
    wire N__28838;
    wire N__28833;
    wire N__28824;
    wire N__28815;
    wire N__28808;
    wire N__28803;
    wire N__28792;
    wire N__28785;
    wire N__28784;
    wire N__28783;
    wire N__28782;
    wire N__28781;
    wire N__28778;
    wire N__28777;
    wire N__28774;
    wire N__28773;
    wire N__28772;
    wire N__28771;
    wire N__28770;
    wire N__28769;
    wire N__28768;
    wire N__28767;
    wire N__28766;
    wire N__28765;
    wire N__28764;
    wire N__28763;
    wire N__28762;
    wire N__28761;
    wire N__28760;
    wire N__28759;
    wire N__28756;
    wire N__28747;
    wire N__28738;
    wire N__28737;
    wire N__28734;
    wire N__28733;
    wire N__28730;
    wire N__28729;
    wire N__28726;
    wire N__28725;
    wire N__28722;
    wire N__28721;
    wire N__28718;
    wire N__28717;
    wire N__28716;
    wire N__28715;
    wire N__28714;
    wire N__28713;
    wire N__28712;
    wire N__28711;
    wire N__28710;
    wire N__28709;
    wire N__28708;
    wire N__28699;
    wire N__28690;
    wire N__28685;
    wire N__28676;
    wire N__28669;
    wire N__28660;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28634;
    wire N__28633;
    wire N__28632;
    wire N__28625;
    wire N__28616;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28600;
    wire N__28599;
    wire N__28596;
    wire N__28595;
    wire N__28594;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28563;
    wire N__28562;
    wire N__28561;
    wire N__28560;
    wire N__28559;
    wire N__28558;
    wire N__28557;
    wire N__28556;
    wire N__28555;
    wire N__28554;
    wire N__28553;
    wire N__28552;
    wire N__28551;
    wire N__28550;
    wire N__28549;
    wire N__28548;
    wire N__28547;
    wire N__28546;
    wire N__28545;
    wire N__28544;
    wire N__28543;
    wire N__28540;
    wire N__28539;
    wire N__28538;
    wire N__28537;
    wire N__28524;
    wire N__28517;
    wire N__28506;
    wire N__28505;
    wire N__28504;
    wire N__28501;
    wire N__28500;
    wire N__28489;
    wire N__28480;
    wire N__28479;
    wire N__28478;
    wire N__28477;
    wire N__28474;
    wire N__28469;
    wire N__28460;
    wire N__28451;
    wire N__28446;
    wire N__28441;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28433;
    wire N__28430;
    wire N__28429;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28411;
    wire N__28408;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28392;
    wire N__28391;
    wire N__28390;
    wire N__28387;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28379;
    wire N__28376;
    wire N__28375;
    wire N__28372;
    wire N__28371;
    wire N__28370;
    wire N__28367;
    wire N__28366;
    wire N__28365;
    wire N__28362;
    wire N__28357;
    wire N__28356;
    wire N__28353;
    wire N__28352;
    wire N__28345;
    wire N__28340;
    wire N__28335;
    wire N__28330;
    wire N__28325;
    wire N__28320;
    wire N__28319;
    wire N__28318;
    wire N__28311;
    wire N__28306;
    wire N__28303;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28291;
    wire N__28290;
    wire N__28289;
    wire N__28288;
    wire N__28287;
    wire N__28278;
    wire N__28269;
    wire N__28268;
    wire N__28265;
    wire N__28264;
    wire N__28261;
    wire N__28252;
    wire N__28247;
    wire N__28244;
    wire N__28243;
    wire N__28242;
    wire N__28237;
    wire N__28230;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28204;
    wire N__28199;
    wire N__28194;
    wire N__28191;
    wire N__28190;
    wire N__28185;
    wire N__28178;
    wire N__28175;
    wire N__28170;
    wire N__28169;
    wire N__28164;
    wire N__28161;
    wire N__28154;
    wire N__28153;
    wire N__28150;
    wire N__28149;
    wire N__28146;
    wire N__28145;
    wire N__28142;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28134;
    wire N__28129;
    wire N__28122;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28105;
    wire N__28104;
    wire N__28103;
    wire N__28090;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28058;
    wire N__28055;
    wire N__28048;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28032;
    wire N__28031;
    wire N__28026;
    wire N__28021;
    wire N__28016;
    wire N__28015;
    wire N__28012;
    wire N__28011;
    wire N__28008;
    wire N__28007;
    wire N__28004;
    wire N__28003;
    wire N__28000;
    wire N__27993;
    wire N__27988;
    wire N__27985;
    wire N__27970;
    wire N__27965;
    wire N__27960;
    wire N__27957;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27931;
    wire N__27926;
    wire N__27919;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27884;
    wire N__27881;
    wire N__27880;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27844;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27823;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27794;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27782;
    wire N__27779;
    wire N__27778;
    wire N__27775;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27742;
    wire N__27741;
    wire N__27738;
    wire N__27733;
    wire N__27728;
    wire N__27725;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27655;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27638;
    wire N__27637;
    wire N__27636;
    wire N__27635;
    wire N__27632;
    wire N__27631;
    wire N__27624;
    wire N__27619;
    wire N__27614;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27581;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27538;
    wire N__27535;
    wire N__27528;
    wire N__27527;
    wire N__27526;
    wire N__27525;
    wire N__27524;
    wire N__27523;
    wire N__27522;
    wire N__27521;
    wire N__27520;
    wire N__27517;
    wire N__27516;
    wire N__27515;
    wire N__27514;
    wire N__27513;
    wire N__27508;
    wire N__27503;
    wire N__27496;
    wire N__27495;
    wire N__27494;
    wire N__27493;
    wire N__27490;
    wire N__27485;
    wire N__27482;
    wire N__27475;
    wire N__27472;
    wire N__27465;
    wire N__27456;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27425;
    wire N__27424;
    wire N__27423;
    wire N__27420;
    wire N__27419;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27411;
    wire N__27410;
    wire N__27409;
    wire N__27408;
    wire N__27407;
    wire N__27406;
    wire N__27405;
    wire N__27404;
    wire N__27403;
    wire N__27402;
    wire N__27401;
    wire N__27400;
    wire N__27397;
    wire N__27390;
    wire N__27387;
    wire N__27386;
    wire N__27385;
    wire N__27382;
    wire N__27375;
    wire N__27370;
    wire N__27369;
    wire N__27368;
    wire N__27367;
    wire N__27364;
    wire N__27353;
    wire N__27348;
    wire N__27345;
    wire N__27340;
    wire N__27333;
    wire N__27326;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27175;
    wire N__27174;
    wire N__27171;
    wire N__27166;
    wire N__27161;
    wire N__27160;
    wire N__27159;
    wire N__27158;
    wire N__27157;
    wire N__27154;
    wire N__27153;
    wire N__27152;
    wire N__27151;
    wire N__27150;
    wire N__27149;
    wire N__27148;
    wire N__27145;
    wire N__27144;
    wire N__27143;
    wire N__27142;
    wire N__27139;
    wire N__27138;
    wire N__27133;
    wire N__27132;
    wire N__27131;
    wire N__27130;
    wire N__27129;
    wire N__27126;
    wire N__27119;
    wire N__27112;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27096;
    wire N__27093;
    wire N__27084;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27037;
    wire N__27036;
    wire N__27033;
    wire N__27032;
    wire N__27029;
    wire N__27028;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__26993;
    wire N__26990;
    wire N__26989;
    wire N__26988;
    wire N__26987;
    wire N__26986;
    wire N__26983;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26951;
    wire N__26950;
    wire N__26949;
    wire N__26948;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26927;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26896;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26892;
    wire N__26891;
    wire N__26888;
    wire N__26887;
    wire N__26886;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26854;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26840;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26828;
    wire N__26825;
    wire N__26820;
    wire N__26819;
    wire N__26818;
    wire N__26817;
    wire N__26816;
    wire N__26815;
    wire N__26812;
    wire N__26807;
    wire N__26798;
    wire N__26795;
    wire N__26790;
    wire N__26785;
    wire N__26782;
    wire N__26775;
    wire N__26772;
    wire N__26753;
    wire N__26752;
    wire N__26747;
    wire N__26744;
    wire N__26743;
    wire N__26742;
    wire N__26741;
    wire N__26740;
    wire N__26739;
    wire N__26738;
    wire N__26737;
    wire N__26736;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26724;
    wire N__26721;
    wire N__26720;
    wire N__26717;
    wire N__26716;
    wire N__26713;
    wire N__26712;
    wire N__26709;
    wire N__26708;
    wire N__26699;
    wire N__26694;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26663;
    wire N__26660;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26630;
    wire N__26627;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26615;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26603;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26591;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26572;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26524;
    wire N__26523;
    wire N__26522;
    wire N__26521;
    wire N__26520;
    wire N__26519;
    wire N__26516;
    wire N__26515;
    wire N__26514;
    wire N__26513;
    wire N__26510;
    wire N__26503;
    wire N__26500;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26493;
    wire N__26490;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26447;
    wire N__26446;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25762;
    wire N__25761;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25739;
    wire N__25736;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25687;
    wire N__25684;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25667;
    wire N__25664;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25653;
    wire N__25650;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25621;
    wire N__25618;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25601;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25540;
    wire N__25537;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25520;
    wire N__25519;
    wire N__25516;
    wire N__25515;
    wire N__25510;
    wire N__25507;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25485;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25460;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25438;
    wire N__25435;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25418;
    wire N__25415;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25403;
    wire N__25400;
    wire N__25399;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25344;
    wire N__25341;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25300;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25246;
    wire N__25245;
    wire N__25244;
    wire N__25241;
    wire N__25236;
    wire N__25233;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25183;
    wire N__25182;
    wire N__25179;
    wire N__25174;
    wire N__25169;
    wire N__25168;
    wire N__25167;
    wire N__25166;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25145;
    wire N__25144;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25120;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25108;
    wire N__25103;
    wire N__25102;
    wire N__25099;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25084;
    wire N__25081;
    wire N__25076;
    wire N__25073;
    wire N__25072;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25049;
    wire N__25046;
    wire N__25045;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25030;
    wire N__25025;
    wire N__25022;
    wire N__25021;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24979;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24956;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24919;
    wire N__24916;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24856;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24798;
    wire N__24795;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24753;
    wire N__24750;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24705;
    wire N__24700;
    wire N__24697;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24676;
    wire N__24671;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24659;
    wire N__24658;
    wire N__24655;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24634;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24602;
    wire N__24601;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24494;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24462;
    wire N__24457;
    wire N__24454;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24436;
    wire N__24435;
    wire N__24434;
    wire N__24433;
    wire N__24432;
    wire N__24431;
    wire N__24428;
    wire N__24427;
    wire N__24426;
    wire N__24423;
    wire N__24422;
    wire N__24419;
    wire N__24418;
    wire N__24417;
    wire N__24412;
    wire N__24409;
    wire N__24408;
    wire N__24401;
    wire N__24398;
    wire N__24393;
    wire N__24386;
    wire N__24383;
    wire N__24378;
    wire N__24373;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24331;
    wire N__24328;
    wire N__24325;
    wire N__24320;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24287;
    wire N__24286;
    wire N__24283;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24262;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24250;
    wire N__24247;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24235;
    wire N__24232;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24197;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24189;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24167;
    wire N__24164;
    wire N__24163;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24130;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24094;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24061;
    wire N__24058;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24043;
    wire N__24040;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24019;
    wire N__24018;
    wire N__24015;
    wire N__24010;
    wire N__24007;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23940;
    wire N__23935;
    wire N__23932;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23907;
    wire N__23902;
    wire N__23899;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23832;
    wire N__23829;
    wire N__23826;
    wire N__23823;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23809;
    wire N__23806;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23782;
    wire N__23779;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23752;
    wire N__23749;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23605;
    wire N__23604;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23596;
    wire N__23593;
    wire N__23592;
    wire N__23589;
    wire N__23588;
    wire N__23585;
    wire N__23580;
    wire N__23571;
    wire N__23564;
    wire N__23561;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23540;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23494;
    wire N__23493;
    wire N__23492;
    wire N__23491;
    wire N__23490;
    wire N__23487;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23479;
    wire N__23476;
    wire N__23475;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23467;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23452;
    wire N__23437;
    wire N__23426;
    wire N__23423;
    wire N__23422;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23396;
    wire N__23393;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23365;
    wire N__23364;
    wire N__23363;
    wire N__23360;
    wire N__23359;
    wire N__23358;
    wire N__23357;
    wire N__23354;
    wire N__23345;
    wire N__23342;
    wire N__23341;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23324;
    wire N__23315;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23284;
    wire N__23281;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23257;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23231;
    wire N__23230;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23156;
    wire N__23155;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23147;
    wire N__23146;
    wire N__23145;
    wire N__23144;
    wire N__23141;
    wire N__23140;
    wire N__23139;
    wire N__23138;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23121;
    wire N__23116;
    wire N__23109;
    wire N__23106;
    wire N__23093;
    wire N__23090;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23050;
    wire N__23049;
    wire N__23046;
    wire N__23041;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23026;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23003;
    wire N__23002;
    wire N__22999;
    wire N__22998;
    wire N__22995;
    wire N__22990;
    wire N__22987;
    wire N__22982;
    wire N__22979;
    wire N__22978;
    wire N__22977;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22943;
    wire N__22942;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22916;
    wire N__22913;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22882;
    wire N__22879;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22820;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22777;
    wire N__22774;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22726;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22659;
    wire N__22654;
    wire N__22651;
    wire N__22646;
    wire N__22643;
    wire N__22642;
    wire N__22639;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22591;
    wire N__22590;
    wire N__22589;
    wire N__22588;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22580;
    wire N__22577;
    wire N__22576;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22568;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22561;
    wire N__22556;
    wire N__22551;
    wire N__22540;
    wire N__22535;
    wire N__22532;
    wire N__22527;
    wire N__22524;
    wire N__22511;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22500;
    wire N__22495;
    wire N__22492;
    wire N__22487;
    wire N__22486;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22471;
    wire N__22466;
    wire N__22465;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22441;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22415;
    wire N__22412;
    wire N__22411;
    wire N__22408;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22378;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22343;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22313;
    wire N__22310;
    wire N__22309;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22213;
    wire N__22210;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22195;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22156;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22139;
    wire N__22138;
    wire N__22135;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22011;
    wire N__22006;
    wire N__22003;
    wire N__21998;
    wire N__21997;
    wire N__21994;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21982;
    wire N__21979;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21955;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21925;
    wire N__21922;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21880;
    wire N__21877;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21821;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21740;
    wire N__21739;
    wire N__21738;
    wire N__21737;
    wire N__21736;
    wire N__21735;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21723;
    wire N__21722;
    wire N__21721;
    wire N__21718;
    wire N__21713;
    wire N__21710;
    wire N__21703;
    wire N__21696;
    wire N__21693;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21640;
    wire N__21637;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21617;
    wire N__21616;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21489;
    wire N__21484;
    wire N__21481;
    wire N__21476;
    wire N__21475;
    wire N__21474;
    wire N__21473;
    wire N__21472;
    wire N__21471;
    wire N__21470;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21444;
    wire N__21443;
    wire N__21434;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21414;
    wire N__21409;
    wire N__21404;
    wire N__21401;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21364;
    wire N__21361;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21340;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21324;
    wire N__21319;
    wire N__21316;
    wire N__21311;
    wire N__21310;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21275;
    wire N__21274;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21239;
    wire N__21236;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21224;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21177;
    wire N__21172;
    wire N__21169;
    wire N__21164;
    wire N__21163;
    wire N__21160;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21110;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21077;
    wire N__21074;
    wire N__21073;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21052;
    wire N__21047;
    wire N__21044;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21032;
    wire N__21029;
    wire N__21028;
    wire N__21025;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20986;
    wire N__20983;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20963;
    wire N__20960;
    wire N__20959;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20935;
    wire N__20930;
    wire N__20927;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20900;
    wire N__20897;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20889;
    wire N__20884;
    wire N__20881;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20802;
    wire N__20797;
    wire N__20794;
    wire N__20789;
    wire N__20786;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20762;
    wire N__20759;
    wire N__20758;
    wire N__20757;
    wire N__20756;
    wire N__20755;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20731;
    wire N__20722;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20710;
    wire N__20709;
    wire N__20706;
    wire N__20701;
    wire N__20696;
    wire N__20693;
    wire N__20692;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20608;
    wire N__20607;
    wire N__20604;
    wire N__20599;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20581;
    wire N__20578;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20536;
    wire N__20535;
    wire N__20532;
    wire N__20527;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20455;
    wire N__20454;
    wire N__20451;
    wire N__20446;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20421;
    wire N__20416;
    wire N__20413;
    wire N__20408;
    wire N__20405;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20393;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20371;
    wire N__20370;
    wire N__20369;
    wire N__20368;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20344;
    wire N__20339;
    wire N__20334;
    wire N__20327;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20321;
    wire N__20320;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20296;
    wire N__20287;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20272;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20230;
    wire N__20227;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20185;
    wire N__20184;
    wire N__20181;
    wire N__20176;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20147;
    wire N__20146;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20129;
    wire N__20128;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20108;
    wire N__20107;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20090;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20071;
    wire N__20068;
    wire N__20063;
    wire N__20062;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20042;
    wire N__20041;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19951;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19771;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19741;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19681;
    wire N__19680;
    wire N__19679;
    wire N__19678;
    wire N__19675;
    wire N__19674;
    wire N__19673;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19667;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19656;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19644;
    wire N__19643;
    wire N__19642;
    wire N__19639;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19621;
    wire N__19618;
    wire N__19609;
    wire N__19602;
    wire N__19589;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19448;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19434;
    wire N__19429;
    wire N__19426;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19318;
    wire N__19317;
    wire N__19314;
    wire N__19309;
    wire N__19306;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19258;
    wire N__19255;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19222;
    wire N__19221;
    wire N__19220;
    wire N__19219;
    wire N__19216;
    wire N__19215;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19207;
    wire N__19206;
    wire N__19205;
    wire N__19204;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19196;
    wire N__19195;
    wire N__19194;
    wire N__19191;
    wire N__19190;
    wire N__19189;
    wire N__19188;
    wire N__19185;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19173;
    wire N__19172;
    wire N__19169;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19161;
    wire N__19158;
    wire N__19151;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19133;
    wire N__19126;
    wire N__19115;
    wire N__19108;
    wire N__19101;
    wire N__19088;
    wire N__19085;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18925;
    wire N__18920;
    wire N__18917;
    wire N__18916;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18849;
    wire N__18844;
    wire N__18841;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18784;
    wire N__18783;
    wire N__18780;
    wire N__18779;
    wire N__18778;
    wire N__18777;
    wire N__18776;
    wire N__18775;
    wire N__18774;
    wire N__18771;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18746;
    wire N__18745;
    wire N__18742;
    wire N__18741;
    wire N__18740;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18723;
    wire N__18714;
    wire N__18707;
    wire N__18700;
    wire N__18693;
    wire N__18688;
    wire N__18677;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18565;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18460;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18445;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18427;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18364;
    wire N__18363;
    wire N__18360;
    wire N__18355;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18331;
    wire N__18328;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18197;
    wire N__18194;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18172;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18145;
    wire N__18144;
    wire N__18143;
    wire N__18142;
    wire N__18139;
    wire N__18138;
    wire N__18135;
    wire N__18134;
    wire N__18133;
    wire N__18130;
    wire N__18129;
    wire N__18128;
    wire N__18125;
    wire N__18124;
    wire N__18121;
    wire N__18120;
    wire N__18119;
    wire N__18116;
    wire N__18111;
    wire N__18110;
    wire N__18109;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18101;
    wire N__18100;
    wire N__18097;
    wire N__18092;
    wire N__18089;
    wire N__18080;
    wire N__18075;
    wire N__18068;
    wire N__18059;
    wire N__18056;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18034;
    wire N__18033;
    wire N__18030;
    wire N__18025;
    wire N__18022;
    wire N__18017;
    wire N__18014;
    wire N__18013;
    wire N__18010;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17995;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17983;
    wire N__17980;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17957;
    wire N__17956;
    wire N__17955;
    wire N__17954;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17948;
    wire N__17947;
    wire N__17946;
    wire N__17945;
    wire N__17942;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17934;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17926;
    wire N__17923;
    wire N__17922;
    wire N__17921;
    wire N__17920;
    wire N__17919;
    wire N__17916;
    wire N__17915;
    wire N__17912;
    wire N__17907;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17868;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17836;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17821;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17782;
    wire N__17779;
    wire N__17778;
    wire N__17777;
    wire N__17776;
    wire N__17775;
    wire N__17774;
    wire N__17773;
    wire N__17772;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17764;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17758;
    wire N__17755;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17745;
    wire N__17744;
    wire N__17741;
    wire N__17740;
    wire N__17737;
    wire N__17736;
    wire N__17735;
    wire N__17732;
    wire N__17731;
    wire N__17726;
    wire N__17721;
    wire N__17716;
    wire N__17709;
    wire N__17700;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17682;
    wire N__17679;
    wire N__17660;
    wire N__17659;
    wire N__17656;
    wire N__17655;
    wire N__17652;
    wire N__17649;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17630;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17513;
    wire N__17510;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17495;
    wire N__17492;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17388;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17320;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17300;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17274;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17217;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17159;
    wire N__17158;
    wire N__17157;
    wire N__17156;
    wire N__17155;
    wire N__17152;
    wire N__17151;
    wire N__17150;
    wire N__17149;
    wire N__17148;
    wire N__17147;
    wire N__17146;
    wire N__17145;
    wire N__17142;
    wire N__17141;
    wire N__17140;
    wire N__17137;
    wire N__17136;
    wire N__17133;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17125;
    wire N__17124;
    wire N__17123;
    wire N__17120;
    wire N__17119;
    wire N__17116;
    wire N__17115;
    wire N__17112;
    wire N__17107;
    wire N__17096;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17074;
    wire N__17065;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17022;
    wire N__17019;
    wire N__17014;
    wire N__17011;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16990;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16974;
    wire N__16971;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16906;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16885;
    wire N__16880;
    wire N__16879;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16840;
    wire N__16837;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16820;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16793;
    wire N__16790;
    wire N__16789;
    wire N__16786;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16767;
    wire N__16764;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16738;
    wire N__16737;
    wire N__16734;
    wire N__16731;
    wire N__16728;
    wire N__16725;
    wire N__16718;
    wire N__16715;
    wire N__16714;
    wire N__16711;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16657;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16618;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16582;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16486;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16453;
    wire N__16450;
    wire N__16449;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16330;
    wire N__16329;
    wire N__16328;
    wire N__16325;
    wire N__16324;
    wire N__16323;
    wire N__16322;
    wire N__16321;
    wire N__16320;
    wire N__16319;
    wire N__16314;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16301;
    wire N__16300;
    wire N__16299;
    wire N__16298;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16290;
    wire N__16289;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16280;
    wire N__16279;
    wire N__16278;
    wire N__16277;
    wire N__16274;
    wire N__16269;
    wire N__16260;
    wire N__16247;
    wire N__16236;
    wire N__16227;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16141;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16129;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16105;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16063;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15993;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15961;
    wire N__15960;
    wire N__15957;
    wire N__15952;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15916;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15906;
    wire N__15901;
    wire N__15898;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15870;
    wire N__15867;
    wire N__15864;
    wire N__15861;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15832;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15691;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15655;
    wire N__15654;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15499;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15469;
    wire N__15466;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15295;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15271;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15226;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15211;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15184;
    wire N__15183;
    wire N__15180;
    wire N__15175;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15086;
    wire N__15083;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14998;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14980;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14914;
    wire N__14911;
    wire N__14910;
    wire N__14907;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14875;
    wire N__14874;
    wire N__14871;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14842;
    wire N__14841;
    wire N__14836;
    wire N__14833;
    wire N__14828;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14763;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14644;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14626;
    wire N__14621;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14581;
    wire N__14580;
    wire N__14577;
    wire N__14572;
    wire N__14569;
    wire N__14564;
    wire N__14561;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14512;
    wire N__14509;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14499;
    wire N__14492;
    wire N__14491;
    wire N__14488;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14478;
    wire N__14475;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14442;
    wire N__14439;
    wire N__14436;
    wire N__14433;
    wire N__14426;
    wire N__14423;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14359;
    wire N__14358;
    wire N__14355;
    wire N__14350;
    wire N__14347;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14304;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14288;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14260;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14245;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14195;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14187;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14157;
    wire N__14154;
    wire N__14151;
    wire N__14148;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14057;
    wire N__14056;
    wire N__14053;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14036;
    wire N__14035;
    wire N__14032;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14002;
    wire N__14001;
    wire N__13998;
    wire N__13993;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13952;
    wire N__13951;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13925;
    wire N__13924;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13911;
    wire N__13908;
    wire N__13905;
    wire N__13898;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13890;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13876;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13819;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13799;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13784;
    wire N__13781;
    wire N__13780;
    wire N__13779;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13760;
    wire N__13759;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13579;
    wire N__13576;
    wire N__13573;
    wire N__13568;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13558;
    wire N__13557;
    wire N__13552;
    wire N__13549;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13510;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13491;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13450;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13436;
    wire N__13435;
    wire N__13434;
    wire N__13431;
    wire N__13430;
    wire N__13429;
    wire N__13428;
    wire N__13427;
    wire N__13426;
    wire N__13421;
    wire N__13416;
    wire N__13407;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13378;
    wire N__13375;
    wire N__13372;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13246;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13231;
    wire N__13226;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13048;
    wire N__13045;
    wire N__13042;
    wire N__13039;
    wire N__13036;
    wire N__13035;
    wire N__13030;
    wire N__13027;
    wire N__13022;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12977;
    wire N__12974;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12862;
    wire N__12859;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12796;
    wire N__12793;
    wire N__12790;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12757;
    wire N__12754;
    wire N__12751;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12706;
    wire N__12705;
    wire N__12702;
    wire N__12697;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12463;
    wire N__12458;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12446;
    wire N__12445;
    wire N__12444;
    wire N__12439;
    wire N__12436;
    wire N__12431;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12423;
    wire N__12418;
    wire N__12415;
    wire N__12410;
    wire N__12409;
    wire N__12408;
    wire N__12403;
    wire N__12400;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12353;
    wire N__12352;
    wire N__12349;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12332;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire LED_c;
    wire n26;
    wire bfn_17_17_0_;
    wire n25;
    wire n3906;
    wire n24;
    wire n3907;
    wire n23;
    wire n3908;
    wire n22;
    wire n3909;
    wire n21;
    wire n3910;
    wire n20;
    wire n3911;
    wire n19;
    wire n3912;
    wire n3913;
    wire n18;
    wire bfn_17_18_0_;
    wire n17;
    wire n3914;
    wire n16;
    wire n3915;
    wire n15;
    wire n3916;
    wire n14;
    wire n3917;
    wire n13;
    wire n3918;
    wire n12;
    wire n3919;
    wire n11_adj_364;
    wire n3920;
    wire n3921;
    wire n10_adj_363;
    wire bfn_17_19_0_;
    wire n9;
    wire n3922;
    wire n8_adj_362;
    wire n3923;
    wire n7;
    wire n3924;
    wire n6;
    wire n3925;
    wire n3926;
    wire n3927;
    wire n3928;
    wire n3929;
    wire bfn_17_20_0_;
    wire n3930;
    wire blink_counter_25;
    wire bfn_17_21_0_;
    wire \eeprom.n4183 ;
    wire \eeprom.n4184 ;
    wire \eeprom.n4185 ;
    wire \eeprom.n4186 ;
    wire \eeprom.n4187 ;
    wire \eeprom.n4188 ;
    wire \eeprom.n4189 ;
    wire \eeprom.n4190 ;
    wire bfn_17_22_0_;
    wire \eeprom.n4191 ;
    wire \eeprom.n4192 ;
    wire \eeprom.n4193 ;
    wire \eeprom.n4194 ;
    wire \eeprom.n4195 ;
    wire \eeprom.n4196 ;
    wire \eeprom.n4197 ;
    wire \eeprom.n4198 ;
    wire bfn_17_23_0_;
    wire \eeprom.n4199 ;
    wire \eeprom.n4200 ;
    wire \eeprom.n4201 ;
    wire \eeprom.n4202 ;
    wire \eeprom.n4203 ;
    wire \eeprom.n4204 ;
    wire bfn_17_24_0_;
    wire \eeprom.n4162 ;
    wire \eeprom.n4163 ;
    wire \eeprom.n4164 ;
    wire \eeprom.n4165 ;
    wire \eeprom.n4166 ;
    wire \eeprom.n4167 ;
    wire \eeprom.n4168 ;
    wire \eeprom.n4169 ;
    wire bfn_17_25_0_;
    wire \eeprom.n4170 ;
    wire \eeprom.n4171 ;
    wire \eeprom.n4172 ;
    wire \eeprom.n4173 ;
    wire \eeprom.n4174 ;
    wire \eeprom.n3372 ;
    wire \eeprom.n4175 ;
    wire \eeprom.n4176 ;
    wire \eeprom.n4177 ;
    wire bfn_17_26_0_;
    wire \eeprom.n4178 ;
    wire \eeprom.n4179 ;
    wire \eeprom.n4180 ;
    wire \eeprom.n4181 ;
    wire \eeprom.n4182 ;
    wire bfn_17_27_0_;
    wire \eeprom.n4142 ;
    wire \eeprom.n4143 ;
    wire \eeprom.n4144 ;
    wire \eeprom.n4145 ;
    wire \eeprom.n4146 ;
    wire \eeprom.n4147 ;
    wire \eeprom.n4148 ;
    wire \eeprom.n4149 ;
    wire bfn_17_28_0_;
    wire \eeprom.n3277 ;
    wire \eeprom.n4150 ;
    wire \eeprom.n4151 ;
    wire \eeprom.n4152 ;
    wire \eeprom.n4153 ;
    wire \eeprom.n4154 ;
    wire \eeprom.n4155 ;
    wire \eeprom.n4156 ;
    wire \eeprom.n4157 ;
    wire bfn_17_29_0_;
    wire \eeprom.n4158 ;
    wire \eeprom.n4159 ;
    wire \eeprom.n4160 ;
    wire \eeprom.n4161 ;
    wire bfn_18_17_0_;
    wire \eeprom.n3966 ;
    wire \eeprom.n3967 ;
    wire \eeprom.n3968 ;
    wire \eeprom.n3969 ;
    wire \eeprom.n3970 ;
    wire \eeprom.n3971 ;
    wire \eeprom.n3972 ;
    wire n5421;
    wire blink_counter_24;
    wire blink_counter_22;
    wire blink_counter_23;
    wire blink_counter_21;
    wire n5420;
    wire \eeprom.n1203 ;
    wire \eeprom.n3713_cascade_ ;
    wire \eeprom.n3618_cascade_ ;
    wire \eeprom.n3615_cascade_ ;
    wire \eeprom.n5221_cascade_ ;
    wire \eeprom.n5225 ;
    wire \eeprom.n3614 ;
    wire \eeprom.n3605 ;
    wire \eeprom.n3471 ;
    wire \eeprom.n32_cascade_ ;
    wire \eeprom.n3529_cascade_ ;
    wire \eeprom.n3481 ;
    wire \eeprom.n3513_cascade_ ;
    wire \eeprom.n3473 ;
    wire \eeprom.n3505_cascade_ ;
    wire \eeprom.n30_adj_273 ;
    wire \eeprom.n3478 ;
    wire \eeprom.n3472 ;
    wire \eeprom.n3484 ;
    wire \eeprom.n3475 ;
    wire \eeprom.n3507_cascade_ ;
    wire \eeprom.n31 ;
    wire \eeprom.n3482 ;
    wire \eeprom.n3514_cascade_ ;
    wire \eeprom.n5323_cascade_ ;
    wire \eeprom.n5321 ;
    wire \eeprom.n4753 ;
    wire \eeprom.n3376 ;
    wire \eeprom.n3380 ;
    wire \eeprom.n3412 ;
    wire \eeprom.n3412_cascade_ ;
    wire \eeprom.n3479 ;
    wire \eeprom.n3375 ;
    wire \eeprom.n3378 ;
    wire \eeprom.n3410 ;
    wire \eeprom.n3477 ;
    wire \eeprom.n3410_cascade_ ;
    wire \eeprom.n3465 ;
    wire \eeprom.n3367 ;
    wire \eeprom.n3267 ;
    wire \eeprom.n3299_cascade_ ;
    wire \eeprom.n3298 ;
    wire \eeprom.n3379 ;
    wire \eeprom.n3299 ;
    wire \eeprom.n3366 ;
    wire \eeprom.n3269 ;
    wire \eeprom.n3301 ;
    wire \eeprom.n3301_cascade_ ;
    wire \eeprom.n3368 ;
    wire \eeprom.n3374 ;
    wire \eeprom.n3406 ;
    wire \eeprom.n3370 ;
    wire \eeprom.n3268 ;
    wire \eeprom.n3300 ;
    wire \eeprom.n3200 ;
    wire \eeprom.n3200_cascade_ ;
    wire \eeprom.n3286 ;
    wire \eeprom.n3280 ;
    wire \eeprom.n3275 ;
    wire \eeprom.n3276 ;
    wire \eeprom.n3279 ;
    wire \eeprom.n3204_cascade_ ;
    wire \eeprom.n3273 ;
    wire \eeprom.n3206_cascade_ ;
    wire \eeprom.n3108_cascade_ ;
    wire \eeprom.n3202 ;
    wire \eeprom.n3201 ;
    wire \eeprom.n3203 ;
    wire \eeprom.n3270 ;
    wire \eeprom.n3203_cascade_ ;
    wire \eeprom.n3113_cascade_ ;
    wire \eeprom.n5305_cascade_ ;
    wire \eeprom.n3034_cascade_ ;
    wire bfn_18_29_0_;
    wire \eeprom.n3085 ;
    wire \eeprom.n4105 ;
    wire \eeprom.n3084 ;
    wire \eeprom.n4106 ;
    wire \eeprom.n3083 ;
    wire \eeprom.n4107 ;
    wire \eeprom.n4108 ;
    wire \eeprom.n3081 ;
    wire \eeprom.n4109 ;
    wire \eeprom.n4110 ;
    wire \eeprom.n3079 ;
    wire \eeprom.n4111 ;
    wire \eeprom.n4112 ;
    wire bfn_18_30_0_;
    wire \eeprom.n3077 ;
    wire \eeprom.n4113 ;
    wire \eeprom.n3076 ;
    wire \eeprom.n4114 ;
    wire \eeprom.n3075 ;
    wire \eeprom.n4115 ;
    wire \eeprom.n4116 ;
    wire \eeprom.n4117 ;
    wire \eeprom.n4118 ;
    wire \eeprom.n4119 ;
    wire \eeprom.n4120 ;
    wire \eeprom.n3070 ;
    wire bfn_18_31_0_;
    wire \eeprom.n3069 ;
    wire \eeprom.n4121 ;
    wire \eeprom.n4122 ;
    wire \eeprom.n3071 ;
    wire \eeprom.n3004 ;
    wire \eeprom.n3613 ;
    wire \eeprom.n1202 ;
    wire \eeprom.n3712_cascade_ ;
    wire \eeprom.n1207 ;
    wire \eeprom.n3618 ;
    wire \eeprom.n3717_cascade_ ;
    wire \eeprom.n1208 ;
    wire \eeprom.n5362_cascade_ ;
    wire \eeprom.n1206 ;
    wire \eeprom.n1205 ;
    wire \eeprom.n3616 ;
    wire \eeprom.n3715_cascade_ ;
    wire \eeprom.n5017 ;
    wire \eeprom.n5019_cascade_ ;
    wire \eeprom.n28_adj_342_cascade_ ;
    wire \eeprom.n3615 ;
    wire \eeprom.n3628_cascade_ ;
    wire \eeprom.n1204 ;
    wire \eeprom.n3714_cascade_ ;
    wire \eeprom.n1201 ;
    wire \eeprom.n3628 ;
    wire \eeprom.n5025_cascade_ ;
    wire \eeprom.n5027_cascade_ ;
    wire \eeprom.n5029_cascade_ ;
    wire \eeprom.n5031_cascade_ ;
    wire \eeprom.n5161 ;
    wire \eeprom.n29_adj_274 ;
    wire \eeprom.n3612 ;
    wire \eeprom.n3617 ;
    wire \eeprom.n3596 ;
    wire \eeprom.n3609_cascade_ ;
    wire \eeprom.n5021_cascade_ ;
    wire \eeprom.n5023 ;
    wire \eeprom.n3474 ;
    wire \eeprom.n3407 ;
    wire \eeprom.n3486 ;
    wire \eeprom.n3468 ;
    wire \eeprom.n3608_cascade_ ;
    wire \eeprom.n3480 ;
    wire \eeprom.n3512_cascade_ ;
    wire \eeprom.n5175 ;
    wire \eeprom.n5177_cascade_ ;
    wire \eeprom.n31_adj_341 ;
    wire \eeprom.n3598 ;
    wire \eeprom.n3483 ;
    wire \eeprom.n3485 ;
    wire \eeprom.n3398 ;
    wire \eeprom.n3397 ;
    wire \eeprom.n3408 ;
    wire \eeprom.n3411 ;
    wire \eeprom.n18_cascade_ ;
    wire \eeprom.n29 ;
    wire \eeprom.n30_cascade_ ;
    wire \eeprom.n3430_cascade_ ;
    wire \eeprom.n3467 ;
    wire \eeprom.n3466 ;
    wire \eeprom.n3498_cascade_ ;
    wire \eeprom.n28_adj_267 ;
    wire \eeprom.n3476 ;
    wire \eeprom.n3373 ;
    wire \eeprom.n3369 ;
    wire \eeprom.n3401 ;
    wire \eeprom.n3400 ;
    wire \eeprom.n3399 ;
    wire \eeprom.n3401_cascade_ ;
    wire \eeprom.n27_adj_263 ;
    wire \eeprom.n3402 ;
    wire \eeprom.n3469 ;
    wire \eeprom.n3307 ;
    wire \eeprom.n3311 ;
    wire \eeprom.n3312 ;
    wire \eeprom.n3309 ;
    wire \eeprom.n28_cascade_ ;
    wire \eeprom.n25 ;
    wire \eeprom.n3385 ;
    wire \eeprom.n3331_cascade_ ;
    wire \eeprom.n3281 ;
    wire \eeprom.n3206 ;
    wire \eeprom.n20_adj_301_cascade_ ;
    wire \eeprom.n16_adj_303 ;
    wire \eeprom.n3212 ;
    wire \eeprom.n28_adj_305_cascade_ ;
    wire \eeprom.n24_adj_304 ;
    wire \eeprom.n3232_cascade_ ;
    wire \eeprom.n3274 ;
    wire \eeprom.n3306 ;
    wire \eeprom.n3305 ;
    wire \eeprom.n3306_cascade_ ;
    wire \eeprom.n3308 ;
    wire \eeprom.n27 ;
    wire \eeprom.n5309 ;
    wire \eeprom.n18_adj_260_cascade_ ;
    wire \eeprom.n24 ;
    wire \eeprom.n22 ;
    wire \eeprom.n26_adj_262_cascade_ ;
    wire \eeprom.n3133_cascade_ ;
    wire \eeprom.n3205 ;
    wire \eeprom.n3272 ;
    wire \eeprom.n3205_cascade_ ;
    wire \eeprom.n3204 ;
    wire \eeprom.n3271 ;
    wire \eeprom.n3207 ;
    wire \eeprom.n3017 ;
    wire \eeprom.n3017_cascade_ ;
    wire \eeprom.n5147_cascade_ ;
    wire \eeprom.n3009 ;
    wire \eeprom.n3002 ;
    wire \eeprom.n3002_cascade_ ;
    wire \eeprom.n20_adj_337 ;
    wire \eeprom.n3078 ;
    wire \eeprom.n3016 ;
    wire \eeprom.n3018 ;
    wire \eeprom.n2914_cascade_ ;
    wire \eeprom.n3073 ;
    wire \eeprom.n3014 ;
    wire \eeprom.n3007 ;
    wire \eeprom.n3074 ;
    wire \eeprom.n3007_cascade_ ;
    wire \eeprom.n3006 ;
    wire \eeprom.n21_adj_336 ;
    wire \eeprom.n3006_cascade_ ;
    wire \eeprom.n18_adj_335 ;
    wire \eeprom.n24_adj_340 ;
    wire \eeprom.n3008 ;
    wire \eeprom.n3005 ;
    wire \eeprom.n3005_cascade_ ;
    wire \eeprom.n3072 ;
    wire \eeprom.n3082 ;
    wire \eeprom.n3010 ;
    wire \eeprom.n3012 ;
    wire \eeprom.n3003 ;
    wire \eeprom.n3086 ;
    wire \eeprom.n3186 ;
    wire bfn_19_30_0_;
    wire \eeprom.n4123 ;
    wire \eeprom.n3117 ;
    wire \eeprom.n3184 ;
    wire \eeprom.n4124 ;
    wire \eeprom.n4125 ;
    wire \eeprom.n4126 ;
    wire \eeprom.n4127 ;
    wire \eeprom.n3113 ;
    wire \eeprom.n3180 ;
    wire \eeprom.n4128 ;
    wire \eeprom.n3179 ;
    wire \eeprom.n4129 ;
    wire \eeprom.n4130 ;
    wire \eeprom.n3111 ;
    wire \eeprom.n3178 ;
    wire bfn_19_31_0_;
    wire \eeprom.n4131 ;
    wire \eeprom.n4132 ;
    wire \eeprom.n3108 ;
    wire \eeprom.n3175 ;
    wire \eeprom.n4133 ;
    wire \eeprom.n3107 ;
    wire \eeprom.n3174 ;
    wire \eeprom.n4134 ;
    wire \eeprom.n3106 ;
    wire \eeprom.n3173 ;
    wire \eeprom.n4135 ;
    wire \eeprom.n3105 ;
    wire \eeprom.n3172 ;
    wire \eeprom.n4136 ;
    wire \eeprom.n3104 ;
    wire \eeprom.n3171 ;
    wire \eeprom.n4137 ;
    wire \eeprom.n4138 ;
    wire \eeprom.n3103 ;
    wire \eeprom.n3170 ;
    wire bfn_19_32_0_;
    wire \eeprom.n3102 ;
    wire \eeprom.n3169 ;
    wire \eeprom.n4139 ;
    wire \eeprom.n3101 ;
    wire \eeprom.n3168 ;
    wire \eeprom.n4140 ;
    wire \eeprom.n3100 ;
    wire \eeprom.n4141 ;
    wire \eeprom.n3199 ;
    wire bfn_20_17_0_;
    wire \eeprom.n4228 ;
    wire \eeprom.n4229 ;
    wire \eeprom.n4230 ;
    wire \eeprom.n4231 ;
    wire \eeprom.n4232 ;
    wire \eeprom.n4233 ;
    wire \eeprom.n5547 ;
    wire \eeprom.n5362 ;
    wire \eeprom.n4234 ;
    wire \eeprom.n4235 ;
    wire \eeprom.n5550 ;
    wire \eeprom.n3717 ;
    wire bfn_20_18_0_;
    wire \eeprom.n4236 ;
    wire \eeprom.n5556 ;
    wire \eeprom.n3715 ;
    wire \eeprom.n4237 ;
    wire \eeprom.n5559 ;
    wire \eeprom.n3714 ;
    wire \eeprom.n4238 ;
    wire \eeprom.n5562 ;
    wire \eeprom.n3713 ;
    wire \eeprom.n4239 ;
    wire \eeprom.n5565 ;
    wire \eeprom.n3712 ;
    wire \eeprom.n4240 ;
    wire \eeprom.n3711 ;
    wire \eeprom.n5568 ;
    wire \eeprom.n4241 ;
    wire \eeprom.n3716 ;
    wire \eeprom.n5553 ;
    wire \eeprom.n3586 ;
    wire bfn_20_19_0_;
    wire \eeprom.n3518 ;
    wire \eeprom.n3585_adj_296 ;
    wire \eeprom.n4205 ;
    wire \eeprom.n3517 ;
    wire \eeprom.n3584 ;
    wire \eeprom.n4206 ;
    wire \eeprom.n3516 ;
    wire \eeprom.n3583 ;
    wire \eeprom.n4207 ;
    wire \eeprom.n3515 ;
    wire \eeprom.n3582 ;
    wire \eeprom.n4208 ;
    wire \eeprom.n3514 ;
    wire \eeprom.n3581_adj_292 ;
    wire \eeprom.n4209 ;
    wire \eeprom.n3513 ;
    wire \eeprom.n3580 ;
    wire \eeprom.n4210 ;
    wire \eeprom.n3512 ;
    wire \eeprom.n3579 ;
    wire \eeprom.n4211 ;
    wire \eeprom.n4212 ;
    wire \eeprom.n3511 ;
    wire \eeprom.n3578 ;
    wire bfn_20_20_0_;
    wire \eeprom.n3510 ;
    wire \eeprom.n3577 ;
    wire \eeprom.n4213 ;
    wire \eeprom.n3509 ;
    wire \eeprom.n3576 ;
    wire \eeprom.n4214 ;
    wire \eeprom.n3508 ;
    wire \eeprom.n3575 ;
    wire \eeprom.n4215 ;
    wire \eeprom.n3507 ;
    wire \eeprom.n3574 ;
    wire \eeprom.n4216 ;
    wire \eeprom.n3506 ;
    wire \eeprom.n3573 ;
    wire \eeprom.n4217 ;
    wire \eeprom.n3505 ;
    wire \eeprom.n3572 ;
    wire \eeprom.n4218 ;
    wire \eeprom.n3504 ;
    wire \eeprom.n3571 ;
    wire \eeprom.n4219 ;
    wire \eeprom.n4220 ;
    wire \eeprom.n3503 ;
    wire \eeprom.n3570 ;
    wire bfn_20_21_0_;
    wire \eeprom.n3569 ;
    wire \eeprom.n4221 ;
    wire \eeprom.n3501 ;
    wire \eeprom.n3568 ;
    wire \eeprom.n4222 ;
    wire \eeprom.n3500 ;
    wire \eeprom.n3567 ;
    wire \eeprom.n4223 ;
    wire \eeprom.n3499 ;
    wire \eeprom.n3566 ;
    wire \eeprom.n4224 ;
    wire \eeprom.n3498 ;
    wire \eeprom.n3565 ;
    wire \eeprom.n4225 ;
    wire \eeprom.n3497 ;
    wire \eeprom.n3564 ;
    wire \eeprom.n4226 ;
    wire \eeprom.n3496 ;
    wire \eeprom.n3529 ;
    wire \eeprom.n4227 ;
    wire \eeprom.n5355 ;
    wire \eeprom.n3382 ;
    wire \eeprom.n3414 ;
    wire \eeprom.n3417 ;
    wire \eeprom.n3414_cascade_ ;
    wire \eeprom.n5291_cascade_ ;
    wire \eeprom.n3405 ;
    wire \eeprom.n4824_cascade_ ;
    wire \eeprom.n3404 ;
    wire \eeprom.n28_adj_261 ;
    wire \eeprom.n3386 ;
    wire \eeprom.n3418 ;
    wire \eeprom.n3384 ;
    wire \eeprom.n3416 ;
    wire \eeprom.n3383 ;
    wire \eeprom.n3313 ;
    wire \eeprom.n3371 ;
    wire \eeprom.n3282 ;
    wire \eeprom.n3381 ;
    wire \eeprom.n3314_cascade_ ;
    wire \eeprom.n3413 ;
    wire \eeprom.n3413_cascade_ ;
    wire \eeprom.n3415 ;
    wire \eeprom.n5289 ;
    wire \eeprom.n3278 ;
    wire \eeprom.n3310 ;
    wire \eeprom.n3331 ;
    wire \eeprom.n3310_cascade_ ;
    wire \eeprom.n3377 ;
    wire \eeprom.n3409 ;
    wire \eeprom.n3284 ;
    wire \eeprom.n3218 ;
    wire \eeprom.n3285 ;
    wire \eeprom.n3317 ;
    wire \eeprom.n3314 ;
    wire \eeprom.n3317_cascade_ ;
    wire \eeprom.n3316 ;
    wire \eeprom.n3318 ;
    wire \eeprom.n5315_cascade_ ;
    wire \eeprom.n5313 ;
    wire \eeprom.n3303 ;
    wire \eeprom.n3304 ;
    wire \eeprom.n4820_cascade_ ;
    wire \eeprom.n3302 ;
    wire \eeprom.n26 ;
    wire \eeprom.n3283 ;
    wire \eeprom.n3232 ;
    wire \eeprom.n3315 ;
    wire \eeprom.n3114 ;
    wire \eeprom.n3181 ;
    wire \eeprom.n3213 ;
    wire \eeprom.n3213_cascade_ ;
    wire \eeprom.n3182 ;
    wire \eeprom.n3115 ;
    wire \eeprom.n3214 ;
    wire \eeprom.n3216 ;
    wire \eeprom.n3214_cascade_ ;
    wire \eeprom.n5205 ;
    wire \eeprom.n5209 ;
    wire \eeprom.n3116 ;
    wire \eeprom.n3183 ;
    wire \eeprom.n3215 ;
    wire \eeprom.n3185 ;
    wire \eeprom.n3118 ;
    wire \eeprom.n3217 ;
    wire \eeprom.n3109 ;
    wire \eeprom.n3176 ;
    wire \eeprom.n3208 ;
    wire \eeprom.n3211 ;
    wire \eeprom.n3208_cascade_ ;
    wire \eeprom.n3210 ;
    wire \eeprom.n26_adj_302 ;
    wire \eeprom.n3080 ;
    wire \eeprom.n3013_cascade_ ;
    wire \eeprom.n3034 ;
    wire \eeprom.n3112 ;
    wire \eeprom.n3011 ;
    wire \eeprom.n5301 ;
    wire \eeprom.n3110 ;
    wire \eeprom.n3133 ;
    wire \eeprom.n3177 ;
    wire \eeprom.n3209 ;
    wire \eeprom.n2910_cascade_ ;
    wire \eeprom.n15_adj_300 ;
    wire \eeprom.n22_adj_331_cascade_ ;
    wire \eeprom.n18_adj_330 ;
    wire \eeprom.n2935_cascade_ ;
    wire \eeprom.n3015 ;
    wire \eeprom.n3013 ;
    wire \eeprom.n3015_cascade_ ;
    wire \eeprom.n5143 ;
    wire \eeprom.n18_adj_290_cascade_ ;
    wire \eeprom.n20_adj_291_cascade_ ;
    wire \eeprom.n2836_cascade_ ;
    wire \eeprom.n2913_cascade_ ;
    wire \eeprom.n5297 ;
    wire \eeprom.n2986 ;
    wire bfn_20_29_0_;
    wire \eeprom.n2985 ;
    wire \eeprom.n4088 ;
    wire \eeprom.n2917 ;
    wire \eeprom.n2984 ;
    wire \eeprom.n4089 ;
    wire \eeprom.n2916 ;
    wire \eeprom.n2983 ;
    wire \eeprom.n4090 ;
    wire \eeprom.n2915 ;
    wire \eeprom.n2982 ;
    wire \eeprom.n4091 ;
    wire \eeprom.n2914 ;
    wire \eeprom.n2981 ;
    wire \eeprom.n4092 ;
    wire \eeprom.n2913 ;
    wire \eeprom.n2980 ;
    wire \eeprom.n4093 ;
    wire \eeprom.n2979 ;
    wire \eeprom.n4094 ;
    wire \eeprom.n4095 ;
    wire \eeprom.n2978 ;
    wire bfn_20_30_0_;
    wire \eeprom.n2910 ;
    wire \eeprom.n2977 ;
    wire \eeprom.n4096 ;
    wire \eeprom.n2909 ;
    wire \eeprom.n2976 ;
    wire \eeprom.n4097 ;
    wire \eeprom.n2908 ;
    wire \eeprom.n2975 ;
    wire \eeprom.n4098 ;
    wire \eeprom.n2974 ;
    wire \eeprom.n4099 ;
    wire \eeprom.n2906 ;
    wire \eeprom.n2973 ;
    wire \eeprom.n4100 ;
    wire \eeprom.n2972 ;
    wire \eeprom.n4101 ;
    wire \eeprom.n2971 ;
    wire \eeprom.n4102 ;
    wire \eeprom.n4103 ;
    wire \eeprom.n2970 ;
    wire bfn_20_31_0_;
    wire \eeprom.n2935 ;
    wire \eeprom.n4104 ;
    wire \eeprom.n3001 ;
    wire \eeprom.enable_N_60_0 ;
    wire \eeprom.enable_N_60_1 ;
    wire \eeprom.enable_N_60_2 ;
    wire \eeprom.enable_N_60_3 ;
    wire \eeprom.enable_N_60_4 ;
    wire \eeprom.n4847_cascade_ ;
    wire \eeprom.enable_N_60_5 ;
    wire \eeprom.enable_N_60_7 ;
    wire \eeprom.enable_N_60_6 ;
    wire \eeprom.n4853_cascade_ ;
    wire \eeprom.enable_N_60_8 ;
    wire \eeprom.enable_N_60_10 ;
    wire \eeprom.enable_N_60_9 ;
    wire \eeprom.n4859_cascade_ ;
    wire \eeprom.enable_N_60_11 ;
    wire \eeprom.n4865_cascade_ ;
    wire \eeprom.enable_N_59_cascade_ ;
    wire \eeprom.enable_N_60_12 ;
    wire \eeprom.enable_N_60_14 ;
    wire \eeprom.enable_N_60_13 ;
    wire \eeprom.n4865 ;
    wire \eeprom.n2211_cascade_ ;
    wire \eeprom.n2214_cascade_ ;
    wire \eeprom.n3720 ;
    wire bfn_21_20_0_;
    wire \eeprom.n4007 ;
    wire \eeprom.n4008 ;
    wire \eeprom.n4009 ;
    wire \eeprom.n4010 ;
    wire \eeprom.n4011 ;
    wire \eeprom.n4012 ;
    wire \eeprom.n4013 ;
    wire \eeprom.n4014 ;
    wire bfn_21_21_0_;
    wire \eeprom.n4015 ;
    wire \eeprom.n4016 ;
    wire \eeprom.n4017 ;
    wire \eeprom.n3403 ;
    wire \eeprom.n3470 ;
    wire \eeprom.n3430 ;
    wire \eeprom.n3502 ;
    wire \eeprom.n2511_cascade_ ;
    wire \eeprom.n2618_cascade_ ;
    wire bfn_21_23_0_;
    wire \eeprom.n2685 ;
    wire \eeprom.n4043 ;
    wire \eeprom.n4044 ;
    wire \eeprom.n4045 ;
    wire \eeprom.n4046 ;
    wire \eeprom.n4047 ;
    wire \eeprom.n4048 ;
    wire \eeprom.n4049 ;
    wire \eeprom.n4050 ;
    wire bfn_21_24_0_;
    wire \eeprom.n4051 ;
    wire \eeprom.n4052 ;
    wire \eeprom.n4053 ;
    wire \eeprom.n4054 ;
    wire \eeprom.n4055 ;
    wire \eeprom.n4056 ;
    wire \eeprom.n2677 ;
    wire \eeprom.n2678 ;
    wire \eeprom.n2710_cascade_ ;
    wire \eeprom.n2686 ;
    wire \eeprom.n2912 ;
    wire \eeprom.n5157_cascade_ ;
    wire \eeprom.n16 ;
    wire \eeprom.n5153 ;
    wire \eeprom.n2918 ;
    wire \eeprom.n2911 ;
    wire \eeprom.n2886 ;
    wire bfn_21_27_0_;
    wire \eeprom.n2885 ;
    wire \eeprom.n4072 ;
    wire \eeprom.n2884 ;
    wire \eeprom.n4073 ;
    wire \eeprom.n2883 ;
    wire \eeprom.n4074 ;
    wire \eeprom.n2882 ;
    wire \eeprom.n4075 ;
    wire \eeprom.n2881 ;
    wire \eeprom.n4076 ;
    wire \eeprom.n2880 ;
    wire \eeprom.n4077 ;
    wire \eeprom.n2879 ;
    wire \eeprom.n4078 ;
    wire \eeprom.n4079 ;
    wire \eeprom.n2878 ;
    wire bfn_21_28_0_;
    wire \eeprom.n2877 ;
    wire \eeprom.n4080 ;
    wire \eeprom.n2876 ;
    wire \eeprom.n4081 ;
    wire \eeprom.n4082 ;
    wire \eeprom.n2874 ;
    wire \eeprom.n4083 ;
    wire \eeprom.n4084 ;
    wire \eeprom.n4085 ;
    wire \eeprom.n4086 ;
    wire \eeprom.n4087 ;
    wire bfn_21_29_0_;
    wire \eeprom.n2902 ;
    wire \eeprom.n2902_cascade_ ;
    wire \eeprom.n19_adj_327 ;
    wire \eeprom.n2872 ;
    wire \eeprom.n2904 ;
    wire \eeprom.n2873 ;
    wire \eeprom.n2905 ;
    wire \eeprom.n2871 ;
    wire \eeprom.n2903 ;
    wire \eeprom.n2875 ;
    wire \eeprom.n2836 ;
    wire \eeprom.n2907 ;
    wire bfn_22_17_0_;
    wire \eeprom.n2285 ;
    wire \eeprom.n3997 ;
    wire \eeprom.n3998 ;
    wire \eeprom.n2283 ;
    wire \eeprom.n3999 ;
    wire \eeprom.n2215 ;
    wire \eeprom.n4000 ;
    wire \eeprom.n2214 ;
    wire \eeprom.n2281 ;
    wire \eeprom.n4001 ;
    wire \eeprom.n4002 ;
    wire \eeprom.n4003 ;
    wire \eeprom.n4004 ;
    wire \eeprom.n2278 ;
    wire bfn_22_18_0_;
    wire \eeprom.n4005 ;
    wire \eeprom.n4006 ;
    wire \eeprom.n2216 ;
    wire \eeprom.n2143_cascade_ ;
    wire \eeprom.n2286 ;
    wire \eeprom.n2218 ;
    wire \eeprom.n5045 ;
    wire \eeprom.n2211 ;
    wire \eeprom.n4797_cascade_ ;
    wire \eeprom.n2242_cascade_ ;
    wire \eeprom.n2282 ;
    wire \eeprom.n5400_cascade_ ;
    wire \eeprom.n2217 ;
    wire \eeprom.n2284 ;
    wire \eeprom.n2280 ;
    wire \eeprom.n2213 ;
    wire \eeprom.n5405 ;
    wire \eeprom.n2316 ;
    wire \eeprom.n2317 ;
    wire \eeprom.n2314 ;
    wire \eeprom.n2318 ;
    wire \eeprom.n5085_cascade_ ;
    wire \eeprom.n2310 ;
    wire \eeprom.n2315 ;
    wire \eeprom.n2313 ;
    wire \eeprom.n5081 ;
    wire \eeprom.n2277 ;
    wire \eeprom.n2309 ;
    wire \eeprom.n2309_cascade_ ;
    wire \eeprom.n2308 ;
    wire \eeprom.n2312 ;
    wire \eeprom.n8_adj_322_cascade_ ;
    wire \eeprom.n7_adj_323 ;
    wire \eeprom.n2341 ;
    wire \eeprom.n2341_cascade_ ;
    wire \eeprom.n5576 ;
    wire \eeprom.n2279 ;
    wire \eeprom.n2311 ;
    wire \eeprom.n5073_cascade_ ;
    wire \eeprom.n4782_cascade_ ;
    wire \eeprom.n12_cascade_ ;
    wire \eeprom.n2440_cascade_ ;
    wire \eeprom.n5071 ;
    wire bfn_22_22_0_;
    wire \eeprom.n4018 ;
    wire \eeprom.n4019 ;
    wire \eeprom.n4020 ;
    wire \eeprom.n4021 ;
    wire \eeprom.n2414 ;
    wire \eeprom.n2481 ;
    wire \eeprom.n4022 ;
    wire \eeprom.n2413 ;
    wire \eeprom.n2480 ;
    wire \eeprom.n4023 ;
    wire \eeprom.n2412 ;
    wire \eeprom.n2479 ;
    wire \eeprom.n4024 ;
    wire \eeprom.n4025 ;
    wire bfn_22_23_0_;
    wire \eeprom.n4026 ;
    wire \eeprom.n2409 ;
    wire \eeprom.n2476 ;
    wire \eeprom.n4027 ;
    wire \eeprom.n4028 ;
    wire \eeprom.n2407 ;
    wire \eeprom.n4029 ;
    wire \eeprom.n2638_cascade_ ;
    wire \eeprom.n2684 ;
    wire \eeprom.n2716_cascade_ ;
    wire \eeprom.n2680 ;
    wire \eeprom.n2679 ;
    wire \eeprom.n2676 ;
    wire \eeprom.n2675 ;
    wire \eeprom.n2673 ;
    wire \eeprom.n2705_cascade_ ;
    wire \eeprom.n17_adj_339 ;
    wire \eeprom.n16_adj_338_cascade_ ;
    wire \eeprom.n2737_cascade_ ;
    wire \eeprom.n2818 ;
    wire bfn_22_25_0_;
    wire \eeprom.n2817 ;
    wire \eeprom.n4057 ;
    wire \eeprom.n2717 ;
    wire \eeprom.n2816 ;
    wire \eeprom.n4058 ;
    wire \eeprom.n2716 ;
    wire \eeprom.n2815 ;
    wire \eeprom.n4059 ;
    wire \eeprom.n2814 ;
    wire \eeprom.n4060 ;
    wire \eeprom.n2813 ;
    wire \eeprom.n4061 ;
    wire \eeprom.n5575 ;
    wire \eeprom.n2812 ;
    wire \eeprom.n4062 ;
    wire \eeprom.n2712 ;
    wire \eeprom.n2811 ;
    wire \eeprom.n4063 ;
    wire \eeprom.n4064 ;
    wire \eeprom.n2711 ;
    wire \eeprom.n2810 ;
    wire bfn_22_26_0_;
    wire \eeprom.n2710 ;
    wire \eeprom.n2809 ;
    wire \eeprom.n4065 ;
    wire \eeprom.n2709 ;
    wire \eeprom.n2808 ;
    wire \eeprom.n4066 ;
    wire \eeprom.n2708 ;
    wire \eeprom.n2807 ;
    wire \eeprom.n4067 ;
    wire \eeprom.n2707 ;
    wire \eeprom.n2806 ;
    wire \eeprom.n4068 ;
    wire \eeprom.n2805 ;
    wire \eeprom.n4069 ;
    wire \eeprom.n2705 ;
    wire \eeprom.n2804 ;
    wire \eeprom.n4070 ;
    wire \eeprom.n2704 ;
    wire \eeprom.n2737 ;
    wire \eeprom.n4071 ;
    wire \eeprom.n2803 ;
    wire \eeprom.n5005_cascade_ ;
    wire \eeprom.n5009_cascade_ ;
    wire \eeprom.n2044_cascade_ ;
    wire \eeprom.n2116_cascade_ ;
    wire bfn_23_18_0_;
    wire \eeprom.n2085 ;
    wire \eeprom.n3980 ;
    wire \eeprom.n2084 ;
    wire \eeprom.n3981 ;
    wire \eeprom.n3982 ;
    wire \eeprom.n2082 ;
    wire \eeprom.n3983 ;
    wire \eeprom.n3984 ;
    wire \eeprom.n2080 ;
    wire \eeprom.n3985 ;
    wire \eeprom.n3986 ;
    wire \eeprom.n3987 ;
    wire bfn_23_19_0_;
    wire \eeprom.n2242 ;
    wire \eeprom.n5501 ;
    wire \eeprom.n2081 ;
    wire \eeprom.n2086 ;
    wire \eeprom.n5061 ;
    wire \eeprom.n2118_cascade_ ;
    wire \eeprom.n4788 ;
    wire \eeprom.n2212 ;
    wire \eeprom.n2019 ;
    wire \eeprom.n3721 ;
    wire \eeprom.n3619 ;
    wire \eeprom.n2219 ;
    wire \eeprom.n3723 ;
    wire \eeprom.n2210 ;
    wire \eeprom.n6_adj_321 ;
    wire \eeprom.n2483 ;
    wire \eeprom.n2416 ;
    wire \eeprom.n2485 ;
    wire \eeprom.n2418 ;
    wire \eeprom.n2477 ;
    wire \eeprom.n2410 ;
    wire \eeprom.n2408 ;
    wire \eeprom.n2475 ;
    wire \eeprom.n2486 ;
    wire \eeprom.n2484 ;
    wire \eeprom.n2417 ;
    wire \eeprom.n2482 ;
    wire \eeprom.n2415 ;
    wire \eeprom.n13_adj_329_cascade_ ;
    wire \eeprom.n2539_cascade_ ;
    wire \eeprom.n2683 ;
    wire \eeprom.n2681 ;
    wire \eeprom.n2713 ;
    wire \eeprom.n2713_cascade_ ;
    wire \eeprom.n2715 ;
    wire \eeprom.n2612 ;
    wire \eeprom.n2611 ;
    wire \eeprom.n2612_cascade_ ;
    wire \eeprom.n2610 ;
    wire \eeprom.n16_adj_334 ;
    wire \eeprom.n2618 ;
    wire \eeprom.n12_adj_333 ;
    wire \eeprom.n2606 ;
    wire \eeprom.n2606_cascade_ ;
    wire \eeprom.n10_adj_332 ;
    wire \eeprom.n2718 ;
    wire \eeprom.n5213 ;
    wire \eeprom.n5215 ;
    wire \eeprom.n4830 ;
    wire \eeprom.n2682 ;
    wire \eeprom.n2714 ;
    wire \eeprom.n2609 ;
    wire \eeprom.n3319 ;
    wire \eeprom.n2608 ;
    wire \eeprom.n2607 ;
    wire \eeprom.n2674 ;
    wire \eeprom.n2607_cascade_ ;
    wire \eeprom.n2638 ;
    wire \eeprom.n2706 ;
    wire \eeprom.n2719 ;
    wire \eeprom.n2919 ;
    wire \eeprom.n2419 ;
    wire \eeprom.n3119 ;
    wire \eeprom.n2186 ;
    wire bfn_24_17_0_;
    wire \eeprom.n2118 ;
    wire \eeprom.n2185 ;
    wire \eeprom.n3988 ;
    wire \eeprom.n2117 ;
    wire \eeprom.n2184 ;
    wire \eeprom.n3989 ;
    wire \eeprom.n2116 ;
    wire \eeprom.n2183 ;
    wire \eeprom.n3990 ;
    wire \eeprom.n2182 ;
    wire \eeprom.n3991 ;
    wire \eeprom.n2114 ;
    wire \eeprom.n2181 ;
    wire \eeprom.n3992 ;
    wire \eeprom.n2180 ;
    wire \eeprom.n3993 ;
    wire \eeprom.n2112 ;
    wire \eeprom.n2179 ;
    wire \eeprom.n3994 ;
    wire \eeprom.n3995 ;
    wire \eeprom.n2178 ;
    wire bfn_24_18_0_;
    wire \eeprom.n2110 ;
    wire \eeprom.n2143 ;
    wire \eeprom.n3996 ;
    wire \eeprom.n2209 ;
    wire \eeprom.n3724 ;
    wire \eeprom.n2015 ;
    wire \eeprom.n2079 ;
    wire \eeprom.n2111 ;
    wire \eeprom.n2018 ;
    wire \eeprom.n1945_cascade_ ;
    wire \eeprom.n2017 ;
    wire \eeprom.n2014 ;
    wire \eeprom.n2016 ;
    wire \eeprom.n2083 ;
    wire \eeprom.n2016_cascade_ ;
    wire \eeprom.n2044 ;
    wire \eeprom.n2115 ;
    wire \eeprom.n2115_cascade_ ;
    wire \eeprom.n2113 ;
    wire \eeprom.n5059 ;
    wire \eeprom.n2013 ;
    wire \eeprom.n2012 ;
    wire \eeprom.n1986 ;
    wire bfn_24_20_0_;
    wire \eeprom.n1985 ;
    wire \eeprom.n3973 ;
    wire \eeprom.n1984 ;
    wire \eeprom.n3974 ;
    wire \eeprom.n1983 ;
    wire \eeprom.n3975 ;
    wire \eeprom.n1982 ;
    wire \eeprom.n3976 ;
    wire \eeprom.n1981 ;
    wire \eeprom.n3977 ;
    wire \eeprom.n1980 ;
    wire \eeprom.n3978 ;
    wire \eeprom.n1945 ;
    wire \eeprom.n3979 ;
    wire \eeprom.n2011 ;
    wire \eeprom.n2411 ;
    wire \eeprom.n2478 ;
    wire \eeprom.n2440 ;
    wire \eeprom.n3419 ;
    wire \eeprom.n5169_cascade_ ;
    wire \eeprom.n5173_cascade_ ;
    wire \eeprom.n11_adj_328 ;
    wire \eeprom.n2615 ;
    wire \eeprom.n2615_cascade_ ;
    wire \eeprom.n2613 ;
    wire \eeprom.n2617 ;
    wire \eeprom.n2614 ;
    wire \eeprom.n5101_cascade_ ;
    wire \eeprom.n2616 ;
    wire \eeprom.n5105 ;
    wire \eeprom.n2586 ;
    wire bfn_24_23_0_;
    wire \eeprom.n2518 ;
    wire \eeprom.n2585 ;
    wire \eeprom.n4030 ;
    wire \eeprom.n2517 ;
    wire \eeprom.n2584 ;
    wire \eeprom.n4031 ;
    wire \eeprom.n2516 ;
    wire \eeprom.n2583 ;
    wire \eeprom.n4032 ;
    wire \eeprom.n2515 ;
    wire \eeprom.n2582 ;
    wire \eeprom.n4033 ;
    wire \eeprom.n2514 ;
    wire \eeprom.n2581 ;
    wire \eeprom.n4034 ;
    wire \eeprom.n2513 ;
    wire \eeprom.n2580 ;
    wire \eeprom.n4035 ;
    wire \eeprom.n2512 ;
    wire \eeprom.n2579 ;
    wire \eeprom.n4036 ;
    wire \eeprom.n4037 ;
    wire \eeprom.n2511 ;
    wire \eeprom.n2578 ;
    wire bfn_24_24_0_;
    wire \eeprom.n2510 ;
    wire \eeprom.n2577 ;
    wire \eeprom.n4038 ;
    wire \eeprom.n2509 ;
    wire \eeprom.n2576 ;
    wire \eeprom.n4039 ;
    wire \eeprom.n2508 ;
    wire \eeprom.n2575 ;
    wire \eeprom.n4040 ;
    wire \eeprom.n2507 ;
    wire \eeprom.n2574 ;
    wire \eeprom.n4041 ;
    wire \eeprom.n2539 ;
    wire \eeprom.n2506 ;
    wire \eeprom.n4042 ;
    wire \eeprom.n2605 ;
    wire \eeprom.n2519 ;
    wire \eeprom.n2619 ;
    wire \eeprom.n2819 ;
    wire \eeprom.n3219 ;
    wire \eeprom.n3019 ;
    wire n1805_cascade_;
    wire n170;
    wire n1800_cascade_;
    wire n164;
    wire n4_adj_361;
    wire n4_adj_361_cascade_;
    wire n162;
    wire n5361_cascade_;
    wire n172;
    wire n22_adj_367_cascade_;
    wire n4_adj_369_cascade_;
    wire n4_cascade_;
    wire n166;
    wire n4;
    wire n168;
    wire n1805;
    wire n158;
    wire n8;
    wire n5461_cascade_;
    wire n1800;
    wire n3585;
    wire n160;
    wire \eeprom.n2119 ;
    wire \eeprom.n2319 ;
    wire bfn_26_21_0_;
    wire \eeprom.n3931 ;
    wire \eeprom.eeprom_counter_2 ;
    wire \eeprom.n3932 ;
    wire \eeprom.n3933 ;
    wire \eeprom.eeprom_counter_4 ;
    wire \eeprom.n3934 ;
    wire \eeprom.n3935 ;
    wire \eeprom.n3936 ;
    wire \eeprom.n3937 ;
    wire \eeprom.n3938 ;
    wire bfn_26_22_0_;
    wire \eeprom.n3939 ;
    wire \eeprom.n3940 ;
    wire \eeprom.n3941 ;
    wire \eeprom.n3942 ;
    wire \eeprom.eeprom_counter_13 ;
    wire \eeprom.n3943 ;
    wire \eeprom.n3944 ;
    wire \eeprom.n3945 ;
    wire \eeprom.n3946 ;
    wire bfn_26_23_0_;
    wire \eeprom.n3947 ;
    wire \eeprom.n3948 ;
    wire \eeprom.n3949 ;
    wire \eeprom.eeprom_counter_20 ;
    wire \eeprom.n3950 ;
    wire \eeprom.n3951 ;
    wire \eeprom.n3952 ;
    wire \eeprom.n3953 ;
    wire \eeprom.n3954 ;
    wire bfn_26_24_0_;
    wire \eeprom.n3955 ;
    wire \eeprom.n3956 ;
    wire \eeprom.n3957 ;
    wire \eeprom.n3958 ;
    wire \eeprom.n3959 ;
    wire \eeprom.n3960 ;
    wire \eeprom.n3961 ;
    wire \eeprom.eeprom_counter_23 ;
    wire \eeprom.eeprom_counter_16 ;
    wire \eeprom.n1919 ;
    wire \eeprom.eeprom_counter_24 ;
    wire \eeprom.eeprom_counter_18 ;
    wire \eeprom.eeprom_counter_17 ;
    wire \eeprom.eeprom_counter_22 ;
    wire \eeprom.eeprom_counter_21 ;
    wire bfn_27_17_0_;
    wire \eeprom.i2c.n3899 ;
    wire \eeprom.i2c.n3900 ;
    wire \eeprom.i2c.n3901 ;
    wire \eeprom.i2c.n3902 ;
    wire \eeprom.i2c.n3903 ;
    wire \eeprom.i2c.n3904 ;
    wire \eeprom.i2c.n3905 ;
    wire n11;
    wire n10_adj_360;
    wire n4733;
    wire \eeprom.i2c.n1913 ;
    wire \eeprom.i2c.n534 ;
    wire \eeprom.i2c.n1829 ;
    wire \eeprom.i2c.n9 ;
    wire \eeprom.i2c.n9_cascade_ ;
    wire n1814;
    wire n1814_cascade_;
    wire \eeprom.i2c.n37 ;
    wire \eeprom.i2c.n37_cascade_ ;
    wire \eeprom.i2c.n33 ;
    wire \eeprom.i2c.n39_cascade_ ;
    wire \eeprom.i2c.n39 ;
    wire \eeprom.i2c.n407_cascade_ ;
    wire \eeprom.n917 ;
    wire \eeprom.eeprom_counter_5 ;
    wire \eeprom.n3722 ;
    wire \eeprom.eeprom_counter_30 ;
    wire \eeprom.n1256_cascade_ ;
    wire \eeprom.n1913 ;
    wire \eeprom.i2c.n13 ;
    wire \eeprom.eeprom_counter_7 ;
    wire \INVeeprom.i2c.i2c_scl_enable_124C_net ;
    wire \eeprom.n1918 ;
    wire \eeprom.eeprom_counter_0 ;
    wire \eeprom.n1912 ;
    wire \eeprom.eeprom_counter_27 ;
    wire \eeprom.n1139_cascade_ ;
    wire \eeprom.eeprom_counter_3 ;
    wire \eeprom.n1916 ;
    wire \eeprom.n5035_cascade_ ;
    wire \eeprom.n5039 ;
    wire \eeprom.eeprom_counter_12 ;
    wire \eeprom.eeprom_counter_1 ;
    wire \eeprom.n892_cascade_ ;
    wire \eeprom.eeprom_counter_10 ;
    wire \eeprom.eeprom_counter_28 ;
    wire \eeprom.n1138_cascade_ ;
    wire \eeprom.n33_adj_289 ;
    wire \eeprom.n33 ;
    wire bfn_27_23_0_;
    wire \eeprom.n32_adj_288 ;
    wire \eeprom.n32_adj_287 ;
    wire \eeprom.n4242 ;
    wire \eeprom.n31_adj_286 ;
    wire \eeprom.n31_adj_285 ;
    wire \eeprom.n4243 ;
    wire \eeprom.n30_adj_277 ;
    wire \eeprom.n30_adj_284 ;
    wire \eeprom.n4244 ;
    wire \eeprom.n29_adj_278 ;
    wire \eeprom.n29_adj_283 ;
    wire \eeprom.n4245 ;
    wire \eeprom.n28_adj_279 ;
    wire \eeprom.n28_adj_282 ;
    wire \eeprom.n4246 ;
    wire \eeprom.n27_adj_280 ;
    wire \eeprom.n4247 ;
    wire \eeprom.n26_adj_276 ;
    wire \eeprom.n26_adj_275 ;
    wire \eeprom.n4248 ;
    wire \eeprom.n4249 ;
    wire bfn_27_24_0_;
    wire \eeprom.n24_adj_269 ;
    wire \eeprom.n4250 ;
    wire \eeprom.n23_adj_268 ;
    wire \eeprom.n23 ;
    wire \eeprom.n4251 ;
    wire \eeprom.n22_adj_265 ;
    wire \eeprom.n4252 ;
    wire \eeprom.n21_adj_264 ;
    wire \eeprom.n21 ;
    wire \eeprom.n4253 ;
    wire \eeprom.n20_adj_259 ;
    wire \eeprom.n20 ;
    wire \eeprom.n4254 ;
    wire \eeprom.n19_adj_320 ;
    wire \eeprom.n4255 ;
    wire \eeprom.n18_adj_326 ;
    wire \eeprom.n4256 ;
    wire \eeprom.n4257 ;
    wire \eeprom.n17 ;
    wire \eeprom.n17_adj_324 ;
    wire bfn_27_25_0_;
    wire \eeprom.n16_adj_294 ;
    wire \eeprom.n16_adj_325 ;
    wire \eeprom.n4258 ;
    wire \eeprom.n15_adj_295 ;
    wire \eeprom.n15 ;
    wire \eeprom.n4259 ;
    wire \eeprom.n14 ;
    wire \eeprom.n4260 ;
    wire \eeprom.n13 ;
    wire \eeprom.n13_adj_318 ;
    wire \eeprom.n4261 ;
    wire \eeprom.n12_adj_298 ;
    wire \eeprom.n12_adj_319 ;
    wire \eeprom.n4262 ;
    wire \eeprom.n11_adj_299 ;
    wire \eeprom.n11 ;
    wire \eeprom.n4263 ;
    wire \eeprom.n10 ;
    wire \eeprom.n10_adj_343 ;
    wire \eeprom.n4264 ;
    wire \eeprom.n4265 ;
    wire \eeprom.n9 ;
    wire \eeprom.n9_adj_308 ;
    wire bfn_27_26_0_;
    wire \eeprom.n8_adj_311 ;
    wire \eeprom.n4266 ;
    wire \eeprom.n7 ;
    wire \eeprom.n4267 ;
    wire \eeprom.n6 ;
    wire \eeprom.n6_adj_306 ;
    wire \eeprom.n4268 ;
    wire \eeprom.n5 ;
    wire \eeprom.n5_adj_317 ;
    wire \eeprom.n4269 ;
    wire \eeprom.n4 ;
    wire \eeprom.n4270 ;
    wire \eeprom.n3 ;
    wire \eeprom.n3_adj_312 ;
    wire \eeprom.n4271 ;
    wire \eeprom.n2 ;
    wire \eeprom.n4272 ;
    wire \eeprom.i2c.counter_3 ;
    wire \eeprom.i2c.counter_5 ;
    wire \eeprom.i2c.counter_4 ;
    wire \eeprom.i2c.counter_7 ;
    wire \eeprom.i2c.counter_6 ;
    wire \eeprom.i2c.n12_cascade_ ;
    wire \eeprom.i2c.n464 ;
    wire n4_adj_358;
    wire n10_cascade_;
    wire state_7_N_162_3;
    wire \eeprom.i2c.n4579 ;
    wire n11_adj_359;
    wire n5458;
    wire n6_adj_365_cascade_;
    wire n471;
    wire state_3;
    wire n3587;
    wire n3587_cascade_;
    wire n10;
    wire n5454;
    wire \eeprom.i2c.counter_1 ;
    wire \eeprom.i2c.counter_2 ;
    wire \eeprom.i2c.counter_0 ;
    wire \eeprom.i2c.n5464_cascade_ ;
    wire \eeprom.i2c.n5451_cascade_ ;
    wire \eeprom.i2c.sda_out ;
    wire \INVeeprom.i2c.sda_out_133C_net ;
    wire \eeprom.i2c.n4513 ;
    wire state_2;
    wire n3595;
    wire state_1;
    wire n3581;
    wire \eeprom.i2c.n407 ;
    wire state_0;
    wire sda_enable;
    wire \INVeeprom.i2c.write_enable_132C_net ;
    wire \eeprom.i2c.n524 ;
    wire \eeprom.i2c.n1901 ;
    wire \eeprom.n892 ;
    wire \eeprom.n1198 ;
    wire bfn_28_21_0_;
    wire \eeprom.n4273 ;
    wire \eeprom.n1139 ;
    wire \eeprom.n1196 ;
    wire \eeprom.n4274 ;
    wire \eeprom.n4275 ;
    wire \eeprom.n4276 ;
    wire \eeprom.n5327 ;
    wire \eeprom.n5328 ;
    wire \eeprom.n4277 ;
    wire \eeprom.n4278 ;
    wire \eeprom.n1192 ;
    wire \eeprom.n1256 ;
    wire \eeprom.n1843_cascade_ ;
    wire \eeprom.n1195 ;
    wire \eeprom.n1915 ;
    wire \eeprom.eeprom_counter_29 ;
    wire \eeprom.n4_adj_310 ;
    wire \eeprom.n1138 ;
    wire \eeprom.n1137_cascade_ ;
    wire \eeprom.n4977 ;
    wire \eeprom.n4983 ;
    wire \eeprom.n1197 ;
    wire \eeprom.n1917 ;
    wire \eeprom.n1194 ;
    wire \eeprom.n1137 ;
    wire \eeprom.n1843 ;
    wire \eeprom.n1914 ;
    wire \eeprom.eeprom_counter_14 ;
    wire \eeprom.n19 ;
    wire \eeprom.n25_adj_271 ;
    wire \eeprom.n3519 ;
    wire \eeprom.n27_adj_281 ;
    wire \eeprom.eeprom_counter_6 ;
    wire \eeprom.n3719 ;
    wire \eeprom.eeprom_counter_19 ;
    wire \eeprom.n14_adj_297 ;
    wire \eeprom.eeprom_counter_26 ;
    wire \eeprom.n7_adj_309 ;
    wire \eeprom.n1140 ;
    wire \eeprom.eeprom_counter_8 ;
    wire \eeprom.n25_adj_272 ;
    wire \eeprom.eeprom_counter_31 ;
    wire \eeprom.n2_adj_307 ;
    wire \eeprom.n1135 ;
    wire CONSTANT_ONE_NET;
    wire n174;
    wire rw;
    wire saved_addr_0;
    wire state_7_N_146_0;
    wire \eeprom.enable ;
    wire \eeprom.i2c.n1832 ;
    wire \eeprom.i2c.n6_adj_255_cascade_ ;
    wire \eeprom.eeprom_counter_9 ;
    wire \eeprom.n24_adj_270 ;
    wire \eeprom.i2c.i2c_clk ;
    wire scl_enable;
    wire scl_c;
    wire \eeprom.eeprom_counter_11 ;
    wire \eeprom.n22_adj_266 ;
    wire \eeprom.eeprom_counter_25 ;
    wire \eeprom.n8 ;
    wire \eeprom.eeprom_counter_15 ;
    wire \eeprom.n18_adj_293 ;
    wire \eeprom.i2c.counter2_0 ;
    wire bfn_30_20_0_;
    wire \eeprom.i2c.counter2_1 ;
    wire \eeprom.i2c.n3962 ;
    wire \eeprom.i2c.counter2_2 ;
    wire \eeprom.i2c.n3963 ;
    wire \eeprom.i2c.counter2_3 ;
    wire \eeprom.i2c.n3964 ;
    wire \eeprom.i2c.n3965 ;
    wire \eeprom.i2c.counter2_4 ;
    wire _gnd_net_;
    wire CLK_N;
    wire \eeprom.i2c.counter2_7__N_133 ;

    defparam CS_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_CLK_pad_iopad (
            .OE(N__30138),
            .DIN(N__30137),
            .DOUT(N__30136),
            .PACKAGEPIN(CS_CLK));
    defparam CS_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_CLK_pad_preio (
            .PADOEN(N__30138),
            .PADOUT(N__30137),
            .PADIN(N__30136),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_pad_iopad (
            .OE(N__30129),
            .DIN(N__30128),
            .DOUT(N__30127),
            .PACKAGEPIN(CS));
    defparam CS_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_pad_preio (
            .PADOEN(N__30129),
            .PADOUT(N__30128),
            .PADIN(N__30127),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam DE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DE_pad_iopad.PULLUP=1'b0;
    IO_PAD DE_pad_iopad (
            .OE(N__30120),
            .DIN(N__30119),
            .DOUT(N__30118),
            .PACKAGEPIN(DE));
    defparam DE_pad_preio.PIN_TYPE=6'b011001;
    defparam DE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DE_pad_preio (
            .PADOEN(N__30120),
            .PADOUT(N__30119),
            .PADIN(N__30118),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHA_pad_iopad.PULLUP=1'b0;
    IO_PAD INHA_pad_iopad (
            .OE(N__30111),
            .DIN(N__30110),
            .DOUT(N__30109),
            .PACKAGEPIN(INHA));
    defparam INHA_pad_preio.PIN_TYPE=6'b011001;
    defparam INHA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHA_pad_preio (
            .PADOEN(N__30111),
            .PADOUT(N__30110),
            .PADIN(N__30109),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHB_pad_iopad.PULLUP=1'b0;
    IO_PAD INHB_pad_iopad (
            .OE(N__30102),
            .DIN(N__30101),
            .DOUT(N__30100),
            .PACKAGEPIN(INHB));
    defparam INHB_pad_preio.PIN_TYPE=6'b011001;
    defparam INHB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHB_pad_preio (
            .PADOEN(N__30102),
            .PADOUT(N__30101),
            .PADIN(N__30100),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHC_pad_iopad.PULLUP=1'b0;
    IO_PAD INHC_pad_iopad (
            .OE(N__30093),
            .DIN(N__30092),
            .DOUT(N__30091),
            .PACKAGEPIN(INHC));
    defparam INHC_pad_preio.PIN_TYPE=6'b011001;
    defparam INHC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHC_pad_preio (
            .PADOEN(N__30093),
            .PADOUT(N__30092),
            .PADIN(N__30091),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLA_pad_iopad.PULLUP=1'b0;
    IO_PAD INLA_pad_iopad (
            .OE(N__30084),
            .DIN(N__30083),
            .DOUT(N__30082),
            .PACKAGEPIN(INLA));
    defparam INLA_pad_preio.PIN_TYPE=6'b011001;
    defparam INLA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLA_pad_preio (
            .PADOEN(N__30084),
            .PADOUT(N__30083),
            .PADIN(N__30082),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLB_pad_iopad.PULLUP=1'b0;
    IO_PAD INLB_pad_iopad (
            .OE(N__30075),
            .DIN(N__30074),
            .DOUT(N__30073),
            .PACKAGEPIN(INLB));
    defparam INLB_pad_preio.PIN_TYPE=6'b011001;
    defparam INLB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLB_pad_preio (
            .PADOEN(N__30075),
            .PADOUT(N__30074),
            .PADIN(N__30073),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLC_pad_iopad.PULLUP=1'b0;
    IO_PAD INLC_pad_iopad (
            .OE(N__30066),
            .DIN(N__30065),
            .DOUT(N__30064),
            .PACKAGEPIN(INLC));
    defparam INLC_pad_preio.PIN_TYPE=6'b011001;
    defparam INLC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLC_pad_preio (
            .PADOEN(N__30066),
            .PADOUT(N__30065),
            .PADIN(N__30064),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__30057),
            .DIN(N__30056),
            .DOUT(N__30055),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__30057),
            .PADOUT(N__30056),
            .PADIN(N__30055),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11906),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__30048),
            .DIN(N__30047),
            .DOUT(N__30046),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__30048),
            .PADOUT(N__30047),
            .PADIN(N__30046),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TX_pad_iopad.PULLUP=1'b0;
    IO_PAD TX_pad_iopad (
            .OE(N__30039),
            .DIN(N__30038),
            .DOUT(N__30037),
            .PACKAGEPIN(TX));
    defparam TX_pad_preio.PIN_TYPE=6'b011001;
    defparam TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TX_pad_preio (
            .PADOEN(N__30039),
            .PADOUT(N__30038),
            .PADIN(N__30037),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__30030),
            .DIN(N__30029),
            .DOUT(N__30028),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__30030),
            .PADOUT(N__30029),
            .PADIN(N__30028),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam scl_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam scl_output_iopad.PULLUP=1'b1;
    IO_PAD scl_output_iopad (
            .OE(N__30021),
            .DIN(N__30020),
            .DOUT(N__30019),
            .PACKAGEPIN(SCL));
    defparam scl_output_preio.PIN_TYPE=6'b101001;
    defparam scl_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO scl_output_preio (
            .PADOEN(N__30021),
            .PADOUT(N__30020),
            .PADIN(N__30019),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29558),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__29585));
    defparam sda_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sda_output_iopad.PULLUP=1'b1;
    IO_PAD sda_output_iopad (
            .OE(N__30012),
            .DIN(N__30011),
            .DOUT(N__30010),
            .PACKAGEPIN(SDA));
    defparam sda_output_preio.PIN_TYPE=6'b101001;
    defparam sda_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO sda_output_preio (
            .PADOEN(N__30012),
            .PADOUT(N__30011),
            .PADIN(N__30010),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26531),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__27311));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__30003),
            .DIN(N__30002),
            .DOUT(N__30001),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__30003),
            .PADOUT(N__30002),
            .PADIN(N__30001),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__7050 (
            .O(N__29984),
            .I(N__29980));
    InMux I__7049 (
            .O(N__29983),
            .I(N__29977));
    LocalMux I__7048 (
            .O(N__29980),
            .I(N__29973));
    LocalMux I__7047 (
            .O(N__29977),
            .I(N__29970));
    InMux I__7046 (
            .O(N__29976),
            .I(N__29967));
    Span4Mux_h I__7045 (
            .O(N__29973),
            .I(N__29962));
    Span4Mux_h I__7044 (
            .O(N__29970),
            .I(N__29962));
    LocalMux I__7043 (
            .O(N__29967),
            .I(\eeprom.eeprom_counter_15 ));
    Odrv4 I__7042 (
            .O(N__29962),
            .I(\eeprom.eeprom_counter_15 ));
    CascadeMux I__7041 (
            .O(N__29957),
            .I(N__29954));
    InMux I__7040 (
            .O(N__29954),
            .I(N__29951));
    LocalMux I__7039 (
            .O(N__29951),
            .I(N__29948));
    Span4Mux_v I__7038 (
            .O(N__29948),
            .I(N__29945));
    Odrv4 I__7037 (
            .O(N__29945),
            .I(\eeprom.n18_adj_293 ));
    InMux I__7036 (
            .O(N__29942),
            .I(N__29938));
    InMux I__7035 (
            .O(N__29941),
            .I(N__29935));
    LocalMux I__7034 (
            .O(N__29938),
            .I(\eeprom.i2c.counter2_0 ));
    LocalMux I__7033 (
            .O(N__29935),
            .I(\eeprom.i2c.counter2_0 ));
    InMux I__7032 (
            .O(N__29930),
            .I(bfn_30_20_0_));
    InMux I__7031 (
            .O(N__29927),
            .I(N__29923));
    InMux I__7030 (
            .O(N__29926),
            .I(N__29920));
    LocalMux I__7029 (
            .O(N__29923),
            .I(\eeprom.i2c.counter2_1 ));
    LocalMux I__7028 (
            .O(N__29920),
            .I(\eeprom.i2c.counter2_1 ));
    InMux I__7027 (
            .O(N__29915),
            .I(\eeprom.i2c.n3962 ));
    InMux I__7026 (
            .O(N__29912),
            .I(N__29908));
    InMux I__7025 (
            .O(N__29911),
            .I(N__29905));
    LocalMux I__7024 (
            .O(N__29908),
            .I(\eeprom.i2c.counter2_2 ));
    LocalMux I__7023 (
            .O(N__29905),
            .I(\eeprom.i2c.counter2_2 ));
    InMux I__7022 (
            .O(N__29900),
            .I(\eeprom.i2c.n3963 ));
    InMux I__7021 (
            .O(N__29897),
            .I(N__29893));
    InMux I__7020 (
            .O(N__29896),
            .I(N__29890));
    LocalMux I__7019 (
            .O(N__29893),
            .I(\eeprom.i2c.counter2_3 ));
    LocalMux I__7018 (
            .O(N__29890),
            .I(\eeprom.i2c.counter2_3 ));
    InMux I__7017 (
            .O(N__29885),
            .I(\eeprom.i2c.n3964 ));
    InMux I__7016 (
            .O(N__29882),
            .I(\eeprom.i2c.n3965 ));
    InMux I__7015 (
            .O(N__29879),
            .I(N__29875));
    InMux I__7014 (
            .O(N__29878),
            .I(N__29872));
    LocalMux I__7013 (
            .O(N__29875),
            .I(\eeprom.i2c.counter2_4 ));
    LocalMux I__7012 (
            .O(N__29872),
            .I(\eeprom.i2c.counter2_4 ));
    ClkMux I__7011 (
            .O(N__29867),
            .I(N__29831));
    ClkMux I__7010 (
            .O(N__29866),
            .I(N__29831));
    ClkMux I__7009 (
            .O(N__29865),
            .I(N__29831));
    ClkMux I__7008 (
            .O(N__29864),
            .I(N__29831));
    ClkMux I__7007 (
            .O(N__29863),
            .I(N__29831));
    ClkMux I__7006 (
            .O(N__29862),
            .I(N__29831));
    ClkMux I__7005 (
            .O(N__29861),
            .I(N__29831));
    ClkMux I__7004 (
            .O(N__29860),
            .I(N__29831));
    ClkMux I__7003 (
            .O(N__29859),
            .I(N__29831));
    ClkMux I__7002 (
            .O(N__29858),
            .I(N__29831));
    ClkMux I__7001 (
            .O(N__29857),
            .I(N__29831));
    ClkMux I__7000 (
            .O(N__29856),
            .I(N__29831));
    GlobalMux I__6999 (
            .O(N__29831),
            .I(N__29828));
    gio2CtrlBuf I__6998 (
            .O(N__29828),
            .I(CLK_N));
    SRMux I__6997 (
            .O(N__29825),
            .I(N__29821));
    InMux I__6996 (
            .O(N__29824),
            .I(N__29818));
    LocalMux I__6995 (
            .O(N__29821),
            .I(N__29813));
    LocalMux I__6994 (
            .O(N__29818),
            .I(N__29810));
    InMux I__6993 (
            .O(N__29817),
            .I(N__29805));
    InMux I__6992 (
            .O(N__29816),
            .I(N__29805));
    Odrv4 I__6991 (
            .O(N__29813),
            .I(\eeprom.i2c.counter2_7__N_133 ));
    Odrv4 I__6990 (
            .O(N__29810),
            .I(\eeprom.i2c.counter2_7__N_133 ));
    LocalMux I__6989 (
            .O(N__29805),
            .I(\eeprom.i2c.counter2_7__N_133 ));
    InMux I__6988 (
            .O(N__29798),
            .I(N__29794));
    InMux I__6987 (
            .O(N__29797),
            .I(N__29791));
    LocalMux I__6986 (
            .O(N__29794),
            .I(state_7_N_146_0));
    LocalMux I__6985 (
            .O(N__29791),
            .I(state_7_N_146_0));
    SRMux I__6984 (
            .O(N__29786),
            .I(N__29782));
    InMux I__6983 (
            .O(N__29785),
            .I(N__29778));
    LocalMux I__6982 (
            .O(N__29782),
            .I(N__29775));
    InMux I__6981 (
            .O(N__29781),
            .I(N__29772));
    LocalMux I__6980 (
            .O(N__29778),
            .I(N__29769));
    Span4Mux_v I__6979 (
            .O(N__29775),
            .I(N__29764));
    LocalMux I__6978 (
            .O(N__29772),
            .I(N__29764));
    Span4Mux_v I__6977 (
            .O(N__29769),
            .I(N__29759));
    Span4Mux_h I__6976 (
            .O(N__29764),
            .I(N__29759));
    Span4Mux_h I__6975 (
            .O(N__29759),
            .I(N__29756));
    Odrv4 I__6974 (
            .O(N__29756),
            .I(\eeprom.enable ));
    CEMux I__6973 (
            .O(N__29753),
            .I(N__29750));
    LocalMux I__6972 (
            .O(N__29750),
            .I(N__29747));
    Span4Mux_h I__6971 (
            .O(N__29747),
            .I(N__29744));
    Odrv4 I__6970 (
            .O(N__29744),
            .I(\eeprom.i2c.n1832 ));
    CascadeMux I__6969 (
            .O(N__29741),
            .I(\eeprom.i2c.n6_adj_255_cascade_ ));
    InMux I__6968 (
            .O(N__29738),
            .I(N__29734));
    InMux I__6967 (
            .O(N__29737),
            .I(N__29731));
    LocalMux I__6966 (
            .O(N__29734),
            .I(N__29727));
    LocalMux I__6965 (
            .O(N__29731),
            .I(N__29724));
    InMux I__6964 (
            .O(N__29730),
            .I(N__29721));
    Span4Mux_v I__6963 (
            .O(N__29727),
            .I(N__29716));
    Span4Mux_v I__6962 (
            .O(N__29724),
            .I(N__29716));
    LocalMux I__6961 (
            .O(N__29721),
            .I(\eeprom.eeprom_counter_9 ));
    Odrv4 I__6960 (
            .O(N__29716),
            .I(\eeprom.eeprom_counter_9 ));
    CascadeMux I__6959 (
            .O(N__29711),
            .I(N__29708));
    InMux I__6958 (
            .O(N__29708),
            .I(N__29705));
    LocalMux I__6957 (
            .O(N__29705),
            .I(N__29702));
    Span4Mux_h I__6956 (
            .O(N__29702),
            .I(N__29699));
    Odrv4 I__6955 (
            .O(N__29699),
            .I(\eeprom.n24_adj_270 ));
    ClkMux I__6954 (
            .O(N__29696),
            .I(N__29690));
    ClkMux I__6953 (
            .O(N__29695),
            .I(N__29684));
    ClkMux I__6952 (
            .O(N__29694),
            .I(N__29680));
    ClkMux I__6951 (
            .O(N__29693),
            .I(N__29677));
    LocalMux I__6950 (
            .O(N__29690),
            .I(N__29674));
    ClkMux I__6949 (
            .O(N__29689),
            .I(N__29671));
    ClkMux I__6948 (
            .O(N__29688),
            .I(N__29668));
    ClkMux I__6947 (
            .O(N__29687),
            .I(N__29665));
    LocalMux I__6946 (
            .O(N__29684),
            .I(N__29662));
    ClkMux I__6945 (
            .O(N__29683),
            .I(N__29659));
    LocalMux I__6944 (
            .O(N__29680),
            .I(N__29651));
    LocalMux I__6943 (
            .O(N__29677),
            .I(N__29651));
    Span4Mux_v I__6942 (
            .O(N__29674),
            .I(N__29646));
    LocalMux I__6941 (
            .O(N__29671),
            .I(N__29646));
    LocalMux I__6940 (
            .O(N__29668),
            .I(N__29641));
    LocalMux I__6939 (
            .O(N__29665),
            .I(N__29641));
    Span4Mux_h I__6938 (
            .O(N__29662),
            .I(N__29636));
    LocalMux I__6937 (
            .O(N__29659),
            .I(N__29636));
    ClkMux I__6936 (
            .O(N__29658),
            .I(N__29633));
    InMux I__6935 (
            .O(N__29657),
            .I(N__29629));
    ClkMux I__6934 (
            .O(N__29656),
            .I(N__29626));
    Span4Mux_v I__6933 (
            .O(N__29651),
            .I(N__29619));
    Span4Mux_v I__6932 (
            .O(N__29646),
            .I(N__29619));
    Span4Mux_h I__6931 (
            .O(N__29641),
            .I(N__29616));
    Span4Mux_v I__6930 (
            .O(N__29636),
            .I(N__29611));
    LocalMux I__6929 (
            .O(N__29633),
            .I(N__29611));
    InMux I__6928 (
            .O(N__29632),
            .I(N__29608));
    LocalMux I__6927 (
            .O(N__29629),
            .I(N__29603));
    LocalMux I__6926 (
            .O(N__29626),
            .I(N__29603));
    InMux I__6925 (
            .O(N__29625),
            .I(N__29598));
    InMux I__6924 (
            .O(N__29624),
            .I(N__29598));
    Odrv4 I__6923 (
            .O(N__29619),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__6922 (
            .O(N__29616),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__6921 (
            .O(N__29611),
            .I(\eeprom.i2c.i2c_clk ));
    LocalMux I__6920 (
            .O(N__29608),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__6919 (
            .O(N__29603),
            .I(\eeprom.i2c.i2c_clk ));
    LocalMux I__6918 (
            .O(N__29598),
            .I(\eeprom.i2c.i2c_clk ));
    IoInMux I__6917 (
            .O(N__29585),
            .I(N__29582));
    LocalMux I__6916 (
            .O(N__29582),
            .I(N__29579));
    IoSpan4Mux I__6915 (
            .O(N__29579),
            .I(N__29575));
    InMux I__6914 (
            .O(N__29578),
            .I(N__29572));
    Span4Mux_s2_h I__6913 (
            .O(N__29575),
            .I(N__29569));
    LocalMux I__6912 (
            .O(N__29572),
            .I(N__29566));
    Span4Mux_v I__6911 (
            .O(N__29569),
            .I(N__29561));
    Span4Mux_v I__6910 (
            .O(N__29566),
            .I(N__29561));
    Odrv4 I__6909 (
            .O(N__29561),
            .I(scl_enable));
    IoInMux I__6908 (
            .O(N__29558),
            .I(N__29555));
    LocalMux I__6907 (
            .O(N__29555),
            .I(N__29552));
    Odrv12 I__6906 (
            .O(N__29552),
            .I(scl_c));
    InMux I__6905 (
            .O(N__29549),
            .I(N__29546));
    LocalMux I__6904 (
            .O(N__29546),
            .I(N__29541));
    InMux I__6903 (
            .O(N__29545),
            .I(N__29538));
    InMux I__6902 (
            .O(N__29544),
            .I(N__29535));
    Span4Mux_h I__6901 (
            .O(N__29541),
            .I(N__29532));
    LocalMux I__6900 (
            .O(N__29538),
            .I(N__29529));
    LocalMux I__6899 (
            .O(N__29535),
            .I(\eeprom.eeprom_counter_11 ));
    Odrv4 I__6898 (
            .O(N__29532),
            .I(\eeprom.eeprom_counter_11 ));
    Odrv4 I__6897 (
            .O(N__29529),
            .I(\eeprom.eeprom_counter_11 ));
    CascadeMux I__6896 (
            .O(N__29522),
            .I(N__29519));
    InMux I__6895 (
            .O(N__29519),
            .I(N__29516));
    LocalMux I__6894 (
            .O(N__29516),
            .I(N__29513));
    Span4Mux_h I__6893 (
            .O(N__29513),
            .I(N__29510));
    Odrv4 I__6892 (
            .O(N__29510),
            .I(\eeprom.n22_adj_266 ));
    CascadeMux I__6891 (
            .O(N__29507),
            .I(N__29504));
    InMux I__6890 (
            .O(N__29504),
            .I(N__29500));
    InMux I__6889 (
            .O(N__29503),
            .I(N__29497));
    LocalMux I__6888 (
            .O(N__29500),
            .I(N__29491));
    LocalMux I__6887 (
            .O(N__29497),
            .I(N__29491));
    InMux I__6886 (
            .O(N__29496),
            .I(N__29488));
    Span4Mux_h I__6885 (
            .O(N__29491),
            .I(N__29485));
    LocalMux I__6884 (
            .O(N__29488),
            .I(\eeprom.eeprom_counter_25 ));
    Odrv4 I__6883 (
            .O(N__29485),
            .I(\eeprom.eeprom_counter_25 ));
    CascadeMux I__6882 (
            .O(N__29480),
            .I(N__29477));
    InMux I__6881 (
            .O(N__29477),
            .I(N__29474));
    LocalMux I__6880 (
            .O(N__29474),
            .I(N__29471));
    Span4Mux_v I__6879 (
            .O(N__29471),
            .I(N__29468));
    Odrv4 I__6878 (
            .O(N__29468),
            .I(\eeprom.n8 ));
    InMux I__6877 (
            .O(N__29465),
            .I(N__29462));
    LocalMux I__6876 (
            .O(N__29462),
            .I(\eeprom.n25_adj_271 ));
    InMux I__6875 (
            .O(N__29459),
            .I(N__29454));
    InMux I__6874 (
            .O(N__29458),
            .I(N__29451));
    InMux I__6873 (
            .O(N__29457),
            .I(N__29448));
    LocalMux I__6872 (
            .O(N__29454),
            .I(N__29445));
    LocalMux I__6871 (
            .O(N__29451),
            .I(N__29442));
    LocalMux I__6870 (
            .O(N__29448),
            .I(N__29439));
    Span4Mux_v I__6869 (
            .O(N__29445),
            .I(N__29436));
    Span4Mux_v I__6868 (
            .O(N__29442),
            .I(N__29431));
    Span4Mux_h I__6867 (
            .O(N__29439),
            .I(N__29431));
    Sp12to4 I__6866 (
            .O(N__29436),
            .I(N__29428));
    Span4Mux_h I__6865 (
            .O(N__29431),
            .I(N__29425));
    Span12Mux_h I__6864 (
            .O(N__29428),
            .I(N__29422));
    Span4Mux_h I__6863 (
            .O(N__29425),
            .I(N__29419));
    Odrv12 I__6862 (
            .O(N__29422),
            .I(\eeprom.n3519 ));
    Odrv4 I__6861 (
            .O(N__29419),
            .I(\eeprom.n3519 ));
    InMux I__6860 (
            .O(N__29414),
            .I(N__29411));
    LocalMux I__6859 (
            .O(N__29411),
            .I(\eeprom.n27_adj_281 ));
    InMux I__6858 (
            .O(N__29408),
            .I(N__29405));
    LocalMux I__6857 (
            .O(N__29405),
            .I(N__29401));
    InMux I__6856 (
            .O(N__29404),
            .I(N__29398));
    Span4Mux_h I__6855 (
            .O(N__29401),
            .I(N__29395));
    LocalMux I__6854 (
            .O(N__29398),
            .I(N__29391));
    Span4Mux_v I__6853 (
            .O(N__29395),
            .I(N__29387));
    InMux I__6852 (
            .O(N__29394),
            .I(N__29384));
    Span4Mux_h I__6851 (
            .O(N__29391),
            .I(N__29381));
    InMux I__6850 (
            .O(N__29390),
            .I(N__29378));
    Odrv4 I__6849 (
            .O(N__29387),
            .I(\eeprom.eeprom_counter_6 ));
    LocalMux I__6848 (
            .O(N__29384),
            .I(\eeprom.eeprom_counter_6 ));
    Odrv4 I__6847 (
            .O(N__29381),
            .I(\eeprom.eeprom_counter_6 ));
    LocalMux I__6846 (
            .O(N__29378),
            .I(\eeprom.eeprom_counter_6 ));
    CascadeMux I__6845 (
            .O(N__29369),
            .I(N__29366));
    InMux I__6844 (
            .O(N__29366),
            .I(N__29363));
    LocalMux I__6843 (
            .O(N__29363),
            .I(N__29360));
    Span4Mux_h I__6842 (
            .O(N__29360),
            .I(N__29357));
    Span4Mux_h I__6841 (
            .O(N__29357),
            .I(N__29354));
    Span4Mux_v I__6840 (
            .O(N__29354),
            .I(N__29351));
    Odrv4 I__6839 (
            .O(N__29351),
            .I(\eeprom.n3719 ));
    InMux I__6838 (
            .O(N__29348),
            .I(N__29344));
    InMux I__6837 (
            .O(N__29347),
            .I(N__29341));
    LocalMux I__6836 (
            .O(N__29344),
            .I(N__29337));
    LocalMux I__6835 (
            .O(N__29341),
            .I(N__29334));
    InMux I__6834 (
            .O(N__29340),
            .I(N__29331));
    Span4Mux_v I__6833 (
            .O(N__29337),
            .I(N__29328));
    Span4Mux_h I__6832 (
            .O(N__29334),
            .I(N__29325));
    LocalMux I__6831 (
            .O(N__29331),
            .I(\eeprom.eeprom_counter_19 ));
    Odrv4 I__6830 (
            .O(N__29328),
            .I(\eeprom.eeprom_counter_19 ));
    Odrv4 I__6829 (
            .O(N__29325),
            .I(\eeprom.eeprom_counter_19 ));
    InMux I__6828 (
            .O(N__29318),
            .I(N__29315));
    LocalMux I__6827 (
            .O(N__29315),
            .I(\eeprom.n14_adj_297 ));
    InMux I__6826 (
            .O(N__29312),
            .I(N__29308));
    InMux I__6825 (
            .O(N__29311),
            .I(N__29305));
    LocalMux I__6824 (
            .O(N__29308),
            .I(N__29299));
    LocalMux I__6823 (
            .O(N__29305),
            .I(N__29299));
    InMux I__6822 (
            .O(N__29304),
            .I(N__29296));
    Odrv4 I__6821 (
            .O(N__29299),
            .I(\eeprom.eeprom_counter_26 ));
    LocalMux I__6820 (
            .O(N__29296),
            .I(\eeprom.eeprom_counter_26 ));
    InMux I__6819 (
            .O(N__29291),
            .I(N__29288));
    LocalMux I__6818 (
            .O(N__29288),
            .I(N__29284));
    InMux I__6817 (
            .O(N__29287),
            .I(N__29281));
    Span4Mux_v I__6816 (
            .O(N__29284),
            .I(N__29276));
    LocalMux I__6815 (
            .O(N__29281),
            .I(N__29276));
    Odrv4 I__6814 (
            .O(N__29276),
            .I(\eeprom.n7_adj_309 ));
    CascadeMux I__6813 (
            .O(N__29273),
            .I(N__29269));
    InMux I__6812 (
            .O(N__29272),
            .I(N__29266));
    InMux I__6811 (
            .O(N__29269),
            .I(N__29263));
    LocalMux I__6810 (
            .O(N__29266),
            .I(N__29260));
    LocalMux I__6809 (
            .O(N__29263),
            .I(N__29257));
    Odrv4 I__6808 (
            .O(N__29260),
            .I(\eeprom.n1140 ));
    Odrv4 I__6807 (
            .O(N__29257),
            .I(\eeprom.n1140 ));
    InMux I__6806 (
            .O(N__29252),
            .I(N__29248));
    InMux I__6805 (
            .O(N__29251),
            .I(N__29245));
    LocalMux I__6804 (
            .O(N__29248),
            .I(N__29241));
    LocalMux I__6803 (
            .O(N__29245),
            .I(N__29238));
    InMux I__6802 (
            .O(N__29244),
            .I(N__29235));
    Span4Mux_h I__6801 (
            .O(N__29241),
            .I(N__29232));
    Span4Mux_h I__6800 (
            .O(N__29238),
            .I(N__29229));
    LocalMux I__6799 (
            .O(N__29235),
            .I(\eeprom.eeprom_counter_8 ));
    Odrv4 I__6798 (
            .O(N__29232),
            .I(\eeprom.eeprom_counter_8 ));
    Odrv4 I__6797 (
            .O(N__29229),
            .I(\eeprom.eeprom_counter_8 ));
    CascadeMux I__6796 (
            .O(N__29222),
            .I(N__29219));
    InMux I__6795 (
            .O(N__29219),
            .I(N__29216));
    LocalMux I__6794 (
            .O(N__29216),
            .I(\eeprom.n25_adj_272 ));
    InMux I__6793 (
            .O(N__29213),
            .I(N__29200));
    InMux I__6792 (
            .O(N__29212),
            .I(N__29187));
    InMux I__6791 (
            .O(N__29211),
            .I(N__29187));
    InMux I__6790 (
            .O(N__29210),
            .I(N__29187));
    InMux I__6789 (
            .O(N__29209),
            .I(N__29187));
    InMux I__6788 (
            .O(N__29208),
            .I(N__29187));
    InMux I__6787 (
            .O(N__29207),
            .I(N__29181));
    InMux I__6786 (
            .O(N__29206),
            .I(N__29165));
    InMux I__6785 (
            .O(N__29205),
            .I(N__29162));
    InMux I__6784 (
            .O(N__29204),
            .I(N__29159));
    InMux I__6783 (
            .O(N__29203),
            .I(N__29156));
    LocalMux I__6782 (
            .O(N__29200),
            .I(N__29153));
    InMux I__6781 (
            .O(N__29199),
            .I(N__29150));
    InMux I__6780 (
            .O(N__29198),
            .I(N__29147));
    LocalMux I__6779 (
            .O(N__29187),
            .I(N__29144));
    InMux I__6778 (
            .O(N__29186),
            .I(N__29141));
    InMux I__6777 (
            .O(N__29185),
            .I(N__29138));
    CascadeMux I__6776 (
            .O(N__29184),
            .I(N__29134));
    LocalMux I__6775 (
            .O(N__29181),
            .I(N__29131));
    InMux I__6774 (
            .O(N__29180),
            .I(N__29124));
    InMux I__6773 (
            .O(N__29179),
            .I(N__29124));
    InMux I__6772 (
            .O(N__29178),
            .I(N__29124));
    InMux I__6771 (
            .O(N__29177),
            .I(N__29117));
    InMux I__6770 (
            .O(N__29176),
            .I(N__29117));
    InMux I__6769 (
            .O(N__29175),
            .I(N__29117));
    InMux I__6768 (
            .O(N__29174),
            .I(N__29112));
    InMux I__6767 (
            .O(N__29173),
            .I(N__29112));
    InMux I__6766 (
            .O(N__29172),
            .I(N__29105));
    InMux I__6765 (
            .O(N__29171),
            .I(N__29105));
    InMux I__6764 (
            .O(N__29170),
            .I(N__29105));
    InMux I__6763 (
            .O(N__29169),
            .I(N__29102));
    InMux I__6762 (
            .O(N__29168),
            .I(N__29099));
    LocalMux I__6761 (
            .O(N__29165),
            .I(N__29091));
    LocalMux I__6760 (
            .O(N__29162),
            .I(N__29087));
    LocalMux I__6759 (
            .O(N__29159),
            .I(N__29084));
    LocalMux I__6758 (
            .O(N__29156),
            .I(N__29081));
    Span4Mux_v I__6757 (
            .O(N__29153),
            .I(N__29072));
    LocalMux I__6756 (
            .O(N__29150),
            .I(N__29072));
    LocalMux I__6755 (
            .O(N__29147),
            .I(N__29072));
    Span4Mux_h I__6754 (
            .O(N__29144),
            .I(N__29072));
    LocalMux I__6753 (
            .O(N__29141),
            .I(N__29069));
    LocalMux I__6752 (
            .O(N__29138),
            .I(N__29066));
    InMux I__6751 (
            .O(N__29137),
            .I(N__29061));
    InMux I__6750 (
            .O(N__29134),
            .I(N__29061));
    Span4Mux_v I__6749 (
            .O(N__29131),
            .I(N__29054));
    LocalMux I__6748 (
            .O(N__29124),
            .I(N__29054));
    LocalMux I__6747 (
            .O(N__29117),
            .I(N__29054));
    LocalMux I__6746 (
            .O(N__29112),
            .I(N__29049));
    LocalMux I__6745 (
            .O(N__29105),
            .I(N__29049));
    LocalMux I__6744 (
            .O(N__29102),
            .I(N__29044));
    LocalMux I__6743 (
            .O(N__29099),
            .I(N__29044));
    InMux I__6742 (
            .O(N__29098),
            .I(N__29037));
    InMux I__6741 (
            .O(N__29097),
            .I(N__29037));
    InMux I__6740 (
            .O(N__29096),
            .I(N__29037));
    InMux I__6739 (
            .O(N__29095),
            .I(N__29034));
    InMux I__6738 (
            .O(N__29094),
            .I(N__29031));
    Span12Mux_h I__6737 (
            .O(N__29091),
            .I(N__29028));
    InMux I__6736 (
            .O(N__29090),
            .I(N__29025));
    Span4Mux_v I__6735 (
            .O(N__29087),
            .I(N__29010));
    Span4Mux_h I__6734 (
            .O(N__29084),
            .I(N__29010));
    Span4Mux_v I__6733 (
            .O(N__29081),
            .I(N__29010));
    Span4Mux_v I__6732 (
            .O(N__29072),
            .I(N__29010));
    Span4Mux_v I__6731 (
            .O(N__29069),
            .I(N__29010));
    Span4Mux_v I__6730 (
            .O(N__29066),
            .I(N__29010));
    LocalMux I__6729 (
            .O(N__29061),
            .I(N__29010));
    Span4Mux_h I__6728 (
            .O(N__29054),
            .I(N__29001));
    Span4Mux_v I__6727 (
            .O(N__29049),
            .I(N__29001));
    Span4Mux_h I__6726 (
            .O(N__29044),
            .I(N__29001));
    LocalMux I__6725 (
            .O(N__29037),
            .I(N__29001));
    LocalMux I__6724 (
            .O(N__29034),
            .I(N__28998));
    LocalMux I__6723 (
            .O(N__29031),
            .I(\eeprom.eeprom_counter_31 ));
    Odrv12 I__6722 (
            .O(N__29028),
            .I(\eeprom.eeprom_counter_31 ));
    LocalMux I__6721 (
            .O(N__29025),
            .I(\eeprom.eeprom_counter_31 ));
    Odrv4 I__6720 (
            .O(N__29010),
            .I(\eeprom.eeprom_counter_31 ));
    Odrv4 I__6719 (
            .O(N__29001),
            .I(\eeprom.eeprom_counter_31 ));
    Odrv4 I__6718 (
            .O(N__28998),
            .I(\eeprom.eeprom_counter_31 ));
    CascadeMux I__6717 (
            .O(N__28985),
            .I(N__28982));
    InMux I__6716 (
            .O(N__28982),
            .I(N__28977));
    InMux I__6715 (
            .O(N__28981),
            .I(N__28974));
    InMux I__6714 (
            .O(N__28980),
            .I(N__28971));
    LocalMux I__6713 (
            .O(N__28977),
            .I(N__28968));
    LocalMux I__6712 (
            .O(N__28974),
            .I(N__28962));
    LocalMux I__6711 (
            .O(N__28971),
            .I(N__28962));
    Span4Mux_v I__6710 (
            .O(N__28968),
            .I(N__28959));
    InMux I__6709 (
            .O(N__28967),
            .I(N__28956));
    Span4Mux_v I__6708 (
            .O(N__28962),
            .I(N__28953));
    Odrv4 I__6707 (
            .O(N__28959),
            .I(\eeprom.n2_adj_307 ));
    LocalMux I__6706 (
            .O(N__28956),
            .I(\eeprom.n2_adj_307 ));
    Odrv4 I__6705 (
            .O(N__28953),
            .I(\eeprom.n2_adj_307 ));
    InMux I__6704 (
            .O(N__28946),
            .I(N__28943));
    LocalMux I__6703 (
            .O(N__28943),
            .I(N__28940));
    Odrv12 I__6702 (
            .O(N__28940),
            .I(\eeprom.n1135 ));
    CascadeMux I__6701 (
            .O(N__28937),
            .I(N__28916));
    CascadeMux I__6700 (
            .O(N__28936),
            .I(N__28912));
    CascadeMux I__6699 (
            .O(N__28935),
            .I(N__28909));
    CascadeMux I__6698 (
            .O(N__28934),
            .I(N__28905));
    CascadeMux I__6697 (
            .O(N__28933),
            .I(N__28901));
    CascadeMux I__6696 (
            .O(N__28932),
            .I(N__28898));
    CascadeMux I__6695 (
            .O(N__28931),
            .I(N__28893));
    CascadeMux I__6694 (
            .O(N__28930),
            .I(N__28889));
    CascadeMux I__6693 (
            .O(N__28929),
            .I(N__28886));
    CascadeMux I__6692 (
            .O(N__28928),
            .I(N__28879));
    CascadeMux I__6691 (
            .O(N__28927),
            .I(N__28870));
    CascadeMux I__6690 (
            .O(N__28926),
            .I(N__28867));
    CascadeMux I__6689 (
            .O(N__28925),
            .I(N__28864));
    CascadeMux I__6688 (
            .O(N__28924),
            .I(N__28861));
    CascadeMux I__6687 (
            .O(N__28923),
            .I(N__28858));
    CascadeMux I__6686 (
            .O(N__28922),
            .I(N__28855));
    CascadeMux I__6685 (
            .O(N__28921),
            .I(N__28852));
    CascadeMux I__6684 (
            .O(N__28920),
            .I(N__28849));
    CascadeMux I__6683 (
            .O(N__28919),
            .I(N__28846));
    InMux I__6682 (
            .O(N__28916),
            .I(N__28838));
    InMux I__6681 (
            .O(N__28915),
            .I(N__28833));
    InMux I__6680 (
            .O(N__28912),
            .I(N__28833));
    InMux I__6679 (
            .O(N__28909),
            .I(N__28824));
    InMux I__6678 (
            .O(N__28908),
            .I(N__28824));
    InMux I__6677 (
            .O(N__28905),
            .I(N__28824));
    InMux I__6676 (
            .O(N__28904),
            .I(N__28824));
    InMux I__6675 (
            .O(N__28901),
            .I(N__28815));
    InMux I__6674 (
            .O(N__28898),
            .I(N__28815));
    InMux I__6673 (
            .O(N__28897),
            .I(N__28815));
    InMux I__6672 (
            .O(N__28896),
            .I(N__28815));
    InMux I__6671 (
            .O(N__28893),
            .I(N__28808));
    InMux I__6670 (
            .O(N__28892),
            .I(N__28808));
    InMux I__6669 (
            .O(N__28889),
            .I(N__28808));
    InMux I__6668 (
            .O(N__28886),
            .I(N__28803));
    InMux I__6667 (
            .O(N__28885),
            .I(N__28803));
    InMux I__6666 (
            .O(N__28884),
            .I(N__28792));
    InMux I__6665 (
            .O(N__28883),
            .I(N__28792));
    InMux I__6664 (
            .O(N__28882),
            .I(N__28792));
    InMux I__6663 (
            .O(N__28879),
            .I(N__28792));
    InMux I__6662 (
            .O(N__28878),
            .I(N__28792));
    InMux I__6661 (
            .O(N__28877),
            .I(N__28785));
    InMux I__6660 (
            .O(N__28876),
            .I(N__28785));
    InMux I__6659 (
            .O(N__28875),
            .I(N__28785));
    CascadeMux I__6658 (
            .O(N__28874),
            .I(N__28778));
    CascadeMux I__6657 (
            .O(N__28873),
            .I(N__28774));
    InMux I__6656 (
            .O(N__28870),
            .I(N__28756));
    InMux I__6655 (
            .O(N__28867),
            .I(N__28747));
    InMux I__6654 (
            .O(N__28864),
            .I(N__28747));
    InMux I__6653 (
            .O(N__28861),
            .I(N__28747));
    InMux I__6652 (
            .O(N__28858),
            .I(N__28747));
    InMux I__6651 (
            .O(N__28855),
            .I(N__28738));
    InMux I__6650 (
            .O(N__28852),
            .I(N__28738));
    InMux I__6649 (
            .O(N__28849),
            .I(N__28738));
    InMux I__6648 (
            .O(N__28846),
            .I(N__28738));
    CascadeMux I__6647 (
            .O(N__28845),
            .I(N__28734));
    CascadeMux I__6646 (
            .O(N__28844),
            .I(N__28730));
    CascadeMux I__6645 (
            .O(N__28843),
            .I(N__28726));
    CascadeMux I__6644 (
            .O(N__28842),
            .I(N__28722));
    CascadeMux I__6643 (
            .O(N__28841),
            .I(N__28718));
    LocalMux I__6642 (
            .O(N__28838),
            .I(N__28699));
    LocalMux I__6641 (
            .O(N__28833),
            .I(N__28699));
    LocalMux I__6640 (
            .O(N__28824),
            .I(N__28699));
    LocalMux I__6639 (
            .O(N__28815),
            .I(N__28699));
    LocalMux I__6638 (
            .O(N__28808),
            .I(N__28690));
    LocalMux I__6637 (
            .O(N__28803),
            .I(N__28690));
    LocalMux I__6636 (
            .O(N__28792),
            .I(N__28690));
    LocalMux I__6635 (
            .O(N__28785),
            .I(N__28690));
    InMux I__6634 (
            .O(N__28784),
            .I(N__28685));
    InMux I__6633 (
            .O(N__28783),
            .I(N__28685));
    InMux I__6632 (
            .O(N__28782),
            .I(N__28676));
    InMux I__6631 (
            .O(N__28781),
            .I(N__28676));
    InMux I__6630 (
            .O(N__28778),
            .I(N__28676));
    InMux I__6629 (
            .O(N__28777),
            .I(N__28676));
    InMux I__6628 (
            .O(N__28774),
            .I(N__28669));
    InMux I__6627 (
            .O(N__28773),
            .I(N__28669));
    InMux I__6626 (
            .O(N__28772),
            .I(N__28669));
    InMux I__6625 (
            .O(N__28771),
            .I(N__28660));
    InMux I__6624 (
            .O(N__28770),
            .I(N__28660));
    InMux I__6623 (
            .O(N__28769),
            .I(N__28660));
    InMux I__6622 (
            .O(N__28768),
            .I(N__28660));
    InMux I__6621 (
            .O(N__28767),
            .I(N__28651));
    InMux I__6620 (
            .O(N__28766),
            .I(N__28651));
    InMux I__6619 (
            .O(N__28765),
            .I(N__28651));
    InMux I__6618 (
            .O(N__28764),
            .I(N__28651));
    CascadeMux I__6617 (
            .O(N__28763),
            .I(N__28648));
    CascadeMux I__6616 (
            .O(N__28762),
            .I(N__28645));
    CascadeMux I__6615 (
            .O(N__28761),
            .I(N__28641));
    CascadeMux I__6614 (
            .O(N__28760),
            .I(N__28638));
    CascadeMux I__6613 (
            .O(N__28759),
            .I(N__28635));
    LocalMux I__6612 (
            .O(N__28756),
            .I(N__28625));
    LocalMux I__6611 (
            .O(N__28747),
            .I(N__28625));
    LocalMux I__6610 (
            .O(N__28738),
            .I(N__28625));
    InMux I__6609 (
            .O(N__28737),
            .I(N__28616));
    InMux I__6608 (
            .O(N__28734),
            .I(N__28616));
    InMux I__6607 (
            .O(N__28733),
            .I(N__28616));
    InMux I__6606 (
            .O(N__28730),
            .I(N__28616));
    InMux I__6605 (
            .O(N__28729),
            .I(N__28607));
    InMux I__6604 (
            .O(N__28726),
            .I(N__28607));
    InMux I__6603 (
            .O(N__28725),
            .I(N__28607));
    InMux I__6602 (
            .O(N__28722),
            .I(N__28607));
    InMux I__6601 (
            .O(N__28721),
            .I(N__28604));
    InMux I__6600 (
            .O(N__28718),
            .I(N__28601));
    CascadeMux I__6599 (
            .O(N__28717),
            .I(N__28596));
    CascadeMux I__6598 (
            .O(N__28716),
            .I(N__28590));
    CascadeMux I__6597 (
            .O(N__28715),
            .I(N__28587));
    CascadeMux I__6596 (
            .O(N__28714),
            .I(N__28583));
    CascadeMux I__6595 (
            .O(N__28713),
            .I(N__28580));
    CascadeMux I__6594 (
            .O(N__28712),
            .I(N__28577));
    CascadeMux I__6593 (
            .O(N__28711),
            .I(N__28573));
    CascadeMux I__6592 (
            .O(N__28710),
            .I(N__28570));
    CascadeMux I__6591 (
            .O(N__28709),
            .I(N__28567));
    CascadeMux I__6590 (
            .O(N__28708),
            .I(N__28564));
    Span4Mux_s3_v I__6589 (
            .O(N__28699),
            .I(N__28540));
    Span4Mux_v I__6588 (
            .O(N__28690),
            .I(N__28524));
    LocalMux I__6587 (
            .O(N__28685),
            .I(N__28524));
    LocalMux I__6586 (
            .O(N__28676),
            .I(N__28524));
    LocalMux I__6585 (
            .O(N__28669),
            .I(N__28524));
    LocalMux I__6584 (
            .O(N__28660),
            .I(N__28524));
    LocalMux I__6583 (
            .O(N__28651),
            .I(N__28524));
    InMux I__6582 (
            .O(N__28648),
            .I(N__28517));
    InMux I__6581 (
            .O(N__28645),
            .I(N__28517));
    InMux I__6580 (
            .O(N__28644),
            .I(N__28517));
    InMux I__6579 (
            .O(N__28641),
            .I(N__28506));
    InMux I__6578 (
            .O(N__28638),
            .I(N__28506));
    InMux I__6577 (
            .O(N__28635),
            .I(N__28506));
    InMux I__6576 (
            .O(N__28634),
            .I(N__28506));
    InMux I__6575 (
            .O(N__28633),
            .I(N__28506));
    CascadeMux I__6574 (
            .O(N__28632),
            .I(N__28501));
    Span4Mux_v I__6573 (
            .O(N__28625),
            .I(N__28489));
    LocalMux I__6572 (
            .O(N__28616),
            .I(N__28489));
    LocalMux I__6571 (
            .O(N__28607),
            .I(N__28489));
    LocalMux I__6570 (
            .O(N__28604),
            .I(N__28489));
    LocalMux I__6569 (
            .O(N__28601),
            .I(N__28489));
    InMux I__6568 (
            .O(N__28600),
            .I(N__28480));
    InMux I__6567 (
            .O(N__28599),
            .I(N__28480));
    InMux I__6566 (
            .O(N__28596),
            .I(N__28480));
    InMux I__6565 (
            .O(N__28595),
            .I(N__28480));
    CascadeMux I__6564 (
            .O(N__28594),
            .I(N__28474));
    InMux I__6563 (
            .O(N__28593),
            .I(N__28469));
    InMux I__6562 (
            .O(N__28590),
            .I(N__28469));
    InMux I__6561 (
            .O(N__28587),
            .I(N__28460));
    InMux I__6560 (
            .O(N__28586),
            .I(N__28460));
    InMux I__6559 (
            .O(N__28583),
            .I(N__28460));
    InMux I__6558 (
            .O(N__28580),
            .I(N__28460));
    InMux I__6557 (
            .O(N__28577),
            .I(N__28451));
    InMux I__6556 (
            .O(N__28576),
            .I(N__28451));
    InMux I__6555 (
            .O(N__28573),
            .I(N__28451));
    InMux I__6554 (
            .O(N__28570),
            .I(N__28451));
    InMux I__6553 (
            .O(N__28567),
            .I(N__28446));
    InMux I__6552 (
            .O(N__28564),
            .I(N__28446));
    InMux I__6551 (
            .O(N__28563),
            .I(N__28441));
    InMux I__6550 (
            .O(N__28562),
            .I(N__28441));
    CascadeMux I__6549 (
            .O(N__28561),
            .I(N__28437));
    CascadeMux I__6548 (
            .O(N__28560),
            .I(N__28434));
    CascadeMux I__6547 (
            .O(N__28559),
            .I(N__28430));
    CascadeMux I__6546 (
            .O(N__28558),
            .I(N__28425));
    CascadeMux I__6545 (
            .O(N__28557),
            .I(N__28422));
    CascadeMux I__6544 (
            .O(N__28556),
            .I(N__28419));
    CascadeMux I__6543 (
            .O(N__28555),
            .I(N__28415));
    CascadeMux I__6542 (
            .O(N__28554),
            .I(N__28412));
    CascadeMux I__6541 (
            .O(N__28553),
            .I(N__28408));
    CascadeMux I__6540 (
            .O(N__28552),
            .I(N__28404));
    CascadeMux I__6539 (
            .O(N__28551),
            .I(N__28401));
    CascadeMux I__6538 (
            .O(N__28550),
            .I(N__28397));
    CascadeMux I__6537 (
            .O(N__28549),
            .I(N__28394));
    CascadeMux I__6536 (
            .O(N__28548),
            .I(N__28387));
    CascadeMux I__6535 (
            .O(N__28547),
            .I(N__28383));
    CascadeMux I__6534 (
            .O(N__28546),
            .I(N__28380));
    CascadeMux I__6533 (
            .O(N__28545),
            .I(N__28376));
    CascadeMux I__6532 (
            .O(N__28544),
            .I(N__28372));
    CascadeMux I__6531 (
            .O(N__28543),
            .I(N__28367));
    Span4Mux_v I__6530 (
            .O(N__28540),
            .I(N__28362));
    InMux I__6529 (
            .O(N__28539),
            .I(N__28357));
    InMux I__6528 (
            .O(N__28538),
            .I(N__28357));
    CascadeMux I__6527 (
            .O(N__28537),
            .I(N__28353));
    Span4Mux_v I__6526 (
            .O(N__28524),
            .I(N__28345));
    LocalMux I__6525 (
            .O(N__28517),
            .I(N__28345));
    LocalMux I__6524 (
            .O(N__28506),
            .I(N__28345));
    InMux I__6523 (
            .O(N__28505),
            .I(N__28340));
    InMux I__6522 (
            .O(N__28504),
            .I(N__28340));
    InMux I__6521 (
            .O(N__28501),
            .I(N__28335));
    InMux I__6520 (
            .O(N__28500),
            .I(N__28335));
    Span4Mux_v I__6519 (
            .O(N__28489),
            .I(N__28330));
    LocalMux I__6518 (
            .O(N__28480),
            .I(N__28330));
    InMux I__6517 (
            .O(N__28479),
            .I(N__28325));
    InMux I__6516 (
            .O(N__28478),
            .I(N__28325));
    InMux I__6515 (
            .O(N__28477),
            .I(N__28320));
    InMux I__6514 (
            .O(N__28474),
            .I(N__28320));
    LocalMux I__6513 (
            .O(N__28469),
            .I(N__28311));
    LocalMux I__6512 (
            .O(N__28460),
            .I(N__28311));
    LocalMux I__6511 (
            .O(N__28451),
            .I(N__28311));
    LocalMux I__6510 (
            .O(N__28446),
            .I(N__28306));
    LocalMux I__6509 (
            .O(N__28441),
            .I(N__28306));
    InMux I__6508 (
            .O(N__28440),
            .I(N__28303));
    InMux I__6507 (
            .O(N__28437),
            .I(N__28298));
    InMux I__6506 (
            .O(N__28434),
            .I(N__28298));
    InMux I__6505 (
            .O(N__28433),
            .I(N__28295));
    InMux I__6504 (
            .O(N__28430),
            .I(N__28292));
    InMux I__6503 (
            .O(N__28429),
            .I(N__28278));
    InMux I__6502 (
            .O(N__28428),
            .I(N__28278));
    InMux I__6501 (
            .O(N__28425),
            .I(N__28278));
    InMux I__6500 (
            .O(N__28422),
            .I(N__28278));
    InMux I__6499 (
            .O(N__28419),
            .I(N__28269));
    InMux I__6498 (
            .O(N__28418),
            .I(N__28269));
    InMux I__6497 (
            .O(N__28415),
            .I(N__28269));
    InMux I__6496 (
            .O(N__28412),
            .I(N__28269));
    CascadeMux I__6495 (
            .O(N__28411),
            .I(N__28265));
    InMux I__6494 (
            .O(N__28408),
            .I(N__28261));
    InMux I__6493 (
            .O(N__28407),
            .I(N__28252));
    InMux I__6492 (
            .O(N__28404),
            .I(N__28252));
    InMux I__6491 (
            .O(N__28401),
            .I(N__28252));
    InMux I__6490 (
            .O(N__28400),
            .I(N__28252));
    InMux I__6489 (
            .O(N__28397),
            .I(N__28247));
    InMux I__6488 (
            .O(N__28394),
            .I(N__28247));
    CascadeMux I__6487 (
            .O(N__28393),
            .I(N__28244));
    InMux I__6486 (
            .O(N__28392),
            .I(N__28237));
    InMux I__6485 (
            .O(N__28391),
            .I(N__28237));
    InMux I__6484 (
            .O(N__28390),
            .I(N__28230));
    InMux I__6483 (
            .O(N__28387),
            .I(N__28230));
    InMux I__6482 (
            .O(N__28386),
            .I(N__28230));
    InMux I__6481 (
            .O(N__28383),
            .I(N__28219));
    InMux I__6480 (
            .O(N__28380),
            .I(N__28219));
    InMux I__6479 (
            .O(N__28379),
            .I(N__28219));
    InMux I__6478 (
            .O(N__28376),
            .I(N__28219));
    InMux I__6477 (
            .O(N__28375),
            .I(N__28219));
    InMux I__6476 (
            .O(N__28372),
            .I(N__28216));
    InMux I__6475 (
            .O(N__28371),
            .I(N__28213));
    InMux I__6474 (
            .O(N__28370),
            .I(N__28204));
    InMux I__6473 (
            .O(N__28367),
            .I(N__28204));
    InMux I__6472 (
            .O(N__28366),
            .I(N__28204));
    InMux I__6471 (
            .O(N__28365),
            .I(N__28204));
    Span4Mux_v I__6470 (
            .O(N__28362),
            .I(N__28199));
    LocalMux I__6469 (
            .O(N__28357),
            .I(N__28199));
    InMux I__6468 (
            .O(N__28356),
            .I(N__28194));
    InMux I__6467 (
            .O(N__28353),
            .I(N__28194));
    CascadeMux I__6466 (
            .O(N__28352),
            .I(N__28191));
    Span4Mux_h I__6465 (
            .O(N__28345),
            .I(N__28185));
    LocalMux I__6464 (
            .O(N__28340),
            .I(N__28185));
    LocalMux I__6463 (
            .O(N__28335),
            .I(N__28178));
    Span4Mux_h I__6462 (
            .O(N__28330),
            .I(N__28178));
    LocalMux I__6461 (
            .O(N__28325),
            .I(N__28178));
    LocalMux I__6460 (
            .O(N__28320),
            .I(N__28175));
    InMux I__6459 (
            .O(N__28319),
            .I(N__28170));
    InMux I__6458 (
            .O(N__28318),
            .I(N__28170));
    Span4Mux_s3_v I__6457 (
            .O(N__28311),
            .I(N__28164));
    Span4Mux_s3_v I__6456 (
            .O(N__28306),
            .I(N__28164));
    LocalMux I__6455 (
            .O(N__28303),
            .I(N__28161));
    LocalMux I__6454 (
            .O(N__28298),
            .I(N__28154));
    LocalMux I__6453 (
            .O(N__28295),
            .I(N__28154));
    LocalMux I__6452 (
            .O(N__28292),
            .I(N__28154));
    CascadeMux I__6451 (
            .O(N__28291),
            .I(N__28150));
    CascadeMux I__6450 (
            .O(N__28290),
            .I(N__28146));
    CascadeMux I__6449 (
            .O(N__28289),
            .I(N__28142));
    CascadeMux I__6448 (
            .O(N__28288),
            .I(N__28138));
    CascadeMux I__6447 (
            .O(N__28287),
            .I(N__28135));
    LocalMux I__6446 (
            .O(N__28278),
            .I(N__28129));
    LocalMux I__6445 (
            .O(N__28269),
            .I(N__28129));
    InMux I__6444 (
            .O(N__28268),
            .I(N__28122));
    InMux I__6443 (
            .O(N__28265),
            .I(N__28122));
    InMux I__6442 (
            .O(N__28264),
            .I(N__28122));
    LocalMux I__6441 (
            .O(N__28261),
            .I(N__28115));
    LocalMux I__6440 (
            .O(N__28252),
            .I(N__28115));
    LocalMux I__6439 (
            .O(N__28247),
            .I(N__28115));
    InMux I__6438 (
            .O(N__28244),
            .I(N__28112));
    InMux I__6437 (
            .O(N__28243),
            .I(N__28109));
    InMux I__6436 (
            .O(N__28242),
            .I(N__28106));
    LocalMux I__6435 (
            .O(N__28237),
            .I(N__28090));
    LocalMux I__6434 (
            .O(N__28230),
            .I(N__28090));
    LocalMux I__6433 (
            .O(N__28219),
            .I(N__28090));
    LocalMux I__6432 (
            .O(N__28216),
            .I(N__28090));
    LocalMux I__6431 (
            .O(N__28213),
            .I(N__28090));
    LocalMux I__6430 (
            .O(N__28204),
            .I(N__28090));
    Span4Mux_v I__6429 (
            .O(N__28199),
            .I(N__28085));
    LocalMux I__6428 (
            .O(N__28194),
            .I(N__28085));
    InMux I__6427 (
            .O(N__28191),
            .I(N__28082));
    InMux I__6426 (
            .O(N__28190),
            .I(N__28079));
    Span4Mux_v I__6425 (
            .O(N__28185),
            .I(N__28076));
    Span4Mux_v I__6424 (
            .O(N__28178),
            .I(N__28069));
    Span4Mux_h I__6423 (
            .O(N__28175),
            .I(N__28069));
    LocalMux I__6422 (
            .O(N__28170),
            .I(N__28069));
    InMux I__6421 (
            .O(N__28169),
            .I(N__28066));
    Sp12to4 I__6420 (
            .O(N__28164),
            .I(N__28063));
    Span4Mux_s3_v I__6419 (
            .O(N__28161),
            .I(N__28058));
    Span4Mux_h I__6418 (
            .O(N__28154),
            .I(N__28058));
    InMux I__6417 (
            .O(N__28153),
            .I(N__28055));
    InMux I__6416 (
            .O(N__28150),
            .I(N__28048));
    InMux I__6415 (
            .O(N__28149),
            .I(N__28048));
    InMux I__6414 (
            .O(N__28146),
            .I(N__28048));
    InMux I__6413 (
            .O(N__28145),
            .I(N__28039));
    InMux I__6412 (
            .O(N__28142),
            .I(N__28039));
    InMux I__6411 (
            .O(N__28141),
            .I(N__28039));
    InMux I__6410 (
            .O(N__28138),
            .I(N__28039));
    InMux I__6409 (
            .O(N__28135),
            .I(N__28036));
    InMux I__6408 (
            .O(N__28134),
            .I(N__28033));
    Span4Mux_h I__6407 (
            .O(N__28129),
            .I(N__28026));
    LocalMux I__6406 (
            .O(N__28122),
            .I(N__28026));
    Span4Mux_v I__6405 (
            .O(N__28115),
            .I(N__28021));
    LocalMux I__6404 (
            .O(N__28112),
            .I(N__28021));
    LocalMux I__6403 (
            .O(N__28109),
            .I(N__28016));
    LocalMux I__6402 (
            .O(N__28106),
            .I(N__28016));
    CascadeMux I__6401 (
            .O(N__28105),
            .I(N__28012));
    CascadeMux I__6400 (
            .O(N__28104),
            .I(N__28008));
    CascadeMux I__6399 (
            .O(N__28103),
            .I(N__28004));
    Span12Mux_v I__6398 (
            .O(N__28090),
            .I(N__28000));
    Span4Mux_h I__6397 (
            .O(N__28085),
            .I(N__27993));
    LocalMux I__6396 (
            .O(N__28082),
            .I(N__27993));
    LocalMux I__6395 (
            .O(N__28079),
            .I(N__27993));
    Span4Mux_h I__6394 (
            .O(N__28076),
            .I(N__27988));
    Span4Mux_v I__6393 (
            .O(N__28069),
            .I(N__27988));
    LocalMux I__6392 (
            .O(N__28066),
            .I(N__27985));
    Span12Mux_s11_h I__6391 (
            .O(N__28063),
            .I(N__27970));
    Sp12to4 I__6390 (
            .O(N__28058),
            .I(N__27970));
    LocalMux I__6389 (
            .O(N__28055),
            .I(N__27970));
    LocalMux I__6388 (
            .O(N__28048),
            .I(N__27970));
    LocalMux I__6387 (
            .O(N__28039),
            .I(N__27970));
    LocalMux I__6386 (
            .O(N__28036),
            .I(N__27970));
    LocalMux I__6385 (
            .O(N__28033),
            .I(N__27970));
    InMux I__6384 (
            .O(N__28032),
            .I(N__27965));
    InMux I__6383 (
            .O(N__28031),
            .I(N__27965));
    Span4Mux_v I__6382 (
            .O(N__28026),
            .I(N__27960));
    Span4Mux_v I__6381 (
            .O(N__28021),
            .I(N__27960));
    Span4Mux_v I__6380 (
            .O(N__28016),
            .I(N__27957));
    InMux I__6379 (
            .O(N__28015),
            .I(N__27942));
    InMux I__6378 (
            .O(N__28012),
            .I(N__27942));
    InMux I__6377 (
            .O(N__28011),
            .I(N__27942));
    InMux I__6376 (
            .O(N__28008),
            .I(N__27942));
    InMux I__6375 (
            .O(N__28007),
            .I(N__27942));
    InMux I__6374 (
            .O(N__28004),
            .I(N__27942));
    InMux I__6373 (
            .O(N__28003),
            .I(N__27942));
    Span12Mux_h I__6372 (
            .O(N__28000),
            .I(N__27939));
    Span4Mux_h I__6371 (
            .O(N__27993),
            .I(N__27936));
    Span4Mux_h I__6370 (
            .O(N__27988),
            .I(N__27931));
    Span4Mux_v I__6369 (
            .O(N__27985),
            .I(N__27931));
    Span12Mux_v I__6368 (
            .O(N__27970),
            .I(N__27926));
    LocalMux I__6367 (
            .O(N__27965),
            .I(N__27926));
    Span4Mux_h I__6366 (
            .O(N__27960),
            .I(N__27919));
    Span4Mux_h I__6365 (
            .O(N__27957),
            .I(N__27919));
    LocalMux I__6364 (
            .O(N__27942),
            .I(N__27919));
    Odrv12 I__6363 (
            .O(N__27939),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6362 (
            .O(N__27936),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6361 (
            .O(N__27931),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6360 (
            .O(N__27926),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6359 (
            .O(N__27919),
            .I(CONSTANT_ONE_NET));
    InMux I__6358 (
            .O(N__27908),
            .I(N__27905));
    LocalMux I__6357 (
            .O(N__27905),
            .I(n174));
    CascadeMux I__6356 (
            .O(N__27902),
            .I(N__27899));
    InMux I__6355 (
            .O(N__27899),
            .I(N__27896));
    LocalMux I__6354 (
            .O(N__27896),
            .I(N__27892));
    InMux I__6353 (
            .O(N__27895),
            .I(N__27889));
    Odrv12 I__6352 (
            .O(N__27892),
            .I(rw));
    LocalMux I__6351 (
            .O(N__27889),
            .I(rw));
    InMux I__6350 (
            .O(N__27884),
            .I(N__27881));
    LocalMux I__6349 (
            .O(N__27881),
            .I(N__27876));
    InMux I__6348 (
            .O(N__27880),
            .I(N__27873));
    InMux I__6347 (
            .O(N__27879),
            .I(N__27870));
    Span4Mux_v I__6346 (
            .O(N__27876),
            .I(N__27867));
    LocalMux I__6345 (
            .O(N__27873),
            .I(N__27864));
    LocalMux I__6344 (
            .O(N__27870),
            .I(saved_addr_0));
    Odrv4 I__6343 (
            .O(N__27867),
            .I(saved_addr_0));
    Odrv4 I__6342 (
            .O(N__27864),
            .I(saved_addr_0));
    InMux I__6341 (
            .O(N__27857),
            .I(\eeprom.n4278 ));
    InMux I__6340 (
            .O(N__27854),
            .I(N__27851));
    LocalMux I__6339 (
            .O(N__27851),
            .I(N__27848));
    Odrv4 I__6338 (
            .O(N__27848),
            .I(\eeprom.n1192 ));
    CascadeMux I__6337 (
            .O(N__27845),
            .I(N__27840));
    CascadeMux I__6336 (
            .O(N__27844),
            .I(N__27837));
    InMux I__6335 (
            .O(N__27843),
            .I(N__27834));
    InMux I__6334 (
            .O(N__27840),
            .I(N__27831));
    InMux I__6333 (
            .O(N__27837),
            .I(N__27828));
    LocalMux I__6332 (
            .O(N__27834),
            .I(N__27823));
    LocalMux I__6331 (
            .O(N__27831),
            .I(N__27823));
    LocalMux I__6330 (
            .O(N__27828),
            .I(\eeprom.n1256 ));
    Odrv4 I__6329 (
            .O(N__27823),
            .I(\eeprom.n1256 ));
    CascadeMux I__6328 (
            .O(N__27818),
            .I(\eeprom.n1843_cascade_ ));
    InMux I__6327 (
            .O(N__27815),
            .I(N__27812));
    LocalMux I__6326 (
            .O(N__27812),
            .I(\eeprom.n1195 ));
    CascadeMux I__6325 (
            .O(N__27809),
            .I(N__27805));
    InMux I__6324 (
            .O(N__27808),
            .I(N__27802));
    InMux I__6323 (
            .O(N__27805),
            .I(N__27799));
    LocalMux I__6322 (
            .O(N__27802),
            .I(N__27794));
    LocalMux I__6321 (
            .O(N__27799),
            .I(N__27794));
    Span4Mux_v I__6320 (
            .O(N__27794),
            .I(N__27790));
    InMux I__6319 (
            .O(N__27793),
            .I(N__27787));
    Odrv4 I__6318 (
            .O(N__27790),
            .I(\eeprom.n1915 ));
    LocalMux I__6317 (
            .O(N__27787),
            .I(\eeprom.n1915 ));
    InMux I__6316 (
            .O(N__27782),
            .I(N__27779));
    LocalMux I__6315 (
            .O(N__27779),
            .I(N__27775));
    InMux I__6314 (
            .O(N__27778),
            .I(N__27771));
    Span4Mux_h I__6313 (
            .O(N__27775),
            .I(N__27768));
    InMux I__6312 (
            .O(N__27774),
            .I(N__27765));
    LocalMux I__6311 (
            .O(N__27771),
            .I(\eeprom.eeprom_counter_29 ));
    Odrv4 I__6310 (
            .O(N__27768),
            .I(\eeprom.eeprom_counter_29 ));
    LocalMux I__6309 (
            .O(N__27765),
            .I(\eeprom.eeprom_counter_29 ));
    InMux I__6308 (
            .O(N__27758),
            .I(N__27755));
    LocalMux I__6307 (
            .O(N__27755),
            .I(N__27752));
    Span4Mux_h I__6306 (
            .O(N__27752),
            .I(N__27749));
    Odrv4 I__6305 (
            .O(N__27749),
            .I(\eeprom.n4_adj_310 ));
    CascadeMux I__6304 (
            .O(N__27746),
            .I(N__27743));
    InMux I__6303 (
            .O(N__27743),
            .I(N__27738));
    InMux I__6302 (
            .O(N__27742),
            .I(N__27733));
    InMux I__6301 (
            .O(N__27741),
            .I(N__27733));
    LocalMux I__6300 (
            .O(N__27738),
            .I(\eeprom.n1138 ));
    LocalMux I__6299 (
            .O(N__27733),
            .I(\eeprom.n1138 ));
    CascadeMux I__6298 (
            .O(N__27728),
            .I(\eeprom.n1137_cascade_ ));
    InMux I__6297 (
            .O(N__27725),
            .I(N__27721));
    InMux I__6296 (
            .O(N__27724),
            .I(N__27718));
    LocalMux I__6295 (
            .O(N__27721),
            .I(\eeprom.n4977 ));
    LocalMux I__6294 (
            .O(N__27718),
            .I(\eeprom.n4977 ));
    InMux I__6293 (
            .O(N__27713),
            .I(N__27710));
    LocalMux I__6292 (
            .O(N__27710),
            .I(\eeprom.n4983 ));
    InMux I__6291 (
            .O(N__27707),
            .I(N__27704));
    LocalMux I__6290 (
            .O(N__27704),
            .I(\eeprom.n1197 ));
    CascadeMux I__6289 (
            .O(N__27701),
            .I(N__27697));
    CascadeMux I__6288 (
            .O(N__27700),
            .I(N__27694));
    InMux I__6287 (
            .O(N__27697),
            .I(N__27691));
    InMux I__6286 (
            .O(N__27694),
            .I(N__27688));
    LocalMux I__6285 (
            .O(N__27691),
            .I(N__27685));
    LocalMux I__6284 (
            .O(N__27688),
            .I(N__27682));
    Span4Mux_h I__6283 (
            .O(N__27685),
            .I(N__27678));
    Span4Mux_h I__6282 (
            .O(N__27682),
            .I(N__27675));
    InMux I__6281 (
            .O(N__27681),
            .I(N__27672));
    Odrv4 I__6280 (
            .O(N__27678),
            .I(\eeprom.n1917 ));
    Odrv4 I__6279 (
            .O(N__27675),
            .I(\eeprom.n1917 ));
    LocalMux I__6278 (
            .O(N__27672),
            .I(\eeprom.n1917 ));
    InMux I__6277 (
            .O(N__27665),
            .I(N__27662));
    LocalMux I__6276 (
            .O(N__27662),
            .I(\eeprom.n1194 ));
    CascadeMux I__6275 (
            .O(N__27659),
            .I(N__27656));
    InMux I__6274 (
            .O(N__27656),
            .I(N__27651));
    InMux I__6273 (
            .O(N__27655),
            .I(N__27648));
    InMux I__6272 (
            .O(N__27654),
            .I(N__27645));
    LocalMux I__6271 (
            .O(N__27651),
            .I(\eeprom.n1137 ));
    LocalMux I__6270 (
            .O(N__27648),
            .I(\eeprom.n1137 ));
    LocalMux I__6269 (
            .O(N__27645),
            .I(\eeprom.n1137 ));
    CascadeMux I__6268 (
            .O(N__27638),
            .I(N__27632));
    InMux I__6267 (
            .O(N__27637),
            .I(N__27624));
    InMux I__6266 (
            .O(N__27636),
            .I(N__27624));
    InMux I__6265 (
            .O(N__27635),
            .I(N__27624));
    InMux I__6264 (
            .O(N__27632),
            .I(N__27619));
    InMux I__6263 (
            .O(N__27631),
            .I(N__27619));
    LocalMux I__6262 (
            .O(N__27624),
            .I(\eeprom.n1843 ));
    LocalMux I__6261 (
            .O(N__27619),
            .I(\eeprom.n1843 ));
    CascadeMux I__6260 (
            .O(N__27614),
            .I(N__27610));
    InMux I__6259 (
            .O(N__27613),
            .I(N__27607));
    InMux I__6258 (
            .O(N__27610),
            .I(N__27604));
    LocalMux I__6257 (
            .O(N__27607),
            .I(N__27601));
    LocalMux I__6256 (
            .O(N__27604),
            .I(N__27598));
    Span4Mux_v I__6255 (
            .O(N__27601),
            .I(N__27594));
    Span4Mux_h I__6254 (
            .O(N__27598),
            .I(N__27591));
    InMux I__6253 (
            .O(N__27597),
            .I(N__27588));
    Odrv4 I__6252 (
            .O(N__27594),
            .I(\eeprom.n1914 ));
    Odrv4 I__6251 (
            .O(N__27591),
            .I(\eeprom.n1914 ));
    LocalMux I__6250 (
            .O(N__27588),
            .I(\eeprom.n1914 ));
    InMux I__6249 (
            .O(N__27581),
            .I(N__27577));
    InMux I__6248 (
            .O(N__27580),
            .I(N__27574));
    LocalMux I__6247 (
            .O(N__27577),
            .I(N__27570));
    LocalMux I__6246 (
            .O(N__27574),
            .I(N__27567));
    InMux I__6245 (
            .O(N__27573),
            .I(N__27564));
    Span4Mux_h I__6244 (
            .O(N__27570),
            .I(N__27561));
    Span4Mux_h I__6243 (
            .O(N__27567),
            .I(N__27558));
    LocalMux I__6242 (
            .O(N__27564),
            .I(\eeprom.eeprom_counter_14 ));
    Odrv4 I__6241 (
            .O(N__27561),
            .I(\eeprom.eeprom_counter_14 ));
    Odrv4 I__6240 (
            .O(N__27558),
            .I(\eeprom.eeprom_counter_14 ));
    CascadeMux I__6239 (
            .O(N__27551),
            .I(N__27548));
    InMux I__6238 (
            .O(N__27548),
            .I(N__27545));
    LocalMux I__6237 (
            .O(N__27545),
            .I(\eeprom.n19 ));
    InMux I__6236 (
            .O(N__27542),
            .I(N__27535));
    InMux I__6235 (
            .O(N__27541),
            .I(N__27528));
    InMux I__6234 (
            .O(N__27540),
            .I(N__27528));
    InMux I__6233 (
            .O(N__27539),
            .I(N__27528));
    CascadeMux I__6232 (
            .O(N__27538),
            .I(N__27517));
    LocalMux I__6231 (
            .O(N__27535),
            .I(N__27508));
    LocalMux I__6230 (
            .O(N__27528),
            .I(N__27508));
    InMux I__6229 (
            .O(N__27527),
            .I(N__27503));
    InMux I__6228 (
            .O(N__27526),
            .I(N__27503));
    InMux I__6227 (
            .O(N__27525),
            .I(N__27496));
    InMux I__6226 (
            .O(N__27524),
            .I(N__27496));
    InMux I__6225 (
            .O(N__27523),
            .I(N__27496));
    CascadeMux I__6224 (
            .O(N__27522),
            .I(N__27490));
    InMux I__6223 (
            .O(N__27521),
            .I(N__27485));
    InMux I__6222 (
            .O(N__27520),
            .I(N__27485));
    InMux I__6221 (
            .O(N__27517),
            .I(N__27482));
    InMux I__6220 (
            .O(N__27516),
            .I(N__27475));
    InMux I__6219 (
            .O(N__27515),
            .I(N__27475));
    InMux I__6218 (
            .O(N__27514),
            .I(N__27475));
    InMux I__6217 (
            .O(N__27513),
            .I(N__27472));
    Span4Mux_v I__6216 (
            .O(N__27508),
            .I(N__27465));
    LocalMux I__6215 (
            .O(N__27503),
            .I(N__27465));
    LocalMux I__6214 (
            .O(N__27496),
            .I(N__27465));
    InMux I__6213 (
            .O(N__27495),
            .I(N__27456));
    InMux I__6212 (
            .O(N__27494),
            .I(N__27456));
    InMux I__6211 (
            .O(N__27493),
            .I(N__27456));
    InMux I__6210 (
            .O(N__27490),
            .I(N__27456));
    LocalMux I__6209 (
            .O(N__27485),
            .I(state_1));
    LocalMux I__6208 (
            .O(N__27482),
            .I(state_1));
    LocalMux I__6207 (
            .O(N__27475),
            .I(state_1));
    LocalMux I__6206 (
            .O(N__27472),
            .I(state_1));
    Odrv4 I__6205 (
            .O(N__27465),
            .I(state_1));
    LocalMux I__6204 (
            .O(N__27456),
            .I(state_1));
    InMux I__6203 (
            .O(N__27443),
            .I(N__27440));
    LocalMux I__6202 (
            .O(N__27440),
            .I(n3581));
    InMux I__6201 (
            .O(N__27437),
            .I(N__27433));
    InMux I__6200 (
            .O(N__27436),
            .I(N__27430));
    LocalMux I__6199 (
            .O(N__27433),
            .I(\eeprom.i2c.n407 ));
    LocalMux I__6198 (
            .O(N__27430),
            .I(\eeprom.i2c.n407 ));
    InMux I__6197 (
            .O(N__27425),
            .I(N__27420));
    CascadeMux I__6196 (
            .O(N__27424),
            .I(N__27415));
    InMux I__6195 (
            .O(N__27423),
            .I(N__27412));
    LocalMux I__6194 (
            .O(N__27420),
            .I(N__27397));
    InMux I__6193 (
            .O(N__27419),
            .I(N__27390));
    InMux I__6192 (
            .O(N__27418),
            .I(N__27390));
    InMux I__6191 (
            .O(N__27415),
            .I(N__27390));
    LocalMux I__6190 (
            .O(N__27412),
            .I(N__27387));
    InMux I__6189 (
            .O(N__27411),
            .I(N__27382));
    InMux I__6188 (
            .O(N__27410),
            .I(N__27375));
    InMux I__6187 (
            .O(N__27409),
            .I(N__27375));
    InMux I__6186 (
            .O(N__27408),
            .I(N__27375));
    InMux I__6185 (
            .O(N__27407),
            .I(N__27370));
    InMux I__6184 (
            .O(N__27406),
            .I(N__27370));
    InMux I__6183 (
            .O(N__27405),
            .I(N__27364));
    InMux I__6182 (
            .O(N__27404),
            .I(N__27353));
    InMux I__6181 (
            .O(N__27403),
            .I(N__27353));
    InMux I__6180 (
            .O(N__27402),
            .I(N__27353));
    InMux I__6179 (
            .O(N__27401),
            .I(N__27353));
    InMux I__6178 (
            .O(N__27400),
            .I(N__27353));
    Span4Mux_v I__6177 (
            .O(N__27397),
            .I(N__27348));
    LocalMux I__6176 (
            .O(N__27390),
            .I(N__27348));
    Span4Mux_h I__6175 (
            .O(N__27387),
            .I(N__27345));
    InMux I__6174 (
            .O(N__27386),
            .I(N__27340));
    InMux I__6173 (
            .O(N__27385),
            .I(N__27340));
    LocalMux I__6172 (
            .O(N__27382),
            .I(N__27333));
    LocalMux I__6171 (
            .O(N__27375),
            .I(N__27333));
    LocalMux I__6170 (
            .O(N__27370),
            .I(N__27333));
    InMux I__6169 (
            .O(N__27369),
            .I(N__27326));
    InMux I__6168 (
            .O(N__27368),
            .I(N__27326));
    InMux I__6167 (
            .O(N__27367),
            .I(N__27326));
    LocalMux I__6166 (
            .O(N__27364),
            .I(state_0));
    LocalMux I__6165 (
            .O(N__27353),
            .I(state_0));
    Odrv4 I__6164 (
            .O(N__27348),
            .I(state_0));
    Odrv4 I__6163 (
            .O(N__27345),
            .I(state_0));
    LocalMux I__6162 (
            .O(N__27340),
            .I(state_0));
    Odrv4 I__6161 (
            .O(N__27333),
            .I(state_0));
    LocalMux I__6160 (
            .O(N__27326),
            .I(state_0));
    IoInMux I__6159 (
            .O(N__27311),
            .I(N__27308));
    LocalMux I__6158 (
            .O(N__27308),
            .I(N__27305));
    Span12Mux_s4_h I__6157 (
            .O(N__27305),
            .I(N__27302));
    Span12Mux_v I__6156 (
            .O(N__27302),
            .I(N__27298));
    InMux I__6155 (
            .O(N__27301),
            .I(N__27295));
    Odrv12 I__6154 (
            .O(N__27298),
            .I(sda_enable));
    LocalMux I__6153 (
            .O(N__27295),
            .I(sda_enable));
    CEMux I__6152 (
            .O(N__27290),
            .I(N__27287));
    LocalMux I__6151 (
            .O(N__27287),
            .I(N__27284));
    Span4Mux_h I__6150 (
            .O(N__27284),
            .I(N__27281));
    Odrv4 I__6149 (
            .O(N__27281),
            .I(\eeprom.i2c.n524 ));
    SRMux I__6148 (
            .O(N__27278),
            .I(N__27275));
    LocalMux I__6147 (
            .O(N__27275),
            .I(N__27272));
    Odrv4 I__6146 (
            .O(N__27272),
            .I(\eeprom.i2c.n1901 ));
    CascadeMux I__6145 (
            .O(N__27269),
            .I(N__27265));
    InMux I__6144 (
            .O(N__27268),
            .I(N__27262));
    InMux I__6143 (
            .O(N__27265),
            .I(N__27259));
    LocalMux I__6142 (
            .O(N__27262),
            .I(\eeprom.n892 ));
    LocalMux I__6141 (
            .O(N__27259),
            .I(\eeprom.n892 ));
    CascadeMux I__6140 (
            .O(N__27254),
            .I(N__27251));
    InMux I__6139 (
            .O(N__27251),
            .I(N__27248));
    LocalMux I__6138 (
            .O(N__27248),
            .I(\eeprom.n1198 ));
    InMux I__6137 (
            .O(N__27245),
            .I(bfn_28_21_0_));
    InMux I__6136 (
            .O(N__27242),
            .I(\eeprom.n4273 ));
    CascadeMux I__6135 (
            .O(N__27239),
            .I(N__27236));
    InMux I__6134 (
            .O(N__27236),
            .I(N__27233));
    LocalMux I__6133 (
            .O(N__27233),
            .I(\eeprom.n1139 ));
    InMux I__6132 (
            .O(N__27230),
            .I(N__27227));
    LocalMux I__6131 (
            .O(N__27227),
            .I(\eeprom.n1196 ));
    InMux I__6130 (
            .O(N__27224),
            .I(\eeprom.n4274 ));
    InMux I__6129 (
            .O(N__27221),
            .I(\eeprom.n4275 ));
    InMux I__6128 (
            .O(N__27218),
            .I(\eeprom.n4276 ));
    InMux I__6127 (
            .O(N__27215),
            .I(N__27212));
    LocalMux I__6126 (
            .O(N__27212),
            .I(\eeprom.n5327 ));
    CascadeMux I__6125 (
            .O(N__27209),
            .I(N__27205));
    InMux I__6124 (
            .O(N__27208),
            .I(N__27202));
    InMux I__6123 (
            .O(N__27205),
            .I(N__27199));
    LocalMux I__6122 (
            .O(N__27202),
            .I(\eeprom.n5328 ));
    LocalMux I__6121 (
            .O(N__27199),
            .I(\eeprom.n5328 ));
    InMux I__6120 (
            .O(N__27194),
            .I(\eeprom.n4277 ));
    InMux I__6119 (
            .O(N__27191),
            .I(N__27188));
    LocalMux I__6118 (
            .O(N__27188),
            .I(n11_adj_359));
    InMux I__6117 (
            .O(N__27185),
            .I(N__27182));
    LocalMux I__6116 (
            .O(N__27182),
            .I(n5458));
    CascadeMux I__6115 (
            .O(N__27179),
            .I(n6_adj_365_cascade_));
    InMux I__6114 (
            .O(N__27176),
            .I(N__27171));
    InMux I__6113 (
            .O(N__27175),
            .I(N__27166));
    InMux I__6112 (
            .O(N__27174),
            .I(N__27166));
    LocalMux I__6111 (
            .O(N__27171),
            .I(n471));
    LocalMux I__6110 (
            .O(N__27166),
            .I(n471));
    CascadeMux I__6109 (
            .O(N__27161),
            .I(N__27154));
    CascadeMux I__6108 (
            .O(N__27160),
            .I(N__27145));
    CascadeMux I__6107 (
            .O(N__27159),
            .I(N__27139));
    InMux I__6106 (
            .O(N__27158),
            .I(N__27133));
    InMux I__6105 (
            .O(N__27157),
            .I(N__27133));
    InMux I__6104 (
            .O(N__27154),
            .I(N__27126));
    InMux I__6103 (
            .O(N__27153),
            .I(N__27119));
    InMux I__6102 (
            .O(N__27152),
            .I(N__27119));
    InMux I__6101 (
            .O(N__27151),
            .I(N__27119));
    InMux I__6100 (
            .O(N__27150),
            .I(N__27112));
    InMux I__6099 (
            .O(N__27149),
            .I(N__27112));
    InMux I__6098 (
            .O(N__27148),
            .I(N__27112));
    InMux I__6097 (
            .O(N__27145),
            .I(N__27107));
    InMux I__6096 (
            .O(N__27144),
            .I(N__27107));
    InMux I__6095 (
            .O(N__27143),
            .I(N__27104));
    InMux I__6094 (
            .O(N__27142),
            .I(N__27101));
    InMux I__6093 (
            .O(N__27139),
            .I(N__27096));
    InMux I__6092 (
            .O(N__27138),
            .I(N__27096));
    LocalMux I__6091 (
            .O(N__27133),
            .I(N__27093));
    InMux I__6090 (
            .O(N__27132),
            .I(N__27084));
    InMux I__6089 (
            .O(N__27131),
            .I(N__27084));
    InMux I__6088 (
            .O(N__27130),
            .I(N__27084));
    InMux I__6087 (
            .O(N__27129),
            .I(N__27084));
    LocalMux I__6086 (
            .O(N__27126),
            .I(state_3));
    LocalMux I__6085 (
            .O(N__27119),
            .I(state_3));
    LocalMux I__6084 (
            .O(N__27112),
            .I(state_3));
    LocalMux I__6083 (
            .O(N__27107),
            .I(state_3));
    LocalMux I__6082 (
            .O(N__27104),
            .I(state_3));
    LocalMux I__6081 (
            .O(N__27101),
            .I(state_3));
    LocalMux I__6080 (
            .O(N__27096),
            .I(state_3));
    Odrv4 I__6079 (
            .O(N__27093),
            .I(state_3));
    LocalMux I__6078 (
            .O(N__27084),
            .I(state_3));
    InMux I__6077 (
            .O(N__27065),
            .I(N__27062));
    LocalMux I__6076 (
            .O(N__27062),
            .I(n3587));
    CascadeMux I__6075 (
            .O(N__27059),
            .I(n3587_cascade_));
    InMux I__6074 (
            .O(N__27056),
            .I(N__27052));
    InMux I__6073 (
            .O(N__27055),
            .I(N__27049));
    LocalMux I__6072 (
            .O(N__27052),
            .I(n10));
    LocalMux I__6071 (
            .O(N__27049),
            .I(n10));
    InMux I__6070 (
            .O(N__27044),
            .I(N__27041));
    LocalMux I__6069 (
            .O(N__27041),
            .I(n5454));
    CascadeMux I__6068 (
            .O(N__27038),
            .I(N__27033));
    InMux I__6067 (
            .O(N__27037),
            .I(N__27029));
    InMux I__6066 (
            .O(N__27036),
            .I(N__27024));
    InMux I__6065 (
            .O(N__27033),
            .I(N__27021));
    InMux I__6064 (
            .O(N__27032),
            .I(N__27018));
    LocalMux I__6063 (
            .O(N__27029),
            .I(N__27015));
    InMux I__6062 (
            .O(N__27028),
            .I(N__27012));
    InMux I__6061 (
            .O(N__27027),
            .I(N__27009));
    LocalMux I__6060 (
            .O(N__27024),
            .I(N__27006));
    LocalMux I__6059 (
            .O(N__27021),
            .I(\eeprom.i2c.counter_1 ));
    LocalMux I__6058 (
            .O(N__27018),
            .I(\eeprom.i2c.counter_1 ));
    Odrv4 I__6057 (
            .O(N__27015),
            .I(\eeprom.i2c.counter_1 ));
    LocalMux I__6056 (
            .O(N__27012),
            .I(\eeprom.i2c.counter_1 ));
    LocalMux I__6055 (
            .O(N__27009),
            .I(\eeprom.i2c.counter_1 ));
    Odrv4 I__6054 (
            .O(N__27006),
            .I(\eeprom.i2c.counter_1 ));
    InMux I__6053 (
            .O(N__26993),
            .I(N__26990));
    LocalMux I__6052 (
            .O(N__26990),
            .I(N__26983));
    InMux I__6051 (
            .O(N__26989),
            .I(N__26979));
    InMux I__6050 (
            .O(N__26988),
            .I(N__26976));
    InMux I__6049 (
            .O(N__26987),
            .I(N__26971));
    InMux I__6048 (
            .O(N__26986),
            .I(N__26971));
    Span4Mux_v I__6047 (
            .O(N__26983),
            .I(N__26968));
    InMux I__6046 (
            .O(N__26982),
            .I(N__26965));
    LocalMux I__6045 (
            .O(N__26979),
            .I(N__26962));
    LocalMux I__6044 (
            .O(N__26976),
            .I(\eeprom.i2c.counter_2 ));
    LocalMux I__6043 (
            .O(N__26971),
            .I(\eeprom.i2c.counter_2 ));
    Odrv4 I__6042 (
            .O(N__26968),
            .I(\eeprom.i2c.counter_2 ));
    LocalMux I__6041 (
            .O(N__26965),
            .I(\eeprom.i2c.counter_2 ));
    Odrv4 I__6040 (
            .O(N__26962),
            .I(\eeprom.i2c.counter_2 ));
    CascadeMux I__6039 (
            .O(N__26951),
            .I(N__26944));
    InMux I__6038 (
            .O(N__26950),
            .I(N__26941));
    InMux I__6037 (
            .O(N__26949),
            .I(N__26936));
    InMux I__6036 (
            .O(N__26948),
            .I(N__26936));
    InMux I__6035 (
            .O(N__26947),
            .I(N__26933));
    InMux I__6034 (
            .O(N__26944),
            .I(N__26930));
    LocalMux I__6033 (
            .O(N__26941),
            .I(N__26927));
    LocalMux I__6032 (
            .O(N__26936),
            .I(\eeprom.i2c.counter_0 ));
    LocalMux I__6031 (
            .O(N__26933),
            .I(\eeprom.i2c.counter_0 ));
    LocalMux I__6030 (
            .O(N__26930),
            .I(\eeprom.i2c.counter_0 ));
    Odrv4 I__6029 (
            .O(N__26927),
            .I(\eeprom.i2c.counter_0 ));
    CascadeMux I__6028 (
            .O(N__26918),
            .I(\eeprom.i2c.n5464_cascade_ ));
    CascadeMux I__6027 (
            .O(N__26915),
            .I(\eeprom.i2c.n5451_cascade_ ));
    InMux I__6026 (
            .O(N__26912),
            .I(N__26909));
    LocalMux I__6025 (
            .O(N__26909),
            .I(\eeprom.i2c.sda_out ));
    CEMux I__6024 (
            .O(N__26906),
            .I(N__26903));
    LocalMux I__6023 (
            .O(N__26903),
            .I(N__26900));
    Odrv12 I__6022 (
            .O(N__26900),
            .I(\eeprom.i2c.n4513 ));
    CascadeMux I__6021 (
            .O(N__26897),
            .I(N__26888));
    CascadeMux I__6020 (
            .O(N__26896),
            .I(N__26882));
    CascadeMux I__6019 (
            .O(N__26895),
            .I(N__26879));
    InMux I__6018 (
            .O(N__26894),
            .I(N__26872));
    InMux I__6017 (
            .O(N__26893),
            .I(N__26872));
    InMux I__6016 (
            .O(N__26892),
            .I(N__26869));
    InMux I__6015 (
            .O(N__26891),
            .I(N__26866));
    InMux I__6014 (
            .O(N__26888),
            .I(N__26861));
    InMux I__6013 (
            .O(N__26887),
            .I(N__26861));
    InMux I__6012 (
            .O(N__26886),
            .I(N__26858));
    CascadeMux I__6011 (
            .O(N__26885),
            .I(N__26855));
    InMux I__6010 (
            .O(N__26882),
            .I(N__26850));
    InMux I__6009 (
            .O(N__26879),
            .I(N__26847));
    CascadeMux I__6008 (
            .O(N__26878),
            .I(N__26844));
    CascadeMux I__6007 (
            .O(N__26877),
            .I(N__26841));
    LocalMux I__6006 (
            .O(N__26872),
            .I(N__26836));
    LocalMux I__6005 (
            .O(N__26869),
            .I(N__26833));
    LocalMux I__6004 (
            .O(N__26866),
            .I(N__26828));
    LocalMux I__6003 (
            .O(N__26861),
            .I(N__26828));
    LocalMux I__6002 (
            .O(N__26858),
            .I(N__26825));
    InMux I__6001 (
            .O(N__26855),
            .I(N__26820));
    InMux I__6000 (
            .O(N__26854),
            .I(N__26820));
    InMux I__5999 (
            .O(N__26853),
            .I(N__26812));
    LocalMux I__5998 (
            .O(N__26850),
            .I(N__26807));
    LocalMux I__5997 (
            .O(N__26847),
            .I(N__26807));
    InMux I__5996 (
            .O(N__26844),
            .I(N__26798));
    InMux I__5995 (
            .O(N__26841),
            .I(N__26798));
    InMux I__5994 (
            .O(N__26840),
            .I(N__26798));
    InMux I__5993 (
            .O(N__26839),
            .I(N__26798));
    Span4Mux_h I__5992 (
            .O(N__26836),
            .I(N__26795));
    Span4Mux_v I__5991 (
            .O(N__26833),
            .I(N__26790));
    Span4Mux_h I__5990 (
            .O(N__26828),
            .I(N__26790));
    Span4Mux_h I__5989 (
            .O(N__26825),
            .I(N__26785));
    LocalMux I__5988 (
            .O(N__26820),
            .I(N__26785));
    InMux I__5987 (
            .O(N__26819),
            .I(N__26782));
    InMux I__5986 (
            .O(N__26818),
            .I(N__26775));
    InMux I__5985 (
            .O(N__26817),
            .I(N__26775));
    InMux I__5984 (
            .O(N__26816),
            .I(N__26775));
    InMux I__5983 (
            .O(N__26815),
            .I(N__26772));
    LocalMux I__5982 (
            .O(N__26812),
            .I(state_2));
    Odrv4 I__5981 (
            .O(N__26807),
            .I(state_2));
    LocalMux I__5980 (
            .O(N__26798),
            .I(state_2));
    Odrv4 I__5979 (
            .O(N__26795),
            .I(state_2));
    Odrv4 I__5978 (
            .O(N__26790),
            .I(state_2));
    Odrv4 I__5977 (
            .O(N__26785),
            .I(state_2));
    LocalMux I__5976 (
            .O(N__26782),
            .I(state_2));
    LocalMux I__5975 (
            .O(N__26775),
            .I(state_2));
    LocalMux I__5974 (
            .O(N__26772),
            .I(state_2));
    InMux I__5973 (
            .O(N__26753),
            .I(N__26747));
    InMux I__5972 (
            .O(N__26752),
            .I(N__26747));
    LocalMux I__5971 (
            .O(N__26747),
            .I(n3595));
    CascadeMux I__5970 (
            .O(N__26744),
            .I(N__26732));
    InMux I__5969 (
            .O(N__26743),
            .I(N__26724));
    InMux I__5968 (
            .O(N__26742),
            .I(N__26724));
    InMux I__5967 (
            .O(N__26741),
            .I(N__26724));
    InMux I__5966 (
            .O(N__26740),
            .I(N__26721));
    CascadeMux I__5965 (
            .O(N__26739),
            .I(N__26717));
    CascadeMux I__5964 (
            .O(N__26738),
            .I(N__26713));
    CascadeMux I__5963 (
            .O(N__26737),
            .I(N__26709));
    InMux I__5962 (
            .O(N__26736),
            .I(N__26699));
    InMux I__5961 (
            .O(N__26735),
            .I(N__26699));
    InMux I__5960 (
            .O(N__26732),
            .I(N__26699));
    InMux I__5959 (
            .O(N__26731),
            .I(N__26699));
    LocalMux I__5958 (
            .O(N__26724),
            .I(N__26694));
    LocalMux I__5957 (
            .O(N__26721),
            .I(N__26694));
    InMux I__5956 (
            .O(N__26720),
            .I(N__26679));
    InMux I__5955 (
            .O(N__26717),
            .I(N__26679));
    InMux I__5954 (
            .O(N__26716),
            .I(N__26679));
    InMux I__5953 (
            .O(N__26713),
            .I(N__26679));
    InMux I__5952 (
            .O(N__26712),
            .I(N__26679));
    InMux I__5951 (
            .O(N__26709),
            .I(N__26679));
    InMux I__5950 (
            .O(N__26708),
            .I(N__26679));
    LocalMux I__5949 (
            .O(N__26699),
            .I(N__26676));
    Span4Mux_v I__5948 (
            .O(N__26694),
            .I(N__26673));
    LocalMux I__5947 (
            .O(N__26679),
            .I(N__26670));
    Span4Mux_v I__5946 (
            .O(N__26676),
            .I(N__26663));
    Span4Mux_h I__5945 (
            .O(N__26673),
            .I(N__26663));
    Span4Mux_v I__5944 (
            .O(N__26670),
            .I(N__26663));
    Sp12to4 I__5943 (
            .O(N__26663),
            .I(N__26660));
    Span12Mux_h I__5942 (
            .O(N__26660),
            .I(N__26656));
    InMux I__5941 (
            .O(N__26659),
            .I(N__26653));
    Odrv12 I__5940 (
            .O(N__26656),
            .I(\eeprom.n2 ));
    LocalMux I__5939 (
            .O(N__26653),
            .I(\eeprom.n2 ));
    InMux I__5938 (
            .O(N__26648),
            .I(\eeprom.n4272 ));
    CascadeMux I__5937 (
            .O(N__26645),
            .I(N__26642));
    InMux I__5936 (
            .O(N__26642),
            .I(N__26638));
    InMux I__5935 (
            .O(N__26641),
            .I(N__26635));
    LocalMux I__5934 (
            .O(N__26638),
            .I(\eeprom.i2c.counter_3 ));
    LocalMux I__5933 (
            .O(N__26635),
            .I(\eeprom.i2c.counter_3 ));
    CascadeMux I__5932 (
            .O(N__26630),
            .I(N__26627));
    InMux I__5931 (
            .O(N__26627),
            .I(N__26623));
    InMux I__5930 (
            .O(N__26626),
            .I(N__26620));
    LocalMux I__5929 (
            .O(N__26623),
            .I(\eeprom.i2c.counter_5 ));
    LocalMux I__5928 (
            .O(N__26620),
            .I(\eeprom.i2c.counter_5 ));
    InMux I__5927 (
            .O(N__26615),
            .I(N__26611));
    InMux I__5926 (
            .O(N__26614),
            .I(N__26608));
    LocalMux I__5925 (
            .O(N__26611),
            .I(\eeprom.i2c.counter_4 ));
    LocalMux I__5924 (
            .O(N__26608),
            .I(\eeprom.i2c.counter_4 ));
    InMux I__5923 (
            .O(N__26603),
            .I(N__26599));
    InMux I__5922 (
            .O(N__26602),
            .I(N__26596));
    LocalMux I__5921 (
            .O(N__26599),
            .I(\eeprom.i2c.counter_7 ));
    LocalMux I__5920 (
            .O(N__26596),
            .I(\eeprom.i2c.counter_7 ));
    InMux I__5919 (
            .O(N__26591),
            .I(N__26587));
    InMux I__5918 (
            .O(N__26590),
            .I(N__26584));
    LocalMux I__5917 (
            .O(N__26587),
            .I(\eeprom.i2c.counter_6 ));
    LocalMux I__5916 (
            .O(N__26584),
            .I(\eeprom.i2c.counter_6 ));
    CascadeMux I__5915 (
            .O(N__26579),
            .I(\eeprom.i2c.n12_cascade_ ));
    CascadeMux I__5914 (
            .O(N__26576),
            .I(N__26573));
    InMux I__5913 (
            .O(N__26573),
            .I(N__26567));
    InMux I__5912 (
            .O(N__26572),
            .I(N__26567));
    LocalMux I__5911 (
            .O(N__26567),
            .I(\eeprom.i2c.n464 ));
    CascadeMux I__5910 (
            .O(N__26564),
            .I(N__26561));
    InMux I__5909 (
            .O(N__26561),
            .I(N__26557));
    InMux I__5908 (
            .O(N__26560),
            .I(N__26554));
    LocalMux I__5907 (
            .O(N__26557),
            .I(N__26551));
    LocalMux I__5906 (
            .O(N__26554),
            .I(N__26547));
    Span4Mux_h I__5905 (
            .O(N__26551),
            .I(N__26544));
    InMux I__5904 (
            .O(N__26550),
            .I(N__26541));
    Odrv4 I__5903 (
            .O(N__26547),
            .I(n4_adj_358));
    Odrv4 I__5902 (
            .O(N__26544),
            .I(n4_adj_358));
    LocalMux I__5901 (
            .O(N__26541),
            .I(n4_adj_358));
    CascadeMux I__5900 (
            .O(N__26534),
            .I(n10_cascade_));
    IoInMux I__5899 (
            .O(N__26531),
            .I(N__26528));
    LocalMux I__5898 (
            .O(N__26528),
            .I(N__26525));
    Span12Mux_s5_h I__5897 (
            .O(N__26525),
            .I(N__26516));
    CascadeMux I__5896 (
            .O(N__26524),
            .I(N__26510));
    InMux I__5895 (
            .O(N__26523),
            .I(N__26503));
    InMux I__5894 (
            .O(N__26522),
            .I(N__26503));
    InMux I__5893 (
            .O(N__26521),
            .I(N__26503));
    CascadeMux I__5892 (
            .O(N__26520),
            .I(N__26500));
    CascadeMux I__5891 (
            .O(N__26519),
            .I(N__26494));
    Span12Mux_v I__5890 (
            .O(N__26516),
            .I(N__26490));
    InMux I__5889 (
            .O(N__26515),
            .I(N__26481));
    InMux I__5888 (
            .O(N__26514),
            .I(N__26481));
    InMux I__5887 (
            .O(N__26513),
            .I(N__26481));
    InMux I__5886 (
            .O(N__26510),
            .I(N__26481));
    LocalMux I__5885 (
            .O(N__26503),
            .I(N__26478));
    InMux I__5884 (
            .O(N__26500),
            .I(N__26475));
    InMux I__5883 (
            .O(N__26499),
            .I(N__26468));
    InMux I__5882 (
            .O(N__26498),
            .I(N__26468));
    InMux I__5881 (
            .O(N__26497),
            .I(N__26468));
    InMux I__5880 (
            .O(N__26494),
            .I(N__26465));
    InMux I__5879 (
            .O(N__26493),
            .I(N__26462));
    Odrv12 I__5878 (
            .O(N__26490),
            .I(state_7_N_162_3));
    LocalMux I__5877 (
            .O(N__26481),
            .I(state_7_N_162_3));
    Odrv4 I__5876 (
            .O(N__26478),
            .I(state_7_N_162_3));
    LocalMux I__5875 (
            .O(N__26475),
            .I(state_7_N_162_3));
    LocalMux I__5874 (
            .O(N__26468),
            .I(state_7_N_162_3));
    LocalMux I__5873 (
            .O(N__26465),
            .I(state_7_N_162_3));
    LocalMux I__5872 (
            .O(N__26462),
            .I(state_7_N_162_3));
    InMux I__5871 (
            .O(N__26447),
            .I(N__26441));
    InMux I__5870 (
            .O(N__26446),
            .I(N__26441));
    LocalMux I__5869 (
            .O(N__26441),
            .I(\eeprom.i2c.n4579 ));
    CascadeMux I__5868 (
            .O(N__26438),
            .I(N__26435));
    InMux I__5867 (
            .O(N__26435),
            .I(N__26432));
    LocalMux I__5866 (
            .O(N__26432),
            .I(\eeprom.n10 ));
    InMux I__5865 (
            .O(N__26429),
            .I(N__26426));
    LocalMux I__5864 (
            .O(N__26426),
            .I(N__26423));
    Span12Mux_h I__5863 (
            .O(N__26423),
            .I(N__26420));
    Odrv12 I__5862 (
            .O(N__26420),
            .I(\eeprom.n10_adj_343 ));
    InMux I__5861 (
            .O(N__26417),
            .I(\eeprom.n4264 ));
    CascadeMux I__5860 (
            .O(N__26414),
            .I(N__26411));
    InMux I__5859 (
            .O(N__26411),
            .I(N__26408));
    LocalMux I__5858 (
            .O(N__26408),
            .I(\eeprom.n9 ));
    CascadeMux I__5857 (
            .O(N__26405),
            .I(N__26402));
    InMux I__5856 (
            .O(N__26402),
            .I(N__26399));
    LocalMux I__5855 (
            .O(N__26399),
            .I(\eeprom.n9_adj_308 ));
    InMux I__5854 (
            .O(N__26396),
            .I(bfn_27_26_0_));
    InMux I__5853 (
            .O(N__26393),
            .I(N__26390));
    LocalMux I__5852 (
            .O(N__26390),
            .I(N__26387));
    Span4Mux_h I__5851 (
            .O(N__26387),
            .I(N__26384));
    Odrv4 I__5850 (
            .O(N__26384),
            .I(\eeprom.n8_adj_311 ));
    InMux I__5849 (
            .O(N__26381),
            .I(\eeprom.n4266 ));
    CascadeMux I__5848 (
            .O(N__26378),
            .I(N__26375));
    InMux I__5847 (
            .O(N__26375),
            .I(N__26372));
    LocalMux I__5846 (
            .O(N__26372),
            .I(\eeprom.n7 ));
    InMux I__5845 (
            .O(N__26369),
            .I(\eeprom.n4267 ));
    CascadeMux I__5844 (
            .O(N__26366),
            .I(N__26363));
    InMux I__5843 (
            .O(N__26363),
            .I(N__26360));
    LocalMux I__5842 (
            .O(N__26360),
            .I(\eeprom.n6 ));
    InMux I__5841 (
            .O(N__26357),
            .I(N__26353));
    InMux I__5840 (
            .O(N__26356),
            .I(N__26350));
    LocalMux I__5839 (
            .O(N__26353),
            .I(N__26345));
    LocalMux I__5838 (
            .O(N__26350),
            .I(N__26345));
    Odrv12 I__5837 (
            .O(N__26345),
            .I(\eeprom.n6_adj_306 ));
    InMux I__5836 (
            .O(N__26342),
            .I(\eeprom.n4268 ));
    CascadeMux I__5835 (
            .O(N__26339),
            .I(N__26336));
    InMux I__5834 (
            .O(N__26336),
            .I(N__26333));
    LocalMux I__5833 (
            .O(N__26333),
            .I(\eeprom.n5 ));
    InMux I__5832 (
            .O(N__26330),
            .I(N__26327));
    LocalMux I__5831 (
            .O(N__26327),
            .I(N__26324));
    Odrv12 I__5830 (
            .O(N__26324),
            .I(\eeprom.n5_adj_317 ));
    InMux I__5829 (
            .O(N__26321),
            .I(\eeprom.n4269 ));
    CascadeMux I__5828 (
            .O(N__26318),
            .I(N__26315));
    InMux I__5827 (
            .O(N__26315),
            .I(N__26312));
    LocalMux I__5826 (
            .O(N__26312),
            .I(\eeprom.n4 ));
    InMux I__5825 (
            .O(N__26309),
            .I(\eeprom.n4270 ));
    CascadeMux I__5824 (
            .O(N__26306),
            .I(N__26303));
    InMux I__5823 (
            .O(N__26303),
            .I(N__26300));
    LocalMux I__5822 (
            .O(N__26300),
            .I(\eeprom.n3 ));
    InMux I__5821 (
            .O(N__26297),
            .I(N__26294));
    LocalMux I__5820 (
            .O(N__26294),
            .I(N__26291));
    Span4Mux_v I__5819 (
            .O(N__26291),
            .I(N__26288));
    Odrv4 I__5818 (
            .O(N__26288),
            .I(\eeprom.n3_adj_312 ));
    InMux I__5817 (
            .O(N__26285),
            .I(\eeprom.n4271 ));
    InMux I__5816 (
            .O(N__26282),
            .I(N__26279));
    LocalMux I__5815 (
            .O(N__26279),
            .I(N__26276));
    Span4Mux_h I__5814 (
            .O(N__26276),
            .I(N__26273));
    Odrv4 I__5813 (
            .O(N__26273),
            .I(\eeprom.n18_adj_326 ));
    InMux I__5812 (
            .O(N__26270),
            .I(\eeprom.n4256 ));
    CascadeMux I__5811 (
            .O(N__26267),
            .I(N__26264));
    InMux I__5810 (
            .O(N__26264),
            .I(N__26261));
    LocalMux I__5809 (
            .O(N__26261),
            .I(\eeprom.n17 ));
    InMux I__5808 (
            .O(N__26258),
            .I(N__26255));
    LocalMux I__5807 (
            .O(N__26255),
            .I(N__26252));
    Odrv12 I__5806 (
            .O(N__26252),
            .I(\eeprom.n17_adj_324 ));
    InMux I__5805 (
            .O(N__26249),
            .I(bfn_27_25_0_));
    CascadeMux I__5804 (
            .O(N__26246),
            .I(N__26243));
    InMux I__5803 (
            .O(N__26243),
            .I(N__26240));
    LocalMux I__5802 (
            .O(N__26240),
            .I(\eeprom.n16_adj_294 ));
    InMux I__5801 (
            .O(N__26237),
            .I(N__26234));
    LocalMux I__5800 (
            .O(N__26234),
            .I(N__26231));
    Odrv12 I__5799 (
            .O(N__26231),
            .I(\eeprom.n16_adj_325 ));
    InMux I__5798 (
            .O(N__26228),
            .I(\eeprom.n4258 ));
    CascadeMux I__5797 (
            .O(N__26225),
            .I(N__26222));
    InMux I__5796 (
            .O(N__26222),
            .I(N__26219));
    LocalMux I__5795 (
            .O(N__26219),
            .I(\eeprom.n15_adj_295 ));
    InMux I__5794 (
            .O(N__26216),
            .I(N__26213));
    LocalMux I__5793 (
            .O(N__26213),
            .I(N__26210));
    Span4Mux_h I__5792 (
            .O(N__26210),
            .I(N__26207));
    Odrv4 I__5791 (
            .O(N__26207),
            .I(\eeprom.n15 ));
    InMux I__5790 (
            .O(N__26204),
            .I(\eeprom.n4259 ));
    InMux I__5789 (
            .O(N__26201),
            .I(N__26198));
    LocalMux I__5788 (
            .O(N__26198),
            .I(N__26195));
    Odrv12 I__5787 (
            .O(N__26195),
            .I(\eeprom.n14 ));
    InMux I__5786 (
            .O(N__26192),
            .I(\eeprom.n4260 ));
    CascadeMux I__5785 (
            .O(N__26189),
            .I(N__26186));
    InMux I__5784 (
            .O(N__26186),
            .I(N__26183));
    LocalMux I__5783 (
            .O(N__26183),
            .I(N__26180));
    Span4Mux_v I__5782 (
            .O(N__26180),
            .I(N__26177));
    Odrv4 I__5781 (
            .O(N__26177),
            .I(\eeprom.n13 ));
    InMux I__5780 (
            .O(N__26174),
            .I(N__26171));
    LocalMux I__5779 (
            .O(N__26171),
            .I(N__26168));
    Span4Mux_v I__5778 (
            .O(N__26168),
            .I(N__26165));
    Odrv4 I__5777 (
            .O(N__26165),
            .I(\eeprom.n13_adj_318 ));
    InMux I__5776 (
            .O(N__26162),
            .I(\eeprom.n4261 ));
    CascadeMux I__5775 (
            .O(N__26159),
            .I(N__26156));
    InMux I__5774 (
            .O(N__26156),
            .I(N__26153));
    LocalMux I__5773 (
            .O(N__26153),
            .I(\eeprom.n12_adj_298 ));
    InMux I__5772 (
            .O(N__26150),
            .I(N__26147));
    LocalMux I__5771 (
            .O(N__26147),
            .I(N__26144));
    Span4Mux_v I__5770 (
            .O(N__26144),
            .I(N__26141));
    Span4Mux_h I__5769 (
            .O(N__26141),
            .I(N__26138));
    Odrv4 I__5768 (
            .O(N__26138),
            .I(\eeprom.n12_adj_319 ));
    InMux I__5767 (
            .O(N__26135),
            .I(\eeprom.n4262 ));
    CascadeMux I__5766 (
            .O(N__26132),
            .I(N__26129));
    InMux I__5765 (
            .O(N__26129),
            .I(N__26126));
    LocalMux I__5764 (
            .O(N__26126),
            .I(\eeprom.n11_adj_299 ));
    InMux I__5763 (
            .O(N__26123),
            .I(N__26120));
    LocalMux I__5762 (
            .O(N__26120),
            .I(N__26117));
    Span4Mux_v I__5761 (
            .O(N__26117),
            .I(N__26114));
    Odrv4 I__5760 (
            .O(N__26114),
            .I(\eeprom.n11 ));
    InMux I__5759 (
            .O(N__26111),
            .I(\eeprom.n4263 ));
    CascadeMux I__5758 (
            .O(N__26108),
            .I(N__26105));
    InMux I__5757 (
            .O(N__26105),
            .I(N__26102));
    LocalMux I__5756 (
            .O(N__26102),
            .I(N__26099));
    Odrv4 I__5755 (
            .O(N__26099),
            .I(\eeprom.n26_adj_276 ));
    InMux I__5754 (
            .O(N__26096),
            .I(N__26093));
    LocalMux I__5753 (
            .O(N__26093),
            .I(N__26090));
    Span4Mux_v I__5752 (
            .O(N__26090),
            .I(N__26087));
    Odrv4 I__5751 (
            .O(N__26087),
            .I(\eeprom.n26_adj_275 ));
    InMux I__5750 (
            .O(N__26084),
            .I(\eeprom.n4248 ));
    InMux I__5749 (
            .O(N__26081),
            .I(bfn_27_24_0_));
    InMux I__5748 (
            .O(N__26078),
            .I(N__26075));
    LocalMux I__5747 (
            .O(N__26075),
            .I(N__26072));
    Span4Mux_h I__5746 (
            .O(N__26072),
            .I(N__26069));
    Odrv4 I__5745 (
            .O(N__26069),
            .I(\eeprom.n24_adj_269 ));
    InMux I__5744 (
            .O(N__26066),
            .I(\eeprom.n4250 ));
    CascadeMux I__5743 (
            .O(N__26063),
            .I(N__26060));
    InMux I__5742 (
            .O(N__26060),
            .I(N__26057));
    LocalMux I__5741 (
            .O(N__26057),
            .I(N__26054));
    Odrv4 I__5740 (
            .O(N__26054),
            .I(\eeprom.n23_adj_268 ));
    InMux I__5739 (
            .O(N__26051),
            .I(N__26048));
    LocalMux I__5738 (
            .O(N__26048),
            .I(N__26045));
    Odrv12 I__5737 (
            .O(N__26045),
            .I(\eeprom.n23 ));
    InMux I__5736 (
            .O(N__26042),
            .I(\eeprom.n4251 ));
    InMux I__5735 (
            .O(N__26039),
            .I(N__26036));
    LocalMux I__5734 (
            .O(N__26036),
            .I(N__26033));
    Span4Mux_h I__5733 (
            .O(N__26033),
            .I(N__26030));
    Odrv4 I__5732 (
            .O(N__26030),
            .I(\eeprom.n22_adj_265 ));
    InMux I__5731 (
            .O(N__26027),
            .I(\eeprom.n4252 ));
    CascadeMux I__5730 (
            .O(N__26024),
            .I(N__26021));
    InMux I__5729 (
            .O(N__26021),
            .I(N__26018));
    LocalMux I__5728 (
            .O(N__26018),
            .I(N__26015));
    Odrv4 I__5727 (
            .O(N__26015),
            .I(\eeprom.n21_adj_264 ));
    InMux I__5726 (
            .O(N__26012),
            .I(N__26009));
    LocalMux I__5725 (
            .O(N__26009),
            .I(N__26006));
    Span4Mux_v I__5724 (
            .O(N__26006),
            .I(N__26003));
    Odrv4 I__5723 (
            .O(N__26003),
            .I(\eeprom.n21 ));
    InMux I__5722 (
            .O(N__26000),
            .I(\eeprom.n4253 ));
    CascadeMux I__5721 (
            .O(N__25997),
            .I(N__25994));
    InMux I__5720 (
            .O(N__25994),
            .I(N__25991));
    LocalMux I__5719 (
            .O(N__25991),
            .I(N__25988));
    Span4Mux_v I__5718 (
            .O(N__25988),
            .I(N__25985));
    Odrv4 I__5717 (
            .O(N__25985),
            .I(\eeprom.n20_adj_259 ));
    InMux I__5716 (
            .O(N__25982),
            .I(N__25979));
    LocalMux I__5715 (
            .O(N__25979),
            .I(N__25976));
    Span4Mux_h I__5714 (
            .O(N__25976),
            .I(N__25973));
    Odrv4 I__5713 (
            .O(N__25973),
            .I(\eeprom.n20 ));
    InMux I__5712 (
            .O(N__25970),
            .I(\eeprom.n4254 ));
    InMux I__5711 (
            .O(N__25967),
            .I(N__25964));
    LocalMux I__5710 (
            .O(N__25964),
            .I(N__25961));
    Span4Mux_h I__5709 (
            .O(N__25961),
            .I(N__25958));
    Odrv4 I__5708 (
            .O(N__25958),
            .I(\eeprom.n19_adj_320 ));
    InMux I__5707 (
            .O(N__25955),
            .I(\eeprom.n4255 ));
    CascadeMux I__5706 (
            .O(N__25952),
            .I(\eeprom.n1138_cascade_ ));
    CascadeMux I__5705 (
            .O(N__25949),
            .I(N__25946));
    InMux I__5704 (
            .O(N__25946),
            .I(N__25943));
    LocalMux I__5703 (
            .O(N__25943),
            .I(N__25940));
    Odrv4 I__5702 (
            .O(N__25940),
            .I(\eeprom.n33_adj_289 ));
    InMux I__5701 (
            .O(N__25937),
            .I(N__25934));
    LocalMux I__5700 (
            .O(N__25934),
            .I(N__25931));
    Odrv12 I__5699 (
            .O(N__25931),
            .I(\eeprom.n33 ));
    InMux I__5698 (
            .O(N__25928),
            .I(bfn_27_23_0_));
    CascadeMux I__5697 (
            .O(N__25925),
            .I(N__25922));
    InMux I__5696 (
            .O(N__25922),
            .I(N__25919));
    LocalMux I__5695 (
            .O(N__25919),
            .I(\eeprom.n32_adj_288 ));
    InMux I__5694 (
            .O(N__25916),
            .I(N__25913));
    LocalMux I__5693 (
            .O(N__25913),
            .I(N__25910));
    Span4Mux_v I__5692 (
            .O(N__25910),
            .I(N__25907));
    Span4Mux_v I__5691 (
            .O(N__25907),
            .I(N__25904));
    Odrv4 I__5690 (
            .O(N__25904),
            .I(\eeprom.n32_adj_287 ));
    InMux I__5689 (
            .O(N__25901),
            .I(\eeprom.n4242 ));
    CascadeMux I__5688 (
            .O(N__25898),
            .I(N__25895));
    InMux I__5687 (
            .O(N__25895),
            .I(N__25892));
    LocalMux I__5686 (
            .O(N__25892),
            .I(N__25889));
    Span4Mux_h I__5685 (
            .O(N__25889),
            .I(N__25886));
    Odrv4 I__5684 (
            .O(N__25886),
            .I(\eeprom.n31_adj_286 ));
    InMux I__5683 (
            .O(N__25883),
            .I(N__25880));
    LocalMux I__5682 (
            .O(N__25880),
            .I(N__25877));
    Span4Mux_v I__5681 (
            .O(N__25877),
            .I(N__25874));
    Odrv4 I__5680 (
            .O(N__25874),
            .I(\eeprom.n31_adj_285 ));
    InMux I__5679 (
            .O(N__25871),
            .I(\eeprom.n4243 ));
    InMux I__5678 (
            .O(N__25868),
            .I(N__25865));
    LocalMux I__5677 (
            .O(N__25865),
            .I(N__25862));
    Odrv4 I__5676 (
            .O(N__25862),
            .I(\eeprom.n30_adj_277 ));
    InMux I__5675 (
            .O(N__25859),
            .I(N__25856));
    LocalMux I__5674 (
            .O(N__25856),
            .I(N__25853));
    Odrv4 I__5673 (
            .O(N__25853),
            .I(\eeprom.n30_adj_284 ));
    InMux I__5672 (
            .O(N__25850),
            .I(\eeprom.n4244 ));
    CascadeMux I__5671 (
            .O(N__25847),
            .I(N__25844));
    InMux I__5670 (
            .O(N__25844),
            .I(N__25841));
    LocalMux I__5669 (
            .O(N__25841),
            .I(N__25838));
    Odrv4 I__5668 (
            .O(N__25838),
            .I(\eeprom.n29_adj_278 ));
    CascadeMux I__5667 (
            .O(N__25835),
            .I(N__25832));
    InMux I__5666 (
            .O(N__25832),
            .I(N__25829));
    LocalMux I__5665 (
            .O(N__25829),
            .I(N__25826));
    Span4Mux_v I__5664 (
            .O(N__25826),
            .I(N__25823));
    Odrv4 I__5663 (
            .O(N__25823),
            .I(\eeprom.n29_adj_283 ));
    InMux I__5662 (
            .O(N__25820),
            .I(\eeprom.n4245 ));
    CascadeMux I__5661 (
            .O(N__25817),
            .I(N__25814));
    InMux I__5660 (
            .O(N__25814),
            .I(N__25811));
    LocalMux I__5659 (
            .O(N__25811),
            .I(N__25808));
    Span4Mux_v I__5658 (
            .O(N__25808),
            .I(N__25805));
    Odrv4 I__5657 (
            .O(N__25805),
            .I(\eeprom.n28_adj_279 ));
    InMux I__5656 (
            .O(N__25802),
            .I(N__25799));
    LocalMux I__5655 (
            .O(N__25799),
            .I(N__25796));
    Span4Mux_h I__5654 (
            .O(N__25796),
            .I(N__25793));
    Span4Mux_v I__5653 (
            .O(N__25793),
            .I(N__25790));
    Odrv4 I__5652 (
            .O(N__25790),
            .I(\eeprom.n28_adj_282 ));
    InMux I__5651 (
            .O(N__25787),
            .I(\eeprom.n4246 ));
    CascadeMux I__5650 (
            .O(N__25784),
            .I(N__25781));
    InMux I__5649 (
            .O(N__25781),
            .I(N__25778));
    LocalMux I__5648 (
            .O(N__25778),
            .I(\eeprom.n27_adj_280 ));
    InMux I__5647 (
            .O(N__25775),
            .I(\eeprom.n4247 ));
    InMux I__5646 (
            .O(N__25772),
            .I(N__25769));
    LocalMux I__5645 (
            .O(N__25769),
            .I(N__25766));
    Span4Mux_h I__5644 (
            .O(N__25766),
            .I(N__25763));
    Span4Mux_h I__5643 (
            .O(N__25763),
            .I(N__25757));
    InMux I__5642 (
            .O(N__25762),
            .I(N__25754));
    InMux I__5641 (
            .O(N__25761),
            .I(N__25751));
    InMux I__5640 (
            .O(N__25760),
            .I(N__25748));
    Odrv4 I__5639 (
            .O(N__25757),
            .I(\eeprom.eeprom_counter_3 ));
    LocalMux I__5638 (
            .O(N__25754),
            .I(\eeprom.eeprom_counter_3 ));
    LocalMux I__5637 (
            .O(N__25751),
            .I(\eeprom.eeprom_counter_3 ));
    LocalMux I__5636 (
            .O(N__25748),
            .I(\eeprom.eeprom_counter_3 ));
    CascadeMux I__5635 (
            .O(N__25739),
            .I(N__25736));
    InMux I__5634 (
            .O(N__25736),
            .I(N__25732));
    InMux I__5633 (
            .O(N__25735),
            .I(N__25729));
    LocalMux I__5632 (
            .O(N__25732),
            .I(N__25726));
    LocalMux I__5631 (
            .O(N__25729),
            .I(N__25723));
    Span4Mux_v I__5630 (
            .O(N__25726),
            .I(N__25719));
    Span4Mux_h I__5629 (
            .O(N__25723),
            .I(N__25716));
    InMux I__5628 (
            .O(N__25722),
            .I(N__25713));
    Odrv4 I__5627 (
            .O(N__25719),
            .I(\eeprom.n1916 ));
    Odrv4 I__5626 (
            .O(N__25716),
            .I(\eeprom.n1916 ));
    LocalMux I__5625 (
            .O(N__25713),
            .I(\eeprom.n1916 ));
    CascadeMux I__5624 (
            .O(N__25706),
            .I(\eeprom.n5035_cascade_ ));
    InMux I__5623 (
            .O(N__25703),
            .I(N__25700));
    LocalMux I__5622 (
            .O(N__25700),
            .I(N__25697));
    Span4Mux_h I__5621 (
            .O(N__25697),
            .I(N__25694));
    Odrv4 I__5620 (
            .O(N__25694),
            .I(\eeprom.n5039 ));
    InMux I__5619 (
            .O(N__25691),
            .I(N__25688));
    LocalMux I__5618 (
            .O(N__25688),
            .I(N__25684));
    InMux I__5617 (
            .O(N__25687),
            .I(N__25680));
    Span4Mux_v I__5616 (
            .O(N__25684),
            .I(N__25677));
    InMux I__5615 (
            .O(N__25683),
            .I(N__25674));
    LocalMux I__5614 (
            .O(N__25680),
            .I(\eeprom.eeprom_counter_12 ));
    Odrv4 I__5613 (
            .O(N__25677),
            .I(\eeprom.eeprom_counter_12 ));
    LocalMux I__5612 (
            .O(N__25674),
            .I(\eeprom.eeprom_counter_12 ));
    InMux I__5611 (
            .O(N__25667),
            .I(N__25664));
    LocalMux I__5610 (
            .O(N__25664),
            .I(N__25660));
    InMux I__5609 (
            .O(N__25663),
            .I(N__25657));
    Span4Mux_h I__5608 (
            .O(N__25660),
            .I(N__25654));
    LocalMux I__5607 (
            .O(N__25657),
            .I(N__25650));
    Span4Mux_v I__5606 (
            .O(N__25654),
            .I(N__25646));
    InMux I__5605 (
            .O(N__25653),
            .I(N__25643));
    Span4Mux_h I__5604 (
            .O(N__25650),
            .I(N__25640));
    InMux I__5603 (
            .O(N__25649),
            .I(N__25637));
    Odrv4 I__5602 (
            .O(N__25646),
            .I(\eeprom.eeprom_counter_1 ));
    LocalMux I__5601 (
            .O(N__25643),
            .I(\eeprom.eeprom_counter_1 ));
    Odrv4 I__5600 (
            .O(N__25640),
            .I(\eeprom.eeprom_counter_1 ));
    LocalMux I__5599 (
            .O(N__25637),
            .I(\eeprom.eeprom_counter_1 ));
    CascadeMux I__5598 (
            .O(N__25628),
            .I(\eeprom.n892_cascade_ ));
    InMux I__5597 (
            .O(N__25625),
            .I(N__25622));
    LocalMux I__5596 (
            .O(N__25622),
            .I(N__25618));
    InMux I__5595 (
            .O(N__25621),
            .I(N__25614));
    Span12Mux_h I__5594 (
            .O(N__25618),
            .I(N__25611));
    InMux I__5593 (
            .O(N__25617),
            .I(N__25608));
    LocalMux I__5592 (
            .O(N__25614),
            .I(\eeprom.eeprom_counter_10 ));
    Odrv12 I__5591 (
            .O(N__25611),
            .I(\eeprom.eeprom_counter_10 ));
    LocalMux I__5590 (
            .O(N__25608),
            .I(\eeprom.eeprom_counter_10 ));
    CascadeMux I__5589 (
            .O(N__25601),
            .I(N__25597));
    CascadeMux I__5588 (
            .O(N__25600),
            .I(N__25594));
    InMux I__5587 (
            .O(N__25597),
            .I(N__25590));
    InMux I__5586 (
            .O(N__25594),
            .I(N__25587));
    InMux I__5585 (
            .O(N__25593),
            .I(N__25584));
    LocalMux I__5584 (
            .O(N__25590),
            .I(N__25581));
    LocalMux I__5583 (
            .O(N__25587),
            .I(N__25578));
    LocalMux I__5582 (
            .O(N__25584),
            .I(\eeprom.eeprom_counter_28 ));
    Odrv4 I__5581 (
            .O(N__25581),
            .I(\eeprom.eeprom_counter_28 ));
    Odrv4 I__5580 (
            .O(N__25578),
            .I(\eeprom.eeprom_counter_28 ));
    CascadeMux I__5579 (
            .O(N__25571),
            .I(\eeprom.n1256_cascade_ ));
    InMux I__5578 (
            .O(N__25568),
            .I(N__25565));
    LocalMux I__5577 (
            .O(N__25565),
            .I(N__25561));
    InMux I__5576 (
            .O(N__25564),
            .I(N__25558));
    Span4Mux_v I__5575 (
            .O(N__25561),
            .I(N__25553));
    LocalMux I__5574 (
            .O(N__25558),
            .I(N__25553));
    Odrv4 I__5573 (
            .O(N__25553),
            .I(\eeprom.n1913 ));
    InMux I__5572 (
            .O(N__25550),
            .I(N__25547));
    LocalMux I__5571 (
            .O(N__25547),
            .I(\eeprom.i2c.n13 ));
    InMux I__5570 (
            .O(N__25544),
            .I(N__25541));
    LocalMux I__5569 (
            .O(N__25541),
            .I(N__25537));
    InMux I__5568 (
            .O(N__25540),
            .I(N__25533));
    Span4Mux_h I__5567 (
            .O(N__25537),
            .I(N__25530));
    InMux I__5566 (
            .O(N__25536),
            .I(N__25527));
    LocalMux I__5565 (
            .O(N__25533),
            .I(\eeprom.eeprom_counter_7 ));
    Odrv4 I__5564 (
            .O(N__25530),
            .I(\eeprom.eeprom_counter_7 ));
    LocalMux I__5563 (
            .O(N__25527),
            .I(\eeprom.eeprom_counter_7 ));
    CascadeMux I__5562 (
            .O(N__25520),
            .I(N__25516));
    InMux I__5561 (
            .O(N__25519),
            .I(N__25510));
    InMux I__5560 (
            .O(N__25516),
            .I(N__25510));
    InMux I__5559 (
            .O(N__25515),
            .I(N__25507));
    LocalMux I__5558 (
            .O(N__25510),
            .I(N__25502));
    LocalMux I__5557 (
            .O(N__25507),
            .I(N__25502));
    Span4Mux_v I__5556 (
            .O(N__25502),
            .I(N__25499));
    Odrv4 I__5555 (
            .O(N__25499),
            .I(\eeprom.n1918 ));
    InMux I__5554 (
            .O(N__25496),
            .I(N__25493));
    LocalMux I__5553 (
            .O(N__25493),
            .I(N__25490));
    Span4Mux_h I__5552 (
            .O(N__25490),
            .I(N__25486));
    CascadeMux I__5551 (
            .O(N__25489),
            .I(N__25481));
    Span4Mux_v I__5550 (
            .O(N__25486),
            .I(N__25478));
    InMux I__5549 (
            .O(N__25485),
            .I(N__25475));
    InMux I__5548 (
            .O(N__25484),
            .I(N__25472));
    InMux I__5547 (
            .O(N__25481),
            .I(N__25469));
    Odrv4 I__5546 (
            .O(N__25478),
            .I(\eeprom.eeprom_counter_0 ));
    LocalMux I__5545 (
            .O(N__25475),
            .I(\eeprom.eeprom_counter_0 ));
    LocalMux I__5544 (
            .O(N__25472),
            .I(\eeprom.eeprom_counter_0 ));
    LocalMux I__5543 (
            .O(N__25469),
            .I(\eeprom.eeprom_counter_0 ));
    InMux I__5542 (
            .O(N__25460),
            .I(N__25456));
    InMux I__5541 (
            .O(N__25459),
            .I(N__25453));
    LocalMux I__5540 (
            .O(N__25456),
            .I(N__25448));
    LocalMux I__5539 (
            .O(N__25453),
            .I(N__25448));
    Span4Mux_v I__5538 (
            .O(N__25448),
            .I(N__25445));
    Odrv4 I__5537 (
            .O(N__25445),
            .I(\eeprom.n1912 ));
    InMux I__5536 (
            .O(N__25442),
            .I(N__25439));
    LocalMux I__5535 (
            .O(N__25439),
            .I(N__25435));
    InMux I__5534 (
            .O(N__25438),
            .I(N__25431));
    Span4Mux_h I__5533 (
            .O(N__25435),
            .I(N__25428));
    InMux I__5532 (
            .O(N__25434),
            .I(N__25425));
    LocalMux I__5531 (
            .O(N__25431),
            .I(\eeprom.eeprom_counter_27 ));
    Odrv4 I__5530 (
            .O(N__25428),
            .I(\eeprom.eeprom_counter_27 ));
    LocalMux I__5529 (
            .O(N__25425),
            .I(\eeprom.eeprom_counter_27 ));
    CascadeMux I__5528 (
            .O(N__25418),
            .I(\eeprom.n1139_cascade_ ));
    InMux I__5527 (
            .O(N__25415),
            .I(N__25411));
    InMux I__5526 (
            .O(N__25414),
            .I(N__25408));
    LocalMux I__5525 (
            .O(N__25411),
            .I(\eeprom.i2c.n37 ));
    LocalMux I__5524 (
            .O(N__25408),
            .I(\eeprom.i2c.n37 ));
    CascadeMux I__5523 (
            .O(N__25403),
            .I(\eeprom.i2c.n37_cascade_ ));
    InMux I__5522 (
            .O(N__25400),
            .I(N__25394));
    InMux I__5521 (
            .O(N__25399),
            .I(N__25394));
    LocalMux I__5520 (
            .O(N__25394),
            .I(\eeprom.i2c.n33 ));
    CascadeMux I__5519 (
            .O(N__25391),
            .I(\eeprom.i2c.n39_cascade_ ));
    InMux I__5518 (
            .O(N__25388),
            .I(N__25385));
    LocalMux I__5517 (
            .O(N__25385),
            .I(\eeprom.i2c.n39 ));
    CascadeMux I__5516 (
            .O(N__25382),
            .I(\eeprom.i2c.n407_cascade_ ));
    CascadeMux I__5515 (
            .O(N__25379),
            .I(N__25376));
    InMux I__5514 (
            .O(N__25376),
            .I(N__25373));
    LocalMux I__5513 (
            .O(N__25373),
            .I(N__25370));
    Span4Mux_h I__5512 (
            .O(N__25370),
            .I(N__25367));
    Span4Mux_h I__5511 (
            .O(N__25367),
            .I(N__25364));
    Odrv4 I__5510 (
            .O(N__25364),
            .I(\eeprom.n917 ));
    InMux I__5509 (
            .O(N__25361),
            .I(N__25357));
    InMux I__5508 (
            .O(N__25360),
            .I(N__25354));
    LocalMux I__5507 (
            .O(N__25357),
            .I(N__25351));
    LocalMux I__5506 (
            .O(N__25354),
            .I(N__25348));
    Span4Mux_h I__5505 (
            .O(N__25351),
            .I(N__25345));
    Span4Mux_h I__5504 (
            .O(N__25348),
            .I(N__25341));
    Span4Mux_h I__5503 (
            .O(N__25345),
            .I(N__25337));
    InMux I__5502 (
            .O(N__25344),
            .I(N__25334));
    Span4Mux_h I__5501 (
            .O(N__25341),
            .I(N__25331));
    InMux I__5500 (
            .O(N__25340),
            .I(N__25328));
    Odrv4 I__5499 (
            .O(N__25337),
            .I(\eeprom.eeprom_counter_5 ));
    LocalMux I__5498 (
            .O(N__25334),
            .I(\eeprom.eeprom_counter_5 ));
    Odrv4 I__5497 (
            .O(N__25331),
            .I(\eeprom.eeprom_counter_5 ));
    LocalMux I__5496 (
            .O(N__25328),
            .I(\eeprom.eeprom_counter_5 ));
    InMux I__5495 (
            .O(N__25319),
            .I(N__25316));
    LocalMux I__5494 (
            .O(N__25316),
            .I(N__25313));
    Span4Mux_h I__5493 (
            .O(N__25313),
            .I(N__25310));
    Span4Mux_h I__5492 (
            .O(N__25310),
            .I(N__25307));
    Odrv4 I__5491 (
            .O(N__25307),
            .I(\eeprom.n3722 ));
    InMux I__5490 (
            .O(N__25304),
            .I(N__25301));
    LocalMux I__5489 (
            .O(N__25301),
            .I(N__25297));
    InMux I__5488 (
            .O(N__25300),
            .I(N__25293));
    Span4Mux_v I__5487 (
            .O(N__25297),
            .I(N__25290));
    InMux I__5486 (
            .O(N__25296),
            .I(N__25287));
    LocalMux I__5485 (
            .O(N__25293),
            .I(\eeprom.eeprom_counter_30 ));
    Odrv4 I__5484 (
            .O(N__25290),
            .I(\eeprom.eeprom_counter_30 ));
    LocalMux I__5483 (
            .O(N__25287),
            .I(\eeprom.eeprom_counter_30 ));
    InMux I__5482 (
            .O(N__25280),
            .I(N__25277));
    LocalMux I__5481 (
            .O(N__25277),
            .I(n4733));
    SRMux I__5480 (
            .O(N__25274),
            .I(N__25271));
    LocalMux I__5479 (
            .O(N__25271),
            .I(N__25268));
    Span4Mux_h I__5478 (
            .O(N__25268),
            .I(N__25265));
    Odrv4 I__5477 (
            .O(N__25265),
            .I(\eeprom.i2c.n1913 ));
    InMux I__5476 (
            .O(N__25262),
            .I(N__25259));
    LocalMux I__5475 (
            .O(N__25259),
            .I(\eeprom.i2c.n534 ));
    CEMux I__5474 (
            .O(N__25256),
            .I(N__25253));
    LocalMux I__5473 (
            .O(N__25253),
            .I(N__25250));
    Odrv12 I__5472 (
            .O(N__25250),
            .I(\eeprom.i2c.n1829 ));
    InMux I__5471 (
            .O(N__25247),
            .I(N__25241));
    InMux I__5470 (
            .O(N__25246),
            .I(N__25236));
    InMux I__5469 (
            .O(N__25245),
            .I(N__25236));
    InMux I__5468 (
            .O(N__25244),
            .I(N__25233));
    LocalMux I__5467 (
            .O(N__25241),
            .I(\eeprom.i2c.n9 ));
    LocalMux I__5466 (
            .O(N__25236),
            .I(\eeprom.i2c.n9 ));
    LocalMux I__5465 (
            .O(N__25233),
            .I(\eeprom.i2c.n9 ));
    CascadeMux I__5464 (
            .O(N__25226),
            .I(\eeprom.i2c.n9_cascade_ ));
    CascadeMux I__5463 (
            .O(N__25223),
            .I(N__25220));
    InMux I__5462 (
            .O(N__25220),
            .I(N__25217));
    LocalMux I__5461 (
            .O(N__25217),
            .I(N__25214));
    Odrv4 I__5460 (
            .O(N__25214),
            .I(n1814));
    CascadeMux I__5459 (
            .O(N__25211),
            .I(n1814_cascade_));
    InMux I__5458 (
            .O(N__25208),
            .I(bfn_27_17_0_));
    InMux I__5457 (
            .O(N__25205),
            .I(\eeprom.i2c.n3899 ));
    InMux I__5456 (
            .O(N__25202),
            .I(\eeprom.i2c.n3900 ));
    InMux I__5455 (
            .O(N__25199),
            .I(\eeprom.i2c.n3901 ));
    InMux I__5454 (
            .O(N__25196),
            .I(\eeprom.i2c.n3902 ));
    InMux I__5453 (
            .O(N__25193),
            .I(\eeprom.i2c.n3903 ));
    InMux I__5452 (
            .O(N__25190),
            .I(\eeprom.i2c.n3904 ));
    InMux I__5451 (
            .O(N__25187),
            .I(\eeprom.i2c.n3905 ));
    InMux I__5450 (
            .O(N__25184),
            .I(N__25179));
    InMux I__5449 (
            .O(N__25183),
            .I(N__25174));
    InMux I__5448 (
            .O(N__25182),
            .I(N__25174));
    LocalMux I__5447 (
            .O(N__25179),
            .I(n11));
    LocalMux I__5446 (
            .O(N__25174),
            .I(n11));
    InMux I__5445 (
            .O(N__25169),
            .I(N__25161));
    InMux I__5444 (
            .O(N__25168),
            .I(N__25161));
    InMux I__5443 (
            .O(N__25167),
            .I(N__25158));
    InMux I__5442 (
            .O(N__25166),
            .I(N__25155));
    LocalMux I__5441 (
            .O(N__25161),
            .I(N__25152));
    LocalMux I__5440 (
            .O(N__25158),
            .I(n10_adj_360));
    LocalMux I__5439 (
            .O(N__25155),
            .I(n10_adj_360));
    Odrv4 I__5438 (
            .O(N__25152),
            .I(n10_adj_360));
    InMux I__5437 (
            .O(N__25145),
            .I(N__25140));
    InMux I__5436 (
            .O(N__25144),
            .I(N__25137));
    InMux I__5435 (
            .O(N__25143),
            .I(N__25134));
    LocalMux I__5434 (
            .O(N__25140),
            .I(N__25127));
    LocalMux I__5433 (
            .O(N__25137),
            .I(N__25127));
    LocalMux I__5432 (
            .O(N__25134),
            .I(N__25127));
    Span12Mux_v I__5431 (
            .O(N__25127),
            .I(N__25124));
    Odrv12 I__5430 (
            .O(N__25124),
            .I(\eeprom.n1919 ));
    CascadeMux I__5429 (
            .O(N__25121),
            .I(N__25116));
    InMux I__5428 (
            .O(N__25120),
            .I(N__25113));
    InMux I__5427 (
            .O(N__25119),
            .I(N__25108));
    InMux I__5426 (
            .O(N__25116),
            .I(N__25108));
    LocalMux I__5425 (
            .O(N__25113),
            .I(\eeprom.eeprom_counter_24 ));
    LocalMux I__5424 (
            .O(N__25108),
            .I(\eeprom.eeprom_counter_24 ));
    InMux I__5423 (
            .O(N__25103),
            .I(N__25099));
    InMux I__5422 (
            .O(N__25102),
            .I(N__25095));
    LocalMux I__5421 (
            .O(N__25099),
            .I(N__25092));
    InMux I__5420 (
            .O(N__25098),
            .I(N__25089));
    LocalMux I__5419 (
            .O(N__25095),
            .I(N__25084));
    Span4Mux_v I__5418 (
            .O(N__25092),
            .I(N__25084));
    LocalMux I__5417 (
            .O(N__25089),
            .I(N__25081));
    Odrv4 I__5416 (
            .O(N__25084),
            .I(\eeprom.eeprom_counter_18 ));
    Odrv4 I__5415 (
            .O(N__25081),
            .I(\eeprom.eeprom_counter_18 ));
    InMux I__5414 (
            .O(N__25076),
            .I(N__25073));
    LocalMux I__5413 (
            .O(N__25073),
            .I(N__25068));
    InMux I__5412 (
            .O(N__25072),
            .I(N__25065));
    InMux I__5411 (
            .O(N__25071),
            .I(N__25062));
    Span4Mux_h I__5410 (
            .O(N__25068),
            .I(N__25059));
    LocalMux I__5409 (
            .O(N__25065),
            .I(N__25056));
    LocalMux I__5408 (
            .O(N__25062),
            .I(\eeprom.eeprom_counter_17 ));
    Odrv4 I__5407 (
            .O(N__25059),
            .I(\eeprom.eeprom_counter_17 ));
    Odrv12 I__5406 (
            .O(N__25056),
            .I(\eeprom.eeprom_counter_17 ));
    InMux I__5405 (
            .O(N__25049),
            .I(N__25046));
    LocalMux I__5404 (
            .O(N__25046),
            .I(N__25041));
    InMux I__5403 (
            .O(N__25045),
            .I(N__25038));
    InMux I__5402 (
            .O(N__25044),
            .I(N__25035));
    Span4Mux_v I__5401 (
            .O(N__25041),
            .I(N__25030));
    LocalMux I__5400 (
            .O(N__25038),
            .I(N__25030));
    LocalMux I__5399 (
            .O(N__25035),
            .I(\eeprom.eeprom_counter_22 ));
    Odrv4 I__5398 (
            .O(N__25030),
            .I(\eeprom.eeprom_counter_22 ));
    InMux I__5397 (
            .O(N__25025),
            .I(N__25022));
    LocalMux I__5396 (
            .O(N__25022),
            .I(N__25017));
    InMux I__5395 (
            .O(N__25021),
            .I(N__25014));
    InMux I__5394 (
            .O(N__25020),
            .I(N__25011));
    Span4Mux_v I__5393 (
            .O(N__25017),
            .I(N__25008));
    LocalMux I__5392 (
            .O(N__25014),
            .I(N__25005));
    LocalMux I__5391 (
            .O(N__25011),
            .I(\eeprom.eeprom_counter_21 ));
    Odrv4 I__5390 (
            .O(N__25008),
            .I(\eeprom.eeprom_counter_21 ));
    Odrv4 I__5389 (
            .O(N__25005),
            .I(\eeprom.eeprom_counter_21 ));
    InMux I__5388 (
            .O(N__24998),
            .I(\eeprom.n3957 ));
    InMux I__5387 (
            .O(N__24995),
            .I(\eeprom.n3958 ));
    InMux I__5386 (
            .O(N__24992),
            .I(\eeprom.n3959 ));
    InMux I__5385 (
            .O(N__24989),
            .I(\eeprom.n3960 ));
    InMux I__5384 (
            .O(N__24986),
            .I(\eeprom.n3961 ));
    InMux I__5383 (
            .O(N__24983),
            .I(N__24980));
    LocalMux I__5382 (
            .O(N__24980),
            .I(N__24975));
    InMux I__5381 (
            .O(N__24979),
            .I(N__24972));
    InMux I__5380 (
            .O(N__24978),
            .I(N__24969));
    Span4Mux_h I__5379 (
            .O(N__24975),
            .I(N__24966));
    LocalMux I__5378 (
            .O(N__24972),
            .I(N__24963));
    LocalMux I__5377 (
            .O(N__24969),
            .I(\eeprom.eeprom_counter_23 ));
    Odrv4 I__5376 (
            .O(N__24966),
            .I(\eeprom.eeprom_counter_23 ));
    Odrv4 I__5375 (
            .O(N__24963),
            .I(\eeprom.eeprom_counter_23 ));
    InMux I__5374 (
            .O(N__24956),
            .I(N__24952));
    CascadeMux I__5373 (
            .O(N__24955),
            .I(N__24949));
    LocalMux I__5372 (
            .O(N__24952),
            .I(N__24945));
    InMux I__5371 (
            .O(N__24949),
            .I(N__24942));
    InMux I__5370 (
            .O(N__24948),
            .I(N__24939));
    Span4Mux_h I__5369 (
            .O(N__24945),
            .I(N__24936));
    LocalMux I__5368 (
            .O(N__24942),
            .I(N__24933));
    LocalMux I__5367 (
            .O(N__24939),
            .I(\eeprom.eeprom_counter_16 ));
    Odrv4 I__5366 (
            .O(N__24936),
            .I(\eeprom.eeprom_counter_16 ));
    Odrv4 I__5365 (
            .O(N__24933),
            .I(\eeprom.eeprom_counter_16 ));
    InMux I__5364 (
            .O(N__24926),
            .I(\eeprom.n3948 ));
    InMux I__5363 (
            .O(N__24923),
            .I(\eeprom.n3949 ));
    CascadeMux I__5362 (
            .O(N__24920),
            .I(N__24916));
    InMux I__5361 (
            .O(N__24919),
            .I(N__24912));
    InMux I__5360 (
            .O(N__24916),
            .I(N__24909));
    InMux I__5359 (
            .O(N__24915),
            .I(N__24906));
    LocalMux I__5358 (
            .O(N__24912),
            .I(N__24903));
    LocalMux I__5357 (
            .O(N__24909),
            .I(N__24900));
    LocalMux I__5356 (
            .O(N__24906),
            .I(\eeprom.eeprom_counter_20 ));
    Odrv4 I__5355 (
            .O(N__24903),
            .I(\eeprom.eeprom_counter_20 ));
    Odrv4 I__5354 (
            .O(N__24900),
            .I(\eeprom.eeprom_counter_20 ));
    InMux I__5353 (
            .O(N__24893),
            .I(\eeprom.n3950 ));
    InMux I__5352 (
            .O(N__24890),
            .I(\eeprom.n3951 ));
    InMux I__5351 (
            .O(N__24887),
            .I(\eeprom.n3952 ));
    InMux I__5350 (
            .O(N__24884),
            .I(\eeprom.n3953 ));
    InMux I__5349 (
            .O(N__24881),
            .I(bfn_26_24_0_));
    InMux I__5348 (
            .O(N__24878),
            .I(\eeprom.n3955 ));
    InMux I__5347 (
            .O(N__24875),
            .I(\eeprom.n3956 ));
    InMux I__5346 (
            .O(N__24872),
            .I(\eeprom.n3939 ));
    InMux I__5345 (
            .O(N__24869),
            .I(\eeprom.n3940 ));
    InMux I__5344 (
            .O(N__24866),
            .I(\eeprom.n3941 ));
    InMux I__5343 (
            .O(N__24863),
            .I(\eeprom.n3942 ));
    InMux I__5342 (
            .O(N__24860),
            .I(N__24857));
    LocalMux I__5341 (
            .O(N__24857),
            .I(N__24852));
    InMux I__5340 (
            .O(N__24856),
            .I(N__24849));
    InMux I__5339 (
            .O(N__24855),
            .I(N__24846));
    Span4Mux_v I__5338 (
            .O(N__24852),
            .I(N__24843));
    LocalMux I__5337 (
            .O(N__24849),
            .I(N__24840));
    LocalMux I__5336 (
            .O(N__24846),
            .I(\eeprom.eeprom_counter_13 ));
    Odrv4 I__5335 (
            .O(N__24843),
            .I(\eeprom.eeprom_counter_13 ));
    Odrv4 I__5334 (
            .O(N__24840),
            .I(\eeprom.eeprom_counter_13 ));
    InMux I__5333 (
            .O(N__24833),
            .I(\eeprom.n3943 ));
    InMux I__5332 (
            .O(N__24830),
            .I(\eeprom.n3944 ));
    InMux I__5331 (
            .O(N__24827),
            .I(\eeprom.n3945 ));
    InMux I__5330 (
            .O(N__24824),
            .I(bfn_26_23_0_));
    InMux I__5329 (
            .O(N__24821),
            .I(\eeprom.n3947 ));
    InMux I__5328 (
            .O(N__24818),
            .I(bfn_26_21_0_));
    InMux I__5327 (
            .O(N__24815),
            .I(\eeprom.n3931 ));
    InMux I__5326 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__5325 (
            .O(N__24809),
            .I(N__24805));
    InMux I__5324 (
            .O(N__24808),
            .I(N__24802));
    Span4Mux_h I__5323 (
            .O(N__24805),
            .I(N__24799));
    LocalMux I__5322 (
            .O(N__24802),
            .I(N__24795));
    Span4Mux_h I__5321 (
            .O(N__24799),
            .I(N__24791));
    InMux I__5320 (
            .O(N__24798),
            .I(N__24788));
    Span4Mux_h I__5319 (
            .O(N__24795),
            .I(N__24785));
    InMux I__5318 (
            .O(N__24794),
            .I(N__24782));
    Odrv4 I__5317 (
            .O(N__24791),
            .I(\eeprom.eeprom_counter_2 ));
    LocalMux I__5316 (
            .O(N__24788),
            .I(\eeprom.eeprom_counter_2 ));
    Odrv4 I__5315 (
            .O(N__24785),
            .I(\eeprom.eeprom_counter_2 ));
    LocalMux I__5314 (
            .O(N__24782),
            .I(\eeprom.eeprom_counter_2 ));
    InMux I__5313 (
            .O(N__24773),
            .I(\eeprom.n3932 ));
    InMux I__5312 (
            .O(N__24770),
            .I(\eeprom.n3933 ));
    InMux I__5311 (
            .O(N__24767),
            .I(N__24764));
    LocalMux I__5310 (
            .O(N__24764),
            .I(N__24760));
    InMux I__5309 (
            .O(N__24763),
            .I(N__24757));
    Span4Mux_h I__5308 (
            .O(N__24760),
            .I(N__24754));
    LocalMux I__5307 (
            .O(N__24757),
            .I(N__24750));
    Span4Mux_v I__5306 (
            .O(N__24754),
            .I(N__24746));
    InMux I__5305 (
            .O(N__24753),
            .I(N__24743));
    Span4Mux_h I__5304 (
            .O(N__24750),
            .I(N__24740));
    InMux I__5303 (
            .O(N__24749),
            .I(N__24737));
    Odrv4 I__5302 (
            .O(N__24746),
            .I(\eeprom.eeprom_counter_4 ));
    LocalMux I__5301 (
            .O(N__24743),
            .I(\eeprom.eeprom_counter_4 ));
    Odrv4 I__5300 (
            .O(N__24740),
            .I(\eeprom.eeprom_counter_4 ));
    LocalMux I__5299 (
            .O(N__24737),
            .I(\eeprom.eeprom_counter_4 ));
    InMux I__5298 (
            .O(N__24728),
            .I(\eeprom.n3934 ));
    InMux I__5297 (
            .O(N__24725),
            .I(\eeprom.n3935 ));
    InMux I__5296 (
            .O(N__24722),
            .I(\eeprom.n3936 ));
    InMux I__5295 (
            .O(N__24719),
            .I(\eeprom.n3937 ));
    InMux I__5294 (
            .O(N__24716),
            .I(bfn_26_22_0_));
    InMux I__5293 (
            .O(N__24713),
            .I(N__24709));
    InMux I__5292 (
            .O(N__24712),
            .I(N__24706));
    LocalMux I__5291 (
            .O(N__24709),
            .I(N__24700));
    LocalMux I__5290 (
            .O(N__24706),
            .I(N__24700));
    InMux I__5289 (
            .O(N__24705),
            .I(N__24697));
    Odrv4 I__5288 (
            .O(N__24700),
            .I(n1805));
    LocalMux I__5287 (
            .O(N__24697),
            .I(n1805));
    InMux I__5286 (
            .O(N__24692),
            .I(N__24689));
    LocalMux I__5285 (
            .O(N__24689),
            .I(n158));
    InMux I__5284 (
            .O(N__24686),
            .I(N__24683));
    LocalMux I__5283 (
            .O(N__24683),
            .I(n8));
    CascadeMux I__5282 (
            .O(N__24680),
            .I(n5461_cascade_));
    InMux I__5281 (
            .O(N__24677),
            .I(N__24671));
    InMux I__5280 (
            .O(N__24676),
            .I(N__24671));
    LocalMux I__5279 (
            .O(N__24671),
            .I(N__24667));
    InMux I__5278 (
            .O(N__24670),
            .I(N__24664));
    Odrv4 I__5277 (
            .O(N__24667),
            .I(n1800));
    LocalMux I__5276 (
            .O(N__24664),
            .I(n1800));
    CascadeMux I__5275 (
            .O(N__24659),
            .I(N__24655));
    InMux I__5274 (
            .O(N__24658),
            .I(N__24650));
    InMux I__5273 (
            .O(N__24655),
            .I(N__24650));
    LocalMux I__5272 (
            .O(N__24650),
            .I(N__24647));
    Odrv4 I__5271 (
            .O(N__24647),
            .I(n3585));
    InMux I__5270 (
            .O(N__24644),
            .I(N__24641));
    LocalMux I__5269 (
            .O(N__24641),
            .I(n160));
    InMux I__5268 (
            .O(N__24638),
            .I(N__24635));
    LocalMux I__5267 (
            .O(N__24635),
            .I(N__24630));
    InMux I__5266 (
            .O(N__24634),
            .I(N__24627));
    InMux I__5265 (
            .O(N__24633),
            .I(N__24624));
    Span4Mux_h I__5264 (
            .O(N__24630),
            .I(N__24619));
    LocalMux I__5263 (
            .O(N__24627),
            .I(N__24619));
    LocalMux I__5262 (
            .O(N__24624),
            .I(N__24616));
    Span4Mux_v I__5261 (
            .O(N__24619),
            .I(N__24613));
    Span4Mux_h I__5260 (
            .O(N__24616),
            .I(N__24610));
    Span4Mux_h I__5259 (
            .O(N__24613),
            .I(N__24607));
    Odrv4 I__5258 (
            .O(N__24610),
            .I(\eeprom.n2119 ));
    Odrv4 I__5257 (
            .O(N__24607),
            .I(\eeprom.n2119 ));
    InMux I__5256 (
            .O(N__24602),
            .I(N__24597));
    InMux I__5255 (
            .O(N__24601),
            .I(N__24594));
    InMux I__5254 (
            .O(N__24600),
            .I(N__24591));
    LocalMux I__5253 (
            .O(N__24597),
            .I(N__24584));
    LocalMux I__5252 (
            .O(N__24594),
            .I(N__24584));
    LocalMux I__5251 (
            .O(N__24591),
            .I(N__24584));
    Odrv12 I__5250 (
            .O(N__24584),
            .I(\eeprom.n2319 ));
    InMux I__5249 (
            .O(N__24581),
            .I(N__24578));
    LocalMux I__5248 (
            .O(N__24578),
            .I(n172));
    CascadeMux I__5247 (
            .O(N__24575),
            .I(n22_adj_367_cascade_));
    CascadeMux I__5246 (
            .O(N__24572),
            .I(n4_adj_369_cascade_));
    CascadeMux I__5245 (
            .O(N__24569),
            .I(n4_cascade_));
    InMux I__5244 (
            .O(N__24566),
            .I(N__24563));
    LocalMux I__5243 (
            .O(N__24563),
            .I(n166));
    CascadeMux I__5242 (
            .O(N__24560),
            .I(N__24557));
    InMux I__5241 (
            .O(N__24557),
            .I(N__24554));
    LocalMux I__5240 (
            .O(N__24554),
            .I(n4));
    InMux I__5239 (
            .O(N__24551),
            .I(N__24548));
    LocalMux I__5238 (
            .O(N__24548),
            .I(n168));
    CascadeMux I__5237 (
            .O(N__24545),
            .I(n1805_cascade_));
    InMux I__5236 (
            .O(N__24542),
            .I(N__24539));
    LocalMux I__5235 (
            .O(N__24539),
            .I(n170));
    CascadeMux I__5234 (
            .O(N__24536),
            .I(n1800_cascade_));
    InMux I__5233 (
            .O(N__24533),
            .I(N__24530));
    LocalMux I__5232 (
            .O(N__24530),
            .I(n164));
    InMux I__5231 (
            .O(N__24527),
            .I(N__24524));
    LocalMux I__5230 (
            .O(N__24524),
            .I(n4_adj_361));
    CascadeMux I__5229 (
            .O(N__24521),
            .I(n4_adj_361_cascade_));
    InMux I__5228 (
            .O(N__24518),
            .I(N__24515));
    LocalMux I__5227 (
            .O(N__24515),
            .I(n162));
    CascadeMux I__5226 (
            .O(N__24512),
            .I(n5361_cascade_));
    CascadeMux I__5225 (
            .O(N__24509),
            .I(N__24505));
    InMux I__5224 (
            .O(N__24508),
            .I(N__24502));
    InMux I__5223 (
            .O(N__24505),
            .I(N__24499));
    LocalMux I__5222 (
            .O(N__24502),
            .I(N__24494));
    LocalMux I__5221 (
            .O(N__24499),
            .I(N__24494));
    Span4Mux_h I__5220 (
            .O(N__24494),
            .I(N__24490));
    InMux I__5219 (
            .O(N__24493),
            .I(N__24487));
    Odrv4 I__5218 (
            .O(N__24490),
            .I(\eeprom.n2508 ));
    LocalMux I__5217 (
            .O(N__24487),
            .I(\eeprom.n2508 ));
    CascadeMux I__5216 (
            .O(N__24482),
            .I(N__24479));
    InMux I__5215 (
            .O(N__24479),
            .I(N__24476));
    LocalMux I__5214 (
            .O(N__24476),
            .I(\eeprom.n2575 ));
    InMux I__5213 (
            .O(N__24473),
            .I(\eeprom.n4040 ));
    InMux I__5212 (
            .O(N__24470),
            .I(N__24466));
    InMux I__5211 (
            .O(N__24469),
            .I(N__24463));
    LocalMux I__5210 (
            .O(N__24466),
            .I(N__24457));
    LocalMux I__5209 (
            .O(N__24463),
            .I(N__24457));
    InMux I__5208 (
            .O(N__24462),
            .I(N__24454));
    Odrv4 I__5207 (
            .O(N__24457),
            .I(\eeprom.n2507 ));
    LocalMux I__5206 (
            .O(N__24454),
            .I(\eeprom.n2507 ));
    CascadeMux I__5205 (
            .O(N__24449),
            .I(N__24446));
    InMux I__5204 (
            .O(N__24446),
            .I(N__24443));
    LocalMux I__5203 (
            .O(N__24443),
            .I(\eeprom.n2574 ));
    InMux I__5202 (
            .O(N__24440),
            .I(\eeprom.n4041 ));
    CascadeMux I__5201 (
            .O(N__24437),
            .I(N__24428));
    CascadeMux I__5200 (
            .O(N__24436),
            .I(N__24423));
    CascadeMux I__5199 (
            .O(N__24435),
            .I(N__24419));
    InMux I__5198 (
            .O(N__24434),
            .I(N__24412));
    InMux I__5197 (
            .O(N__24433),
            .I(N__24412));
    CascadeMux I__5196 (
            .O(N__24432),
            .I(N__24409));
    InMux I__5195 (
            .O(N__24431),
            .I(N__24401));
    InMux I__5194 (
            .O(N__24428),
            .I(N__24401));
    InMux I__5193 (
            .O(N__24427),
            .I(N__24401));
    InMux I__5192 (
            .O(N__24426),
            .I(N__24398));
    InMux I__5191 (
            .O(N__24423),
            .I(N__24393));
    InMux I__5190 (
            .O(N__24422),
            .I(N__24393));
    InMux I__5189 (
            .O(N__24419),
            .I(N__24386));
    InMux I__5188 (
            .O(N__24418),
            .I(N__24386));
    InMux I__5187 (
            .O(N__24417),
            .I(N__24386));
    LocalMux I__5186 (
            .O(N__24412),
            .I(N__24383));
    InMux I__5185 (
            .O(N__24409),
            .I(N__24378));
    InMux I__5184 (
            .O(N__24408),
            .I(N__24378));
    LocalMux I__5183 (
            .O(N__24401),
            .I(N__24373));
    LocalMux I__5182 (
            .O(N__24398),
            .I(N__24373));
    LocalMux I__5181 (
            .O(N__24393),
            .I(\eeprom.n2539 ));
    LocalMux I__5180 (
            .O(N__24386),
            .I(\eeprom.n2539 ));
    Odrv4 I__5179 (
            .O(N__24383),
            .I(\eeprom.n2539 ));
    LocalMux I__5178 (
            .O(N__24378),
            .I(\eeprom.n2539 ));
    Odrv4 I__5177 (
            .O(N__24373),
            .I(\eeprom.n2539 ));
    CascadeMux I__5176 (
            .O(N__24362),
            .I(N__24359));
    InMux I__5175 (
            .O(N__24359),
            .I(N__24356));
    LocalMux I__5174 (
            .O(N__24356),
            .I(N__24352));
    CascadeMux I__5173 (
            .O(N__24355),
            .I(N__24349));
    Span4Mux_v I__5172 (
            .O(N__24352),
            .I(N__24346));
    InMux I__5171 (
            .O(N__24349),
            .I(N__24343));
    Odrv4 I__5170 (
            .O(N__24346),
            .I(\eeprom.n2506 ));
    LocalMux I__5169 (
            .O(N__24343),
            .I(\eeprom.n2506 ));
    InMux I__5168 (
            .O(N__24338),
            .I(\eeprom.n4042 ));
    InMux I__5167 (
            .O(N__24335),
            .I(N__24332));
    LocalMux I__5166 (
            .O(N__24332),
            .I(N__24328));
    InMux I__5165 (
            .O(N__24331),
            .I(N__24325));
    Odrv4 I__5164 (
            .O(N__24328),
            .I(\eeprom.n2605 ));
    LocalMux I__5163 (
            .O(N__24325),
            .I(\eeprom.n2605 ));
    InMux I__5162 (
            .O(N__24320),
            .I(N__24316));
    InMux I__5161 (
            .O(N__24319),
            .I(N__24313));
    LocalMux I__5160 (
            .O(N__24316),
            .I(N__24309));
    LocalMux I__5159 (
            .O(N__24313),
            .I(N__24306));
    CascadeMux I__5158 (
            .O(N__24312),
            .I(N__24303));
    Span4Mux_h I__5157 (
            .O(N__24309),
            .I(N__24300));
    Span4Mux_h I__5156 (
            .O(N__24306),
            .I(N__24297));
    InMux I__5155 (
            .O(N__24303),
            .I(N__24294));
    Odrv4 I__5154 (
            .O(N__24300),
            .I(\eeprom.n2519 ));
    Odrv4 I__5153 (
            .O(N__24297),
            .I(\eeprom.n2519 ));
    LocalMux I__5152 (
            .O(N__24294),
            .I(\eeprom.n2519 ));
    InMux I__5151 (
            .O(N__24287),
            .I(N__24283));
    InMux I__5150 (
            .O(N__24286),
            .I(N__24279));
    LocalMux I__5149 (
            .O(N__24283),
            .I(N__24276));
    InMux I__5148 (
            .O(N__24282),
            .I(N__24273));
    LocalMux I__5147 (
            .O(N__24279),
            .I(N__24270));
    Span4Mux_v I__5146 (
            .O(N__24276),
            .I(N__24267));
    LocalMux I__5145 (
            .O(N__24273),
            .I(N__24262));
    Span4Mux_v I__5144 (
            .O(N__24270),
            .I(N__24262));
    Odrv4 I__5143 (
            .O(N__24267),
            .I(\eeprom.n2619 ));
    Odrv4 I__5142 (
            .O(N__24262),
            .I(\eeprom.n2619 ));
    InMux I__5141 (
            .O(N__24257),
            .I(N__24250));
    InMux I__5140 (
            .O(N__24256),
            .I(N__24250));
    InMux I__5139 (
            .O(N__24255),
            .I(N__24247));
    LocalMux I__5138 (
            .O(N__24250),
            .I(N__24242));
    LocalMux I__5137 (
            .O(N__24247),
            .I(N__24242));
    Span4Mux_v I__5136 (
            .O(N__24242),
            .I(N__24239));
    Odrv4 I__5135 (
            .O(N__24239),
            .I(\eeprom.n2819 ));
    InMux I__5134 (
            .O(N__24236),
            .I(N__24232));
    InMux I__5133 (
            .O(N__24235),
            .I(N__24228));
    LocalMux I__5132 (
            .O(N__24232),
            .I(N__24225));
    InMux I__5131 (
            .O(N__24231),
            .I(N__24222));
    LocalMux I__5130 (
            .O(N__24228),
            .I(N__24219));
    Span4Mux_v I__5129 (
            .O(N__24225),
            .I(N__24214));
    LocalMux I__5128 (
            .O(N__24222),
            .I(N__24214));
    Span4Mux_h I__5127 (
            .O(N__24219),
            .I(N__24211));
    Span4Mux_h I__5126 (
            .O(N__24214),
            .I(N__24208));
    Span4Mux_h I__5125 (
            .O(N__24211),
            .I(N__24205));
    Span4Mux_h I__5124 (
            .O(N__24208),
            .I(N__24202));
    Odrv4 I__5123 (
            .O(N__24205),
            .I(\eeprom.n3219 ));
    Odrv4 I__5122 (
            .O(N__24202),
            .I(\eeprom.n3219 ));
    InMux I__5121 (
            .O(N__24197),
            .I(N__24193));
    InMux I__5120 (
            .O(N__24196),
            .I(N__24190));
    LocalMux I__5119 (
            .O(N__24193),
            .I(N__24184));
    LocalMux I__5118 (
            .O(N__24190),
            .I(N__24184));
    InMux I__5117 (
            .O(N__24189),
            .I(N__24181));
    Span4Mux_h I__5116 (
            .O(N__24184),
            .I(N__24178));
    LocalMux I__5115 (
            .O(N__24181),
            .I(N__24175));
    Span4Mux_h I__5114 (
            .O(N__24178),
            .I(N__24172));
    Odrv12 I__5113 (
            .O(N__24175),
            .I(\eeprom.n3019 ));
    Odrv4 I__5112 (
            .O(N__24172),
            .I(\eeprom.n3019 ));
    CascadeMux I__5111 (
            .O(N__24167),
            .I(N__24164));
    InMux I__5110 (
            .O(N__24164),
            .I(N__24159));
    InMux I__5109 (
            .O(N__24163),
            .I(N__24156));
    InMux I__5108 (
            .O(N__24162),
            .I(N__24153));
    LocalMux I__5107 (
            .O(N__24159),
            .I(N__24150));
    LocalMux I__5106 (
            .O(N__24156),
            .I(\eeprom.n2516 ));
    LocalMux I__5105 (
            .O(N__24153),
            .I(\eeprom.n2516 ));
    Odrv4 I__5104 (
            .O(N__24150),
            .I(\eeprom.n2516 ));
    InMux I__5103 (
            .O(N__24143),
            .I(N__24140));
    LocalMux I__5102 (
            .O(N__24140),
            .I(\eeprom.n2583 ));
    InMux I__5101 (
            .O(N__24137),
            .I(\eeprom.n4032 ));
    CascadeMux I__5100 (
            .O(N__24134),
            .I(N__24131));
    InMux I__5099 (
            .O(N__24131),
            .I(N__24126));
    CascadeMux I__5098 (
            .O(N__24130),
            .I(N__24123));
    InMux I__5097 (
            .O(N__24129),
            .I(N__24120));
    LocalMux I__5096 (
            .O(N__24126),
            .I(N__24117));
    InMux I__5095 (
            .O(N__24123),
            .I(N__24114));
    LocalMux I__5094 (
            .O(N__24120),
            .I(\eeprom.n2515 ));
    Odrv4 I__5093 (
            .O(N__24117),
            .I(\eeprom.n2515 ));
    LocalMux I__5092 (
            .O(N__24114),
            .I(\eeprom.n2515 ));
    InMux I__5091 (
            .O(N__24107),
            .I(N__24104));
    LocalMux I__5090 (
            .O(N__24104),
            .I(\eeprom.n2582 ));
    InMux I__5089 (
            .O(N__24101),
            .I(\eeprom.n4033 ));
    CascadeMux I__5088 (
            .O(N__24098),
            .I(N__24095));
    InMux I__5087 (
            .O(N__24095),
            .I(N__24090));
    InMux I__5086 (
            .O(N__24094),
            .I(N__24087));
    InMux I__5085 (
            .O(N__24093),
            .I(N__24084));
    LocalMux I__5084 (
            .O(N__24090),
            .I(N__24081));
    LocalMux I__5083 (
            .O(N__24087),
            .I(\eeprom.n2514 ));
    LocalMux I__5082 (
            .O(N__24084),
            .I(\eeprom.n2514 ));
    Odrv4 I__5081 (
            .O(N__24081),
            .I(\eeprom.n2514 ));
    InMux I__5080 (
            .O(N__24074),
            .I(N__24071));
    LocalMux I__5079 (
            .O(N__24071),
            .I(\eeprom.n2581 ));
    InMux I__5078 (
            .O(N__24068),
            .I(\eeprom.n4034 ));
    CascadeMux I__5077 (
            .O(N__24065),
            .I(N__24062));
    InMux I__5076 (
            .O(N__24062),
            .I(N__24058));
    InMux I__5075 (
            .O(N__24061),
            .I(N__24054));
    LocalMux I__5074 (
            .O(N__24058),
            .I(N__24051));
    InMux I__5073 (
            .O(N__24057),
            .I(N__24048));
    LocalMux I__5072 (
            .O(N__24054),
            .I(N__24043));
    Span4Mux_h I__5071 (
            .O(N__24051),
            .I(N__24043));
    LocalMux I__5070 (
            .O(N__24048),
            .I(N__24040));
    Odrv4 I__5069 (
            .O(N__24043),
            .I(\eeprom.n2513 ));
    Odrv4 I__5068 (
            .O(N__24040),
            .I(\eeprom.n2513 ));
    InMux I__5067 (
            .O(N__24035),
            .I(N__24032));
    LocalMux I__5066 (
            .O(N__24032),
            .I(\eeprom.n2580 ));
    InMux I__5065 (
            .O(N__24029),
            .I(\eeprom.n4035 ));
    CascadeMux I__5064 (
            .O(N__24026),
            .I(N__24023));
    InMux I__5063 (
            .O(N__24023),
            .I(N__24020));
    LocalMux I__5062 (
            .O(N__24020),
            .I(N__24015));
    InMux I__5061 (
            .O(N__24019),
            .I(N__24010));
    InMux I__5060 (
            .O(N__24018),
            .I(N__24010));
    Span4Mux_h I__5059 (
            .O(N__24015),
            .I(N__24007));
    LocalMux I__5058 (
            .O(N__24010),
            .I(\eeprom.n2512 ));
    Odrv4 I__5057 (
            .O(N__24007),
            .I(\eeprom.n2512 ));
    InMux I__5056 (
            .O(N__24002),
            .I(N__23999));
    LocalMux I__5055 (
            .O(N__23999),
            .I(\eeprom.n2579 ));
    InMux I__5054 (
            .O(N__23996),
            .I(\eeprom.n4036 ));
    CascadeMux I__5053 (
            .O(N__23993),
            .I(N__23990));
    InMux I__5052 (
            .O(N__23990),
            .I(N__23986));
    InMux I__5051 (
            .O(N__23989),
            .I(N__23983));
    LocalMux I__5050 (
            .O(N__23986),
            .I(N__23980));
    LocalMux I__5049 (
            .O(N__23983),
            .I(N__23977));
    Span4Mux_h I__5048 (
            .O(N__23980),
            .I(N__23974));
    Odrv4 I__5047 (
            .O(N__23977),
            .I(\eeprom.n2511 ));
    Odrv4 I__5046 (
            .O(N__23974),
            .I(\eeprom.n2511 ));
    InMux I__5045 (
            .O(N__23969),
            .I(N__23966));
    LocalMux I__5044 (
            .O(N__23966),
            .I(N__23963));
    Span4Mux_h I__5043 (
            .O(N__23963),
            .I(N__23960));
    Odrv4 I__5042 (
            .O(N__23960),
            .I(\eeprom.n2578 ));
    InMux I__5041 (
            .O(N__23957),
            .I(bfn_24_24_0_));
    CascadeMux I__5040 (
            .O(N__23954),
            .I(N__23951));
    InMux I__5039 (
            .O(N__23951),
            .I(N__23948));
    LocalMux I__5038 (
            .O(N__23948),
            .I(N__23944));
    InMux I__5037 (
            .O(N__23947),
            .I(N__23941));
    Sp12to4 I__5036 (
            .O(N__23944),
            .I(N__23935));
    LocalMux I__5035 (
            .O(N__23941),
            .I(N__23935));
    InMux I__5034 (
            .O(N__23940),
            .I(N__23932));
    Odrv12 I__5033 (
            .O(N__23935),
            .I(\eeprom.n2510 ));
    LocalMux I__5032 (
            .O(N__23932),
            .I(\eeprom.n2510 ));
    InMux I__5031 (
            .O(N__23927),
            .I(N__23924));
    LocalMux I__5030 (
            .O(N__23924),
            .I(\eeprom.n2577 ));
    InMux I__5029 (
            .O(N__23921),
            .I(\eeprom.n4038 ));
    CascadeMux I__5028 (
            .O(N__23918),
            .I(N__23914));
    InMux I__5027 (
            .O(N__23917),
            .I(N__23911));
    InMux I__5026 (
            .O(N__23914),
            .I(N__23908));
    LocalMux I__5025 (
            .O(N__23911),
            .I(N__23902));
    LocalMux I__5024 (
            .O(N__23908),
            .I(N__23902));
    InMux I__5023 (
            .O(N__23907),
            .I(N__23899));
    Odrv4 I__5022 (
            .O(N__23902),
            .I(\eeprom.n2509 ));
    LocalMux I__5021 (
            .O(N__23899),
            .I(\eeprom.n2509 ));
    InMux I__5020 (
            .O(N__23894),
            .I(N__23891));
    LocalMux I__5019 (
            .O(N__23891),
            .I(\eeprom.n2576 ));
    InMux I__5018 (
            .O(N__23888),
            .I(\eeprom.n4039 ));
    CascadeMux I__5017 (
            .O(N__23885),
            .I(\eeprom.n5173_cascade_ ));
    InMux I__5016 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__5015 (
            .O(N__23879),
            .I(\eeprom.n11_adj_328 ));
    CascadeMux I__5014 (
            .O(N__23876),
            .I(N__23872));
    CascadeMux I__5013 (
            .O(N__23875),
            .I(N__23869));
    InMux I__5012 (
            .O(N__23872),
            .I(N__23866));
    InMux I__5011 (
            .O(N__23869),
            .I(N__23863));
    LocalMux I__5010 (
            .O(N__23866),
            .I(N__23860));
    LocalMux I__5009 (
            .O(N__23863),
            .I(N__23857));
    Span4Mux_v I__5008 (
            .O(N__23860),
            .I(N__23854));
    Odrv4 I__5007 (
            .O(N__23857),
            .I(\eeprom.n2615 ));
    Odrv4 I__5006 (
            .O(N__23854),
            .I(\eeprom.n2615 ));
    CascadeMux I__5005 (
            .O(N__23849),
            .I(\eeprom.n2615_cascade_ ));
    CascadeMux I__5004 (
            .O(N__23846),
            .I(N__23843));
    InMux I__5003 (
            .O(N__23843),
            .I(N__23839));
    InMux I__5002 (
            .O(N__23842),
            .I(N__23836));
    LocalMux I__5001 (
            .O(N__23839),
            .I(N__23833));
    LocalMux I__5000 (
            .O(N__23836),
            .I(N__23829));
    Span4Mux_v I__4999 (
            .O(N__23833),
            .I(N__23826));
    InMux I__4998 (
            .O(N__23832),
            .I(N__23823));
    Odrv4 I__4997 (
            .O(N__23829),
            .I(\eeprom.n2613 ));
    Odrv4 I__4996 (
            .O(N__23826),
            .I(\eeprom.n2613 ));
    LocalMux I__4995 (
            .O(N__23823),
            .I(\eeprom.n2613 ));
    CascadeMux I__4994 (
            .O(N__23816),
            .I(N__23813));
    InMux I__4993 (
            .O(N__23813),
            .I(N__23810));
    LocalMux I__4992 (
            .O(N__23810),
            .I(N__23806));
    InMux I__4991 (
            .O(N__23809),
            .I(N__23802));
    Span4Mux_h I__4990 (
            .O(N__23806),
            .I(N__23799));
    InMux I__4989 (
            .O(N__23805),
            .I(N__23796));
    LocalMux I__4988 (
            .O(N__23802),
            .I(\eeprom.n2617 ));
    Odrv4 I__4987 (
            .O(N__23799),
            .I(\eeprom.n2617 ));
    LocalMux I__4986 (
            .O(N__23796),
            .I(\eeprom.n2617 ));
    CascadeMux I__4985 (
            .O(N__23789),
            .I(N__23786));
    InMux I__4984 (
            .O(N__23786),
            .I(N__23783));
    LocalMux I__4983 (
            .O(N__23783),
            .I(N__23779));
    InMux I__4982 (
            .O(N__23782),
            .I(N__23775));
    Span4Mux_h I__4981 (
            .O(N__23779),
            .I(N__23772));
    InMux I__4980 (
            .O(N__23778),
            .I(N__23769));
    LocalMux I__4979 (
            .O(N__23775),
            .I(\eeprom.n2614 ));
    Odrv4 I__4978 (
            .O(N__23772),
            .I(\eeprom.n2614 ));
    LocalMux I__4977 (
            .O(N__23769),
            .I(\eeprom.n2614 ));
    CascadeMux I__4976 (
            .O(N__23762),
            .I(\eeprom.n5101_cascade_ ));
    CascadeMux I__4975 (
            .O(N__23759),
            .I(N__23756));
    InMux I__4974 (
            .O(N__23756),
            .I(N__23753));
    LocalMux I__4973 (
            .O(N__23753),
            .I(N__23749));
    InMux I__4972 (
            .O(N__23752),
            .I(N__23745));
    Span4Mux_h I__4971 (
            .O(N__23749),
            .I(N__23742));
    InMux I__4970 (
            .O(N__23748),
            .I(N__23739));
    LocalMux I__4969 (
            .O(N__23745),
            .I(\eeprom.n2616 ));
    Odrv4 I__4968 (
            .O(N__23742),
            .I(\eeprom.n2616 ));
    LocalMux I__4967 (
            .O(N__23739),
            .I(\eeprom.n2616 ));
    CascadeMux I__4966 (
            .O(N__23732),
            .I(N__23729));
    InMux I__4965 (
            .O(N__23729),
            .I(N__23726));
    LocalMux I__4964 (
            .O(N__23726),
            .I(\eeprom.n5105 ));
    InMux I__4963 (
            .O(N__23723),
            .I(N__23720));
    LocalMux I__4962 (
            .O(N__23720),
            .I(N__23717));
    Span4Mux_v I__4961 (
            .O(N__23717),
            .I(N__23714));
    Odrv4 I__4960 (
            .O(N__23714),
            .I(\eeprom.n2586 ));
    InMux I__4959 (
            .O(N__23711),
            .I(bfn_24_23_0_));
    CascadeMux I__4958 (
            .O(N__23708),
            .I(N__23704));
    CascadeMux I__4957 (
            .O(N__23707),
            .I(N__23701));
    InMux I__4956 (
            .O(N__23704),
            .I(N__23697));
    InMux I__4955 (
            .O(N__23701),
            .I(N__23694));
    InMux I__4954 (
            .O(N__23700),
            .I(N__23691));
    LocalMux I__4953 (
            .O(N__23697),
            .I(N__23688));
    LocalMux I__4952 (
            .O(N__23694),
            .I(\eeprom.n2518 ));
    LocalMux I__4951 (
            .O(N__23691),
            .I(\eeprom.n2518 ));
    Odrv4 I__4950 (
            .O(N__23688),
            .I(\eeprom.n2518 ));
    InMux I__4949 (
            .O(N__23681),
            .I(N__23678));
    LocalMux I__4948 (
            .O(N__23678),
            .I(\eeprom.n2585 ));
    InMux I__4947 (
            .O(N__23675),
            .I(\eeprom.n4030 ));
    CascadeMux I__4946 (
            .O(N__23672),
            .I(N__23668));
    CascadeMux I__4945 (
            .O(N__23671),
            .I(N__23665));
    InMux I__4944 (
            .O(N__23668),
            .I(N__23661));
    InMux I__4943 (
            .O(N__23665),
            .I(N__23658));
    InMux I__4942 (
            .O(N__23664),
            .I(N__23655));
    LocalMux I__4941 (
            .O(N__23661),
            .I(N__23652));
    LocalMux I__4940 (
            .O(N__23658),
            .I(\eeprom.n2517 ));
    LocalMux I__4939 (
            .O(N__23655),
            .I(\eeprom.n2517 ));
    Odrv4 I__4938 (
            .O(N__23652),
            .I(\eeprom.n2517 ));
    InMux I__4937 (
            .O(N__23645),
            .I(N__23642));
    LocalMux I__4936 (
            .O(N__23642),
            .I(\eeprom.n2584 ));
    InMux I__4935 (
            .O(N__23639),
            .I(\eeprom.n4031 ));
    InMux I__4934 (
            .O(N__23636),
            .I(N__23633));
    LocalMux I__4933 (
            .O(N__23633),
            .I(\eeprom.n1982 ));
    InMux I__4932 (
            .O(N__23630),
            .I(\eeprom.n3976 ));
    InMux I__4931 (
            .O(N__23627),
            .I(N__23624));
    LocalMux I__4930 (
            .O(N__23624),
            .I(\eeprom.n1981 ));
    InMux I__4929 (
            .O(N__23621),
            .I(\eeprom.n3977 ));
    CascadeMux I__4928 (
            .O(N__23618),
            .I(N__23615));
    InMux I__4927 (
            .O(N__23615),
            .I(N__23612));
    LocalMux I__4926 (
            .O(N__23612),
            .I(\eeprom.n1980 ));
    InMux I__4925 (
            .O(N__23609),
            .I(\eeprom.n3978 ));
    CascadeMux I__4924 (
            .O(N__23606),
            .I(N__23600));
    CascadeMux I__4923 (
            .O(N__23605),
            .I(N__23597));
    CascadeMux I__4922 (
            .O(N__23604),
            .I(N__23593));
    CascadeMux I__4921 (
            .O(N__23603),
            .I(N__23589));
    InMux I__4920 (
            .O(N__23600),
            .I(N__23585));
    InMux I__4919 (
            .O(N__23597),
            .I(N__23580));
    InMux I__4918 (
            .O(N__23596),
            .I(N__23580));
    InMux I__4917 (
            .O(N__23593),
            .I(N__23571));
    InMux I__4916 (
            .O(N__23592),
            .I(N__23571));
    InMux I__4915 (
            .O(N__23589),
            .I(N__23571));
    InMux I__4914 (
            .O(N__23588),
            .I(N__23571));
    LocalMux I__4913 (
            .O(N__23585),
            .I(\eeprom.n1945 ));
    LocalMux I__4912 (
            .O(N__23580),
            .I(\eeprom.n1945 ));
    LocalMux I__4911 (
            .O(N__23571),
            .I(\eeprom.n1945 ));
    InMux I__4910 (
            .O(N__23564),
            .I(\eeprom.n3979 ));
    InMux I__4909 (
            .O(N__23561),
            .I(N__23557));
    CascadeMux I__4908 (
            .O(N__23560),
            .I(N__23554));
    LocalMux I__4907 (
            .O(N__23557),
            .I(N__23551));
    InMux I__4906 (
            .O(N__23554),
            .I(N__23548));
    Span4Mux_h I__4905 (
            .O(N__23551),
            .I(N__23545));
    LocalMux I__4904 (
            .O(N__23548),
            .I(\eeprom.n2011 ));
    Odrv4 I__4903 (
            .O(N__23545),
            .I(\eeprom.n2011 ));
    InMux I__4902 (
            .O(N__23540),
            .I(N__23536));
    CascadeMux I__4901 (
            .O(N__23539),
            .I(N__23533));
    LocalMux I__4900 (
            .O(N__23536),
            .I(N__23530));
    InMux I__4899 (
            .O(N__23533),
            .I(N__23527));
    Span4Mux_h I__4898 (
            .O(N__23530),
            .I(N__23523));
    LocalMux I__4897 (
            .O(N__23527),
            .I(N__23520));
    InMux I__4896 (
            .O(N__23526),
            .I(N__23517));
    Odrv4 I__4895 (
            .O(N__23523),
            .I(\eeprom.n2411 ));
    Odrv4 I__4894 (
            .O(N__23520),
            .I(\eeprom.n2411 ));
    LocalMux I__4893 (
            .O(N__23517),
            .I(\eeprom.n2411 ));
    CascadeMux I__4892 (
            .O(N__23510),
            .I(N__23507));
    InMux I__4891 (
            .O(N__23507),
            .I(N__23504));
    LocalMux I__4890 (
            .O(N__23504),
            .I(N__23501));
    Span4Mux_h I__4889 (
            .O(N__23501),
            .I(N__23498));
    Odrv4 I__4888 (
            .O(N__23498),
            .I(\eeprom.n2478 ));
    InMux I__4887 (
            .O(N__23495),
            .I(N__23487));
    InMux I__4886 (
            .O(N__23494),
            .I(N__23483));
    CascadeMux I__4885 (
            .O(N__23493),
            .I(N__23480));
    CascadeMux I__4884 (
            .O(N__23492),
            .I(N__23476));
    CascadeMux I__4883 (
            .O(N__23491),
            .I(N__23471));
    CascadeMux I__4882 (
            .O(N__23490),
            .I(N__23468));
    LocalMux I__4881 (
            .O(N__23487),
            .I(N__23463));
    InMux I__4880 (
            .O(N__23486),
            .I(N__23460));
    LocalMux I__4879 (
            .O(N__23483),
            .I(N__23457));
    InMux I__4878 (
            .O(N__23480),
            .I(N__23452));
    InMux I__4877 (
            .O(N__23479),
            .I(N__23452));
    InMux I__4876 (
            .O(N__23476),
            .I(N__23437));
    InMux I__4875 (
            .O(N__23475),
            .I(N__23437));
    InMux I__4874 (
            .O(N__23474),
            .I(N__23437));
    InMux I__4873 (
            .O(N__23471),
            .I(N__23437));
    InMux I__4872 (
            .O(N__23468),
            .I(N__23437));
    InMux I__4871 (
            .O(N__23467),
            .I(N__23437));
    InMux I__4870 (
            .O(N__23466),
            .I(N__23437));
    Odrv4 I__4869 (
            .O(N__23463),
            .I(\eeprom.n2440 ));
    LocalMux I__4868 (
            .O(N__23460),
            .I(\eeprom.n2440 ));
    Odrv4 I__4867 (
            .O(N__23457),
            .I(\eeprom.n2440 ));
    LocalMux I__4866 (
            .O(N__23452),
            .I(\eeprom.n2440 ));
    LocalMux I__4865 (
            .O(N__23437),
            .I(\eeprom.n2440 ));
    InMux I__4864 (
            .O(N__23426),
            .I(N__23423));
    LocalMux I__4863 (
            .O(N__23423),
            .I(N__23418));
    InMux I__4862 (
            .O(N__23422),
            .I(N__23415));
    InMux I__4861 (
            .O(N__23421),
            .I(N__23412));
    Span4Mux_v I__4860 (
            .O(N__23418),
            .I(N__23407));
    LocalMux I__4859 (
            .O(N__23415),
            .I(N__23407));
    LocalMux I__4858 (
            .O(N__23412),
            .I(N__23404));
    Span4Mux_h I__4857 (
            .O(N__23407),
            .I(N__23401));
    Odrv12 I__4856 (
            .O(N__23404),
            .I(\eeprom.n3419 ));
    Odrv4 I__4855 (
            .O(N__23401),
            .I(\eeprom.n3419 ));
    CascadeMux I__4854 (
            .O(N__23396),
            .I(\eeprom.n5169_cascade_ ));
    CascadeMux I__4853 (
            .O(N__23393),
            .I(N__23389));
    InMux I__4852 (
            .O(N__23392),
            .I(N__23386));
    InMux I__4851 (
            .O(N__23389),
            .I(N__23383));
    LocalMux I__4850 (
            .O(N__23386),
            .I(N__23380));
    LocalMux I__4849 (
            .O(N__23383),
            .I(\eeprom.n2016 ));
    Odrv4 I__4848 (
            .O(N__23380),
            .I(\eeprom.n2016 ));
    InMux I__4847 (
            .O(N__23375),
            .I(N__23372));
    LocalMux I__4846 (
            .O(N__23372),
            .I(\eeprom.n2083 ));
    CascadeMux I__4845 (
            .O(N__23369),
            .I(\eeprom.n2016_cascade_ ));
    CascadeMux I__4844 (
            .O(N__23366),
            .I(N__23360));
    InMux I__4843 (
            .O(N__23365),
            .I(N__23354));
    InMux I__4842 (
            .O(N__23364),
            .I(N__23345));
    InMux I__4841 (
            .O(N__23363),
            .I(N__23345));
    InMux I__4840 (
            .O(N__23360),
            .I(N__23345));
    InMux I__4839 (
            .O(N__23359),
            .I(N__23345));
    CascadeMux I__4838 (
            .O(N__23358),
            .I(N__23342));
    InMux I__4837 (
            .O(N__23357),
            .I(N__23337));
    LocalMux I__4836 (
            .O(N__23354),
            .I(N__23334));
    LocalMux I__4835 (
            .O(N__23345),
            .I(N__23331));
    InMux I__4834 (
            .O(N__23342),
            .I(N__23324));
    InMux I__4833 (
            .O(N__23341),
            .I(N__23324));
    InMux I__4832 (
            .O(N__23340),
            .I(N__23324));
    LocalMux I__4831 (
            .O(N__23337),
            .I(\eeprom.n2044 ));
    Odrv4 I__4830 (
            .O(N__23334),
            .I(\eeprom.n2044 ));
    Odrv4 I__4829 (
            .O(N__23331),
            .I(\eeprom.n2044 ));
    LocalMux I__4828 (
            .O(N__23324),
            .I(\eeprom.n2044 ));
    CascadeMux I__4827 (
            .O(N__23315),
            .I(N__23311));
    CascadeMux I__4826 (
            .O(N__23314),
            .I(N__23308));
    InMux I__4825 (
            .O(N__23311),
            .I(N__23305));
    InMux I__4824 (
            .O(N__23308),
            .I(N__23302));
    LocalMux I__4823 (
            .O(N__23305),
            .I(N__23299));
    LocalMux I__4822 (
            .O(N__23302),
            .I(N__23296));
    Odrv4 I__4821 (
            .O(N__23299),
            .I(\eeprom.n2115 ));
    Odrv4 I__4820 (
            .O(N__23296),
            .I(\eeprom.n2115 ));
    CascadeMux I__4819 (
            .O(N__23291),
            .I(\eeprom.n2115_cascade_ ));
    CascadeMux I__4818 (
            .O(N__23288),
            .I(N__23285));
    InMux I__4817 (
            .O(N__23285),
            .I(N__23281));
    InMux I__4816 (
            .O(N__23284),
            .I(N__23277));
    LocalMux I__4815 (
            .O(N__23281),
            .I(N__23274));
    InMux I__4814 (
            .O(N__23280),
            .I(N__23271));
    LocalMux I__4813 (
            .O(N__23277),
            .I(\eeprom.n2113 ));
    Odrv4 I__4812 (
            .O(N__23274),
            .I(\eeprom.n2113 ));
    LocalMux I__4811 (
            .O(N__23271),
            .I(\eeprom.n2113 ));
    InMux I__4810 (
            .O(N__23264),
            .I(N__23261));
    LocalMux I__4809 (
            .O(N__23261),
            .I(\eeprom.n5059 ));
    InMux I__4808 (
            .O(N__23258),
            .I(N__23253));
    InMux I__4807 (
            .O(N__23257),
            .I(N__23250));
    CascadeMux I__4806 (
            .O(N__23256),
            .I(N__23247));
    LocalMux I__4805 (
            .O(N__23253),
            .I(N__23242));
    LocalMux I__4804 (
            .O(N__23250),
            .I(N__23242));
    InMux I__4803 (
            .O(N__23247),
            .I(N__23239));
    Span4Mux_h I__4802 (
            .O(N__23242),
            .I(N__23236));
    LocalMux I__4801 (
            .O(N__23239),
            .I(\eeprom.n2013 ));
    Odrv4 I__4800 (
            .O(N__23236),
            .I(\eeprom.n2013 ));
    InMux I__4799 (
            .O(N__23231),
            .I(N__23226));
    InMux I__4798 (
            .O(N__23230),
            .I(N__23223));
    InMux I__4797 (
            .O(N__23229),
            .I(N__23220));
    LocalMux I__4796 (
            .O(N__23226),
            .I(N__23217));
    LocalMux I__4795 (
            .O(N__23223),
            .I(\eeprom.n2012 ));
    LocalMux I__4794 (
            .O(N__23220),
            .I(\eeprom.n2012 ));
    Odrv4 I__4793 (
            .O(N__23217),
            .I(\eeprom.n2012 ));
    InMux I__4792 (
            .O(N__23210),
            .I(N__23207));
    LocalMux I__4791 (
            .O(N__23207),
            .I(N__23204));
    Odrv4 I__4790 (
            .O(N__23204),
            .I(\eeprom.n1986 ));
    InMux I__4789 (
            .O(N__23201),
            .I(bfn_24_20_0_));
    InMux I__4788 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__4787 (
            .O(N__23195),
            .I(\eeprom.n1985 ));
    InMux I__4786 (
            .O(N__23192),
            .I(\eeprom.n3973 ));
    InMux I__4785 (
            .O(N__23189),
            .I(N__23186));
    LocalMux I__4784 (
            .O(N__23186),
            .I(\eeprom.n1984 ));
    InMux I__4783 (
            .O(N__23183),
            .I(\eeprom.n3974 ));
    InMux I__4782 (
            .O(N__23180),
            .I(N__23177));
    LocalMux I__4781 (
            .O(N__23177),
            .I(N__23174));
    Odrv4 I__4780 (
            .O(N__23174),
            .I(\eeprom.n1983 ));
    InMux I__4779 (
            .O(N__23171),
            .I(\eeprom.n3975 ));
    InMux I__4778 (
            .O(N__23168),
            .I(N__23164));
    InMux I__4777 (
            .O(N__23167),
            .I(N__23161));
    LocalMux I__4776 (
            .O(N__23164),
            .I(\eeprom.n2110 ));
    LocalMux I__4775 (
            .O(N__23161),
            .I(\eeprom.n2110 ));
    CascadeMux I__4774 (
            .O(N__23156),
            .I(N__23151));
    CascadeMux I__4773 (
            .O(N__23155),
            .I(N__23148));
    CascadeMux I__4772 (
            .O(N__23154),
            .I(N__23141));
    InMux I__4771 (
            .O(N__23151),
            .I(N__23134));
    InMux I__4770 (
            .O(N__23148),
            .I(N__23131));
    InMux I__4769 (
            .O(N__23147),
            .I(N__23128));
    InMux I__4768 (
            .O(N__23146),
            .I(N__23121));
    InMux I__4767 (
            .O(N__23145),
            .I(N__23121));
    InMux I__4766 (
            .O(N__23144),
            .I(N__23121));
    InMux I__4765 (
            .O(N__23141),
            .I(N__23116));
    InMux I__4764 (
            .O(N__23140),
            .I(N__23116));
    InMux I__4763 (
            .O(N__23139),
            .I(N__23109));
    InMux I__4762 (
            .O(N__23138),
            .I(N__23109));
    InMux I__4761 (
            .O(N__23137),
            .I(N__23109));
    LocalMux I__4760 (
            .O(N__23134),
            .I(N__23106));
    LocalMux I__4759 (
            .O(N__23131),
            .I(\eeprom.n2143 ));
    LocalMux I__4758 (
            .O(N__23128),
            .I(\eeprom.n2143 ));
    LocalMux I__4757 (
            .O(N__23121),
            .I(\eeprom.n2143 ));
    LocalMux I__4756 (
            .O(N__23116),
            .I(\eeprom.n2143 ));
    LocalMux I__4755 (
            .O(N__23109),
            .I(\eeprom.n2143 ));
    Odrv4 I__4754 (
            .O(N__23106),
            .I(\eeprom.n2143 ));
    InMux I__4753 (
            .O(N__23093),
            .I(\eeprom.n3996 ));
    CascadeMux I__4752 (
            .O(N__23090),
            .I(N__23086));
    CascadeMux I__4751 (
            .O(N__23089),
            .I(N__23083));
    InMux I__4750 (
            .O(N__23086),
            .I(N__23080));
    InMux I__4749 (
            .O(N__23083),
            .I(N__23077));
    LocalMux I__4748 (
            .O(N__23080),
            .I(N__23074));
    LocalMux I__4747 (
            .O(N__23077),
            .I(N__23071));
    Odrv12 I__4746 (
            .O(N__23074),
            .I(\eeprom.n2209 ));
    Odrv4 I__4745 (
            .O(N__23071),
            .I(\eeprom.n2209 ));
    InMux I__4744 (
            .O(N__23066),
            .I(N__23063));
    LocalMux I__4743 (
            .O(N__23063),
            .I(N__23060));
    Span4Mux_v I__4742 (
            .O(N__23060),
            .I(N__23057));
    Odrv4 I__4741 (
            .O(N__23057),
            .I(\eeprom.n3724 ));
    CascadeMux I__4740 (
            .O(N__23054),
            .I(N__23051));
    InMux I__4739 (
            .O(N__23051),
            .I(N__23046));
    InMux I__4738 (
            .O(N__23050),
            .I(N__23041));
    InMux I__4737 (
            .O(N__23049),
            .I(N__23041));
    LocalMux I__4736 (
            .O(N__23046),
            .I(\eeprom.n2015 ));
    LocalMux I__4735 (
            .O(N__23041),
            .I(\eeprom.n2015 ));
    CascadeMux I__4734 (
            .O(N__23036),
            .I(N__23033));
    InMux I__4733 (
            .O(N__23033),
            .I(N__23030));
    LocalMux I__4732 (
            .O(N__23030),
            .I(\eeprom.n2079 ));
    CascadeMux I__4731 (
            .O(N__23027),
            .I(N__23022));
    InMux I__4730 (
            .O(N__23026),
            .I(N__23019));
    InMux I__4729 (
            .O(N__23025),
            .I(N__23016));
    InMux I__4728 (
            .O(N__23022),
            .I(N__23013));
    LocalMux I__4727 (
            .O(N__23019),
            .I(N__23010));
    LocalMux I__4726 (
            .O(N__23016),
            .I(\eeprom.n2111 ));
    LocalMux I__4725 (
            .O(N__23013),
            .I(\eeprom.n2111 ));
    Odrv4 I__4724 (
            .O(N__23010),
            .I(\eeprom.n2111 ));
    CascadeMux I__4723 (
            .O(N__23003),
            .I(N__22999));
    CascadeMux I__4722 (
            .O(N__23002),
            .I(N__22995));
    InMux I__4721 (
            .O(N__22999),
            .I(N__22990));
    InMux I__4720 (
            .O(N__22998),
            .I(N__22990));
    InMux I__4719 (
            .O(N__22995),
            .I(N__22987));
    LocalMux I__4718 (
            .O(N__22990),
            .I(\eeprom.n2018 ));
    LocalMux I__4717 (
            .O(N__22987),
            .I(\eeprom.n2018 ));
    CascadeMux I__4716 (
            .O(N__22982),
            .I(\eeprom.n1945_cascade_ ));
    CascadeMux I__4715 (
            .O(N__22979),
            .I(N__22973));
    CascadeMux I__4714 (
            .O(N__22978),
            .I(N__22970));
    InMux I__4713 (
            .O(N__22977),
            .I(N__22967));
    CascadeMux I__4712 (
            .O(N__22976),
            .I(N__22964));
    InMux I__4711 (
            .O(N__22973),
            .I(N__22959));
    InMux I__4710 (
            .O(N__22970),
            .I(N__22959));
    LocalMux I__4709 (
            .O(N__22967),
            .I(N__22956));
    InMux I__4708 (
            .O(N__22964),
            .I(N__22953));
    LocalMux I__4707 (
            .O(N__22959),
            .I(N__22950));
    Odrv4 I__4706 (
            .O(N__22956),
            .I(\eeprom.n2017 ));
    LocalMux I__4705 (
            .O(N__22953),
            .I(\eeprom.n2017 ));
    Odrv4 I__4704 (
            .O(N__22950),
            .I(\eeprom.n2017 ));
    CascadeMux I__4703 (
            .O(N__22943),
            .I(N__22938));
    CascadeMux I__4702 (
            .O(N__22942),
            .I(N__22935));
    InMux I__4701 (
            .O(N__22941),
            .I(N__22932));
    InMux I__4700 (
            .O(N__22938),
            .I(N__22929));
    InMux I__4699 (
            .O(N__22935),
            .I(N__22926));
    LocalMux I__4698 (
            .O(N__22932),
            .I(N__22923));
    LocalMux I__4697 (
            .O(N__22929),
            .I(\eeprom.n2014 ));
    LocalMux I__4696 (
            .O(N__22926),
            .I(\eeprom.n2014 ));
    Odrv4 I__4695 (
            .O(N__22923),
            .I(\eeprom.n2014 ));
    CascadeMux I__4694 (
            .O(N__22916),
            .I(N__22913));
    InMux I__4693 (
            .O(N__22913),
            .I(N__22909));
    InMux I__4692 (
            .O(N__22912),
            .I(N__22906));
    LocalMux I__4691 (
            .O(N__22909),
            .I(N__22903));
    LocalMux I__4690 (
            .O(N__22906),
            .I(\eeprom.n2118 ));
    Odrv4 I__4689 (
            .O(N__22903),
            .I(\eeprom.n2118 ));
    InMux I__4688 (
            .O(N__22898),
            .I(N__22895));
    LocalMux I__4687 (
            .O(N__22895),
            .I(N__22892));
    Span4Mux_h I__4686 (
            .O(N__22892),
            .I(N__22889));
    Odrv4 I__4685 (
            .O(N__22889),
            .I(\eeprom.n2185 ));
    InMux I__4684 (
            .O(N__22886),
            .I(\eeprom.n3988 ));
    CascadeMux I__4683 (
            .O(N__22883),
            .I(N__22879));
    InMux I__4682 (
            .O(N__22882),
            .I(N__22875));
    InMux I__4681 (
            .O(N__22879),
            .I(N__22872));
    InMux I__4680 (
            .O(N__22878),
            .I(N__22869));
    LocalMux I__4679 (
            .O(N__22875),
            .I(\eeprom.n2117 ));
    LocalMux I__4678 (
            .O(N__22872),
            .I(\eeprom.n2117 ));
    LocalMux I__4677 (
            .O(N__22869),
            .I(\eeprom.n2117 ));
    CascadeMux I__4676 (
            .O(N__22862),
            .I(N__22859));
    InMux I__4675 (
            .O(N__22859),
            .I(N__22856));
    LocalMux I__4674 (
            .O(N__22856),
            .I(N__22853));
    Span4Mux_h I__4673 (
            .O(N__22853),
            .I(N__22850));
    Odrv4 I__4672 (
            .O(N__22850),
            .I(\eeprom.n2184 ));
    InMux I__4671 (
            .O(N__22847),
            .I(\eeprom.n3989 ));
    CascadeMux I__4670 (
            .O(N__22844),
            .I(N__22841));
    InMux I__4669 (
            .O(N__22841),
            .I(N__22838));
    LocalMux I__4668 (
            .O(N__22838),
            .I(N__22834));
    CascadeMux I__4667 (
            .O(N__22837),
            .I(N__22831));
    Span4Mux_v I__4666 (
            .O(N__22834),
            .I(N__22828));
    InMux I__4665 (
            .O(N__22831),
            .I(N__22825));
    Odrv4 I__4664 (
            .O(N__22828),
            .I(\eeprom.n2116 ));
    LocalMux I__4663 (
            .O(N__22825),
            .I(\eeprom.n2116 ));
    InMux I__4662 (
            .O(N__22820),
            .I(N__22816));
    InMux I__4661 (
            .O(N__22819),
            .I(N__22813));
    LocalMux I__4660 (
            .O(N__22816),
            .I(N__22810));
    LocalMux I__4659 (
            .O(N__22813),
            .I(N__22807));
    Span4Mux_v I__4658 (
            .O(N__22810),
            .I(N__22804));
    Span4Mux_h I__4657 (
            .O(N__22807),
            .I(N__22801));
    Odrv4 I__4656 (
            .O(N__22804),
            .I(\eeprom.n2183 ));
    Odrv4 I__4655 (
            .O(N__22801),
            .I(\eeprom.n2183 ));
    InMux I__4654 (
            .O(N__22796),
            .I(\eeprom.n3990 ));
    InMux I__4653 (
            .O(N__22793),
            .I(N__22790));
    LocalMux I__4652 (
            .O(N__22790),
            .I(N__22787));
    Span4Mux_h I__4651 (
            .O(N__22787),
            .I(N__22784));
    Odrv4 I__4650 (
            .O(N__22784),
            .I(\eeprom.n2182 ));
    InMux I__4649 (
            .O(N__22781),
            .I(\eeprom.n3991 ));
    CascadeMux I__4648 (
            .O(N__22778),
            .I(N__22774));
    InMux I__4647 (
            .O(N__22777),
            .I(N__22770));
    InMux I__4646 (
            .O(N__22774),
            .I(N__22767));
    InMux I__4645 (
            .O(N__22773),
            .I(N__22764));
    LocalMux I__4644 (
            .O(N__22770),
            .I(\eeprom.n2114 ));
    LocalMux I__4643 (
            .O(N__22767),
            .I(\eeprom.n2114 ));
    LocalMux I__4642 (
            .O(N__22764),
            .I(\eeprom.n2114 ));
    InMux I__4641 (
            .O(N__22757),
            .I(N__22754));
    LocalMux I__4640 (
            .O(N__22754),
            .I(N__22751));
    Span4Mux_v I__4639 (
            .O(N__22751),
            .I(N__22748));
    Odrv4 I__4638 (
            .O(N__22748),
            .I(\eeprom.n2181 ));
    InMux I__4637 (
            .O(N__22745),
            .I(\eeprom.n3992 ));
    InMux I__4636 (
            .O(N__22742),
            .I(N__22739));
    LocalMux I__4635 (
            .O(N__22739),
            .I(N__22736));
    Odrv4 I__4634 (
            .O(N__22736),
            .I(\eeprom.n2180 ));
    InMux I__4633 (
            .O(N__22733),
            .I(\eeprom.n3993 ));
    InMux I__4632 (
            .O(N__22730),
            .I(N__22727));
    LocalMux I__4631 (
            .O(N__22727),
            .I(N__22722));
    CascadeMux I__4630 (
            .O(N__22726),
            .I(N__22719));
    CascadeMux I__4629 (
            .O(N__22725),
            .I(N__22716));
    Span4Mux_h I__4628 (
            .O(N__22722),
            .I(N__22713));
    InMux I__4627 (
            .O(N__22719),
            .I(N__22710));
    InMux I__4626 (
            .O(N__22716),
            .I(N__22707));
    Odrv4 I__4625 (
            .O(N__22713),
            .I(\eeprom.n2112 ));
    LocalMux I__4624 (
            .O(N__22710),
            .I(\eeprom.n2112 ));
    LocalMux I__4623 (
            .O(N__22707),
            .I(\eeprom.n2112 ));
    CascadeMux I__4622 (
            .O(N__22700),
            .I(N__22697));
    InMux I__4621 (
            .O(N__22697),
            .I(N__22694));
    LocalMux I__4620 (
            .O(N__22694),
            .I(N__22691));
    Span4Mux_h I__4619 (
            .O(N__22691),
            .I(N__22688));
    Odrv4 I__4618 (
            .O(N__22688),
            .I(\eeprom.n2179 ));
    InMux I__4617 (
            .O(N__22685),
            .I(\eeprom.n3994 ));
    CascadeMux I__4616 (
            .O(N__22682),
            .I(N__22679));
    InMux I__4615 (
            .O(N__22679),
            .I(N__22676));
    LocalMux I__4614 (
            .O(N__22676),
            .I(\eeprom.n2178 ));
    InMux I__4613 (
            .O(N__22673),
            .I(bfn_24_18_0_));
    InMux I__4612 (
            .O(N__22670),
            .I(N__22667));
    LocalMux I__4611 (
            .O(N__22667),
            .I(N__22663));
    InMux I__4610 (
            .O(N__22666),
            .I(N__22660));
    Span4Mux_v I__4609 (
            .O(N__22663),
            .I(N__22654));
    LocalMux I__4608 (
            .O(N__22660),
            .I(N__22654));
    InMux I__4607 (
            .O(N__22659),
            .I(N__22651));
    Sp12to4 I__4606 (
            .O(N__22654),
            .I(N__22646));
    LocalMux I__4605 (
            .O(N__22651),
            .I(N__22646));
    Odrv12 I__4604 (
            .O(N__22646),
            .I(\eeprom.n3319 ));
    InMux I__4603 (
            .O(N__22643),
            .I(N__22639));
    InMux I__4602 (
            .O(N__22642),
            .I(N__22635));
    LocalMux I__4601 (
            .O(N__22639),
            .I(N__22632));
    InMux I__4600 (
            .O(N__22638),
            .I(N__22629));
    LocalMux I__4599 (
            .O(N__22635),
            .I(\eeprom.n2608 ));
    Odrv4 I__4598 (
            .O(N__22632),
            .I(\eeprom.n2608 ));
    LocalMux I__4597 (
            .O(N__22629),
            .I(\eeprom.n2608 ));
    CascadeMux I__4596 (
            .O(N__22622),
            .I(N__22619));
    InMux I__4595 (
            .O(N__22619),
            .I(N__22616));
    LocalMux I__4594 (
            .O(N__22616),
            .I(N__22612));
    InMux I__4593 (
            .O(N__22615),
            .I(N__22609));
    Odrv4 I__4592 (
            .O(N__22612),
            .I(\eeprom.n2607 ));
    LocalMux I__4591 (
            .O(N__22609),
            .I(\eeprom.n2607 ));
    InMux I__4590 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__4589 (
            .O(N__22601),
            .I(N__22598));
    Odrv4 I__4588 (
            .O(N__22598),
            .I(\eeprom.n2674 ));
    CascadeMux I__4587 (
            .O(N__22595),
            .I(\eeprom.n2607_cascade_ ));
    CascadeMux I__4586 (
            .O(N__22592),
            .I(N__22584));
    CascadeMux I__4585 (
            .O(N__22591),
            .I(N__22581));
    CascadeMux I__4584 (
            .O(N__22590),
            .I(N__22577));
    CascadeMux I__4583 (
            .O(N__22589),
            .I(N__22572));
    CascadeMux I__4582 (
            .O(N__22588),
            .I(N__22569));
    CascadeMux I__4581 (
            .O(N__22587),
            .I(N__22565));
    InMux I__4580 (
            .O(N__22584),
            .I(N__22556));
    InMux I__4579 (
            .O(N__22581),
            .I(N__22556));
    InMux I__4578 (
            .O(N__22580),
            .I(N__22551));
    InMux I__4577 (
            .O(N__22577),
            .I(N__22551));
    InMux I__4576 (
            .O(N__22576),
            .I(N__22540));
    InMux I__4575 (
            .O(N__22575),
            .I(N__22540));
    InMux I__4574 (
            .O(N__22572),
            .I(N__22540));
    InMux I__4573 (
            .O(N__22569),
            .I(N__22540));
    InMux I__4572 (
            .O(N__22568),
            .I(N__22540));
    InMux I__4571 (
            .O(N__22565),
            .I(N__22535));
    InMux I__4570 (
            .O(N__22564),
            .I(N__22535));
    InMux I__4569 (
            .O(N__22563),
            .I(N__22532));
    InMux I__4568 (
            .O(N__22562),
            .I(N__22527));
    InMux I__4567 (
            .O(N__22561),
            .I(N__22527));
    LocalMux I__4566 (
            .O(N__22556),
            .I(N__22524));
    LocalMux I__4565 (
            .O(N__22551),
            .I(\eeprom.n2638 ));
    LocalMux I__4564 (
            .O(N__22540),
            .I(\eeprom.n2638 ));
    LocalMux I__4563 (
            .O(N__22535),
            .I(\eeprom.n2638 ));
    LocalMux I__4562 (
            .O(N__22532),
            .I(\eeprom.n2638 ));
    LocalMux I__4561 (
            .O(N__22527),
            .I(\eeprom.n2638 ));
    Odrv4 I__4560 (
            .O(N__22524),
            .I(\eeprom.n2638 ));
    InMux I__4559 (
            .O(N__22511),
            .I(N__22507));
    InMux I__4558 (
            .O(N__22510),
            .I(N__22504));
    LocalMux I__4557 (
            .O(N__22507),
            .I(N__22501));
    LocalMux I__4556 (
            .O(N__22504),
            .I(N__22495));
    Span4Mux_h I__4555 (
            .O(N__22501),
            .I(N__22495));
    InMux I__4554 (
            .O(N__22500),
            .I(N__22492));
    Odrv4 I__4553 (
            .O(N__22495),
            .I(\eeprom.n2706 ));
    LocalMux I__4552 (
            .O(N__22492),
            .I(\eeprom.n2706 ));
    InMux I__4551 (
            .O(N__22487),
            .I(N__22482));
    InMux I__4550 (
            .O(N__22486),
            .I(N__22479));
    InMux I__4549 (
            .O(N__22485),
            .I(N__22476));
    LocalMux I__4548 (
            .O(N__22482),
            .I(N__22471));
    LocalMux I__4547 (
            .O(N__22479),
            .I(N__22471));
    LocalMux I__4546 (
            .O(N__22476),
            .I(\eeprom.n2719 ));
    Odrv4 I__4545 (
            .O(N__22471),
            .I(\eeprom.n2719 ));
    InMux I__4544 (
            .O(N__22466),
            .I(N__22461));
    InMux I__4543 (
            .O(N__22465),
            .I(N__22458));
    InMux I__4542 (
            .O(N__22464),
            .I(N__22455));
    LocalMux I__4541 (
            .O(N__22461),
            .I(N__22448));
    LocalMux I__4540 (
            .O(N__22458),
            .I(N__22448));
    LocalMux I__4539 (
            .O(N__22455),
            .I(N__22448));
    Span4Mux_v I__4538 (
            .O(N__22448),
            .I(N__22445));
    Odrv4 I__4537 (
            .O(N__22445),
            .I(\eeprom.n2919 ));
    InMux I__4536 (
            .O(N__22442),
            .I(N__22437));
    InMux I__4535 (
            .O(N__22441),
            .I(N__22434));
    CascadeMux I__4534 (
            .O(N__22440),
            .I(N__22431));
    LocalMux I__4533 (
            .O(N__22437),
            .I(N__22428));
    LocalMux I__4532 (
            .O(N__22434),
            .I(N__22425));
    InMux I__4531 (
            .O(N__22431),
            .I(N__22422));
    Span4Mux_h I__4530 (
            .O(N__22428),
            .I(N__22415));
    Span4Mux_h I__4529 (
            .O(N__22425),
            .I(N__22415));
    LocalMux I__4528 (
            .O(N__22422),
            .I(N__22415));
    Odrv4 I__4527 (
            .O(N__22415),
            .I(\eeprom.n2419 ));
    InMux I__4526 (
            .O(N__22412),
            .I(N__22408));
    InMux I__4525 (
            .O(N__22411),
            .I(N__22404));
    LocalMux I__4524 (
            .O(N__22408),
            .I(N__22401));
    InMux I__4523 (
            .O(N__22407),
            .I(N__22398));
    LocalMux I__4522 (
            .O(N__22404),
            .I(N__22395));
    Span4Mux_v I__4521 (
            .O(N__22401),
            .I(N__22392));
    LocalMux I__4520 (
            .O(N__22398),
            .I(N__22389));
    Span4Mux_h I__4519 (
            .O(N__22395),
            .I(N__22386));
    Span4Mux_h I__4518 (
            .O(N__22392),
            .I(N__22383));
    Span4Mux_h I__4517 (
            .O(N__22389),
            .I(N__22378));
    Span4Mux_v I__4516 (
            .O(N__22386),
            .I(N__22378));
    Odrv4 I__4515 (
            .O(N__22383),
            .I(\eeprom.n3119 ));
    Odrv4 I__4514 (
            .O(N__22378),
            .I(\eeprom.n3119 ));
    InMux I__4513 (
            .O(N__22373),
            .I(N__22370));
    LocalMux I__4512 (
            .O(N__22370),
            .I(N__22367));
    Span4Mux_h I__4511 (
            .O(N__22367),
            .I(N__22364));
    Odrv4 I__4510 (
            .O(N__22364),
            .I(\eeprom.n2186 ));
    InMux I__4509 (
            .O(N__22361),
            .I(bfn_24_17_0_));
    InMux I__4508 (
            .O(N__22358),
            .I(N__22354));
    InMux I__4507 (
            .O(N__22357),
            .I(N__22351));
    LocalMux I__4506 (
            .O(N__22354),
            .I(N__22348));
    LocalMux I__4505 (
            .O(N__22351),
            .I(\eeprom.n2612 ));
    Odrv4 I__4504 (
            .O(N__22348),
            .I(\eeprom.n2612 ));
    InMux I__4503 (
            .O(N__22343),
            .I(N__22339));
    InMux I__4502 (
            .O(N__22342),
            .I(N__22336));
    LocalMux I__4501 (
            .O(N__22339),
            .I(N__22333));
    LocalMux I__4500 (
            .O(N__22336),
            .I(N__22330));
    Span4Mux_v I__4499 (
            .O(N__22333),
            .I(N__22326));
    Span4Mux_h I__4498 (
            .O(N__22330),
            .I(N__22323));
    InMux I__4497 (
            .O(N__22329),
            .I(N__22320));
    Odrv4 I__4496 (
            .O(N__22326),
            .I(\eeprom.n2611 ));
    Odrv4 I__4495 (
            .O(N__22323),
            .I(\eeprom.n2611 ));
    LocalMux I__4494 (
            .O(N__22320),
            .I(\eeprom.n2611 ));
    CascadeMux I__4493 (
            .O(N__22313),
            .I(\eeprom.n2612_cascade_ ));
    CascadeMux I__4492 (
            .O(N__22310),
            .I(N__22305));
    CascadeMux I__4491 (
            .O(N__22309),
            .I(N__22302));
    InMux I__4490 (
            .O(N__22308),
            .I(N__22299));
    InMux I__4489 (
            .O(N__22305),
            .I(N__22294));
    InMux I__4488 (
            .O(N__22302),
            .I(N__22294));
    LocalMux I__4487 (
            .O(N__22299),
            .I(N__22291));
    LocalMux I__4486 (
            .O(N__22294),
            .I(N__22288));
    Span4Mux_h I__4485 (
            .O(N__22291),
            .I(N__22285));
    Odrv4 I__4484 (
            .O(N__22288),
            .I(\eeprom.n2610 ));
    Odrv4 I__4483 (
            .O(N__22285),
            .I(\eeprom.n2610 ));
    InMux I__4482 (
            .O(N__22280),
            .I(N__22277));
    LocalMux I__4481 (
            .O(N__22277),
            .I(\eeprom.n16_adj_334 ));
    InMux I__4480 (
            .O(N__22274),
            .I(N__22270));
    CascadeMux I__4479 (
            .O(N__22273),
            .I(N__22267));
    LocalMux I__4478 (
            .O(N__22270),
            .I(N__22264));
    InMux I__4477 (
            .O(N__22267),
            .I(N__22261));
    Span4Mux_v I__4476 (
            .O(N__22264),
            .I(N__22258));
    LocalMux I__4475 (
            .O(N__22261),
            .I(\eeprom.n2618 ));
    Odrv4 I__4474 (
            .O(N__22258),
            .I(\eeprom.n2618 ));
    CascadeMux I__4473 (
            .O(N__22253),
            .I(N__22250));
    InMux I__4472 (
            .O(N__22250),
            .I(N__22247));
    LocalMux I__4471 (
            .O(N__22247),
            .I(\eeprom.n12_adj_333 ));
    InMux I__4470 (
            .O(N__22244),
            .I(N__22240));
    InMux I__4469 (
            .O(N__22243),
            .I(N__22237));
    LocalMux I__4468 (
            .O(N__22240),
            .I(N__22234));
    LocalMux I__4467 (
            .O(N__22237),
            .I(N__22231));
    Span4Mux_v I__4466 (
            .O(N__22234),
            .I(N__22228));
    Odrv4 I__4465 (
            .O(N__22231),
            .I(\eeprom.n2606 ));
    Odrv4 I__4464 (
            .O(N__22228),
            .I(\eeprom.n2606 ));
    CascadeMux I__4463 (
            .O(N__22223),
            .I(\eeprom.n2606_cascade_ ));
    InMux I__4462 (
            .O(N__22220),
            .I(N__22217));
    LocalMux I__4461 (
            .O(N__22217),
            .I(\eeprom.n10_adj_332 ));
    InMux I__4460 (
            .O(N__22214),
            .I(N__22210));
    InMux I__4459 (
            .O(N__22213),
            .I(N__22206));
    LocalMux I__4458 (
            .O(N__22210),
            .I(N__22203));
    InMux I__4457 (
            .O(N__22209),
            .I(N__22200));
    LocalMux I__4456 (
            .O(N__22206),
            .I(N__22195));
    Span4Mux_v I__4455 (
            .O(N__22203),
            .I(N__22195));
    LocalMux I__4454 (
            .O(N__22200),
            .I(\eeprom.n2718 ));
    Odrv4 I__4453 (
            .O(N__22195),
            .I(\eeprom.n2718 ));
    CascadeMux I__4452 (
            .O(N__22190),
            .I(N__22187));
    InMux I__4451 (
            .O(N__22187),
            .I(N__22184));
    LocalMux I__4450 (
            .O(N__22184),
            .I(\eeprom.n5213 ));
    InMux I__4449 (
            .O(N__22181),
            .I(N__22178));
    LocalMux I__4448 (
            .O(N__22178),
            .I(\eeprom.n5215 ));
    InMux I__4447 (
            .O(N__22175),
            .I(N__22172));
    LocalMux I__4446 (
            .O(N__22172),
            .I(\eeprom.n4830 ));
    InMux I__4445 (
            .O(N__22169),
            .I(N__22166));
    LocalMux I__4444 (
            .O(N__22166),
            .I(N__22163));
    Span4Mux_v I__4443 (
            .O(N__22163),
            .I(N__22160));
    Odrv4 I__4442 (
            .O(N__22160),
            .I(\eeprom.n2682 ));
    InMux I__4441 (
            .O(N__22157),
            .I(N__22152));
    InMux I__4440 (
            .O(N__22156),
            .I(N__22149));
    InMux I__4439 (
            .O(N__22155),
            .I(N__22146));
    LocalMux I__4438 (
            .O(N__22152),
            .I(\eeprom.n2714 ));
    LocalMux I__4437 (
            .O(N__22149),
            .I(\eeprom.n2714 ));
    LocalMux I__4436 (
            .O(N__22146),
            .I(\eeprom.n2714 ));
    InMux I__4435 (
            .O(N__22139),
            .I(N__22135));
    InMux I__4434 (
            .O(N__22138),
            .I(N__22131));
    LocalMux I__4433 (
            .O(N__22135),
            .I(N__22128));
    InMux I__4432 (
            .O(N__22134),
            .I(N__22125));
    LocalMux I__4431 (
            .O(N__22131),
            .I(\eeprom.n2609 ));
    Odrv4 I__4430 (
            .O(N__22128),
            .I(\eeprom.n2609 ));
    LocalMux I__4429 (
            .O(N__22125),
            .I(\eeprom.n2609 ));
    InMux I__4428 (
            .O(N__22118),
            .I(N__22115));
    LocalMux I__4427 (
            .O(N__22115),
            .I(\eeprom.n2482 ));
    CascadeMux I__4426 (
            .O(N__22112),
            .I(N__22109));
    InMux I__4425 (
            .O(N__22109),
            .I(N__22105));
    CascadeMux I__4424 (
            .O(N__22108),
            .I(N__22102));
    LocalMux I__4423 (
            .O(N__22105),
            .I(N__22099));
    InMux I__4422 (
            .O(N__22102),
            .I(N__22096));
    Span4Mux_h I__4421 (
            .O(N__22099),
            .I(N__22092));
    LocalMux I__4420 (
            .O(N__22096),
            .I(N__22089));
    InMux I__4419 (
            .O(N__22095),
            .I(N__22086));
    Odrv4 I__4418 (
            .O(N__22092),
            .I(\eeprom.n2415 ));
    Odrv4 I__4417 (
            .O(N__22089),
            .I(\eeprom.n2415 ));
    LocalMux I__4416 (
            .O(N__22086),
            .I(\eeprom.n2415 ));
    CascadeMux I__4415 (
            .O(N__22079),
            .I(\eeprom.n13_adj_329_cascade_ ));
    CascadeMux I__4414 (
            .O(N__22076),
            .I(\eeprom.n2539_cascade_ ));
    CascadeMux I__4413 (
            .O(N__22073),
            .I(N__22070));
    InMux I__4412 (
            .O(N__22070),
            .I(N__22067));
    LocalMux I__4411 (
            .O(N__22067),
            .I(N__22064));
    Span4Mux_h I__4410 (
            .O(N__22064),
            .I(N__22061));
    Odrv4 I__4409 (
            .O(N__22061),
            .I(\eeprom.n2683 ));
    InMux I__4408 (
            .O(N__22058),
            .I(N__22055));
    LocalMux I__4407 (
            .O(N__22055),
            .I(N__22052));
    Span4Mux_h I__4406 (
            .O(N__22052),
            .I(N__22049));
    Odrv4 I__4405 (
            .O(N__22049),
            .I(\eeprom.n2681 ));
    InMux I__4404 (
            .O(N__22046),
            .I(N__22043));
    LocalMux I__4403 (
            .O(N__22043),
            .I(N__22039));
    InMux I__4402 (
            .O(N__22042),
            .I(N__22036));
    Span4Mux_h I__4401 (
            .O(N__22039),
            .I(N__22031));
    LocalMux I__4400 (
            .O(N__22036),
            .I(N__22031));
    Odrv4 I__4399 (
            .O(N__22031),
            .I(\eeprom.n2713 ));
    CascadeMux I__4398 (
            .O(N__22028),
            .I(\eeprom.n2713_cascade_ ));
    InMux I__4397 (
            .O(N__22025),
            .I(N__22021));
    InMux I__4396 (
            .O(N__22024),
            .I(N__22018));
    LocalMux I__4395 (
            .O(N__22021),
            .I(N__22015));
    LocalMux I__4394 (
            .O(N__22018),
            .I(N__22012));
    Span4Mux_h I__4393 (
            .O(N__22015),
            .I(N__22006));
    Span4Mux_h I__4392 (
            .O(N__22012),
            .I(N__22006));
    InMux I__4391 (
            .O(N__22011),
            .I(N__22003));
    Odrv4 I__4390 (
            .O(N__22006),
            .I(\eeprom.n2715 ));
    LocalMux I__4389 (
            .O(N__22003),
            .I(\eeprom.n2715 ));
    CascadeMux I__4388 (
            .O(N__21998),
            .I(N__21994));
    CascadeMux I__4387 (
            .O(N__21997),
            .I(N__21990));
    InMux I__4386 (
            .O(N__21994),
            .I(N__21987));
    InMux I__4385 (
            .O(N__21993),
            .I(N__21982));
    InMux I__4384 (
            .O(N__21990),
            .I(N__21982));
    LocalMux I__4383 (
            .O(N__21987),
            .I(N__21979));
    LocalMux I__4382 (
            .O(N__21982),
            .I(\eeprom.n2219 ));
    Odrv4 I__4381 (
            .O(N__21979),
            .I(\eeprom.n2219 ));
    CascadeMux I__4380 (
            .O(N__21974),
            .I(N__21971));
    InMux I__4379 (
            .O(N__21971),
            .I(N__21968));
    LocalMux I__4378 (
            .O(N__21968),
            .I(N__21965));
    Span4Mux_v I__4377 (
            .O(N__21965),
            .I(N__21962));
    Odrv4 I__4376 (
            .O(N__21962),
            .I(\eeprom.n3723 ));
    CascadeMux I__4375 (
            .O(N__21959),
            .I(N__21956));
    InMux I__4374 (
            .O(N__21956),
            .I(N__21951));
    InMux I__4373 (
            .O(N__21955),
            .I(N__21948));
    InMux I__4372 (
            .O(N__21954),
            .I(N__21945));
    LocalMux I__4371 (
            .O(N__21951),
            .I(\eeprom.n2210 ));
    LocalMux I__4370 (
            .O(N__21948),
            .I(\eeprom.n2210 ));
    LocalMux I__4369 (
            .O(N__21945),
            .I(\eeprom.n2210 ));
    InMux I__4368 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__4367 (
            .O(N__21935),
            .I(\eeprom.n6_adj_321 ));
    InMux I__4366 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__4365 (
            .O(N__21929),
            .I(\eeprom.n2483 ));
    InMux I__4364 (
            .O(N__21926),
            .I(N__21922));
    CascadeMux I__4363 (
            .O(N__21925),
            .I(N__21918));
    LocalMux I__4362 (
            .O(N__21922),
            .I(N__21915));
    CascadeMux I__4361 (
            .O(N__21921),
            .I(N__21912));
    InMux I__4360 (
            .O(N__21918),
            .I(N__21909));
    Span4Mux_h I__4359 (
            .O(N__21915),
            .I(N__21906));
    InMux I__4358 (
            .O(N__21912),
            .I(N__21903));
    LocalMux I__4357 (
            .O(N__21909),
            .I(N__21900));
    Odrv4 I__4356 (
            .O(N__21906),
            .I(\eeprom.n2416 ));
    LocalMux I__4355 (
            .O(N__21903),
            .I(\eeprom.n2416 ));
    Odrv4 I__4354 (
            .O(N__21900),
            .I(\eeprom.n2416 ));
    InMux I__4353 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__4352 (
            .O(N__21890),
            .I(\eeprom.n2485 ));
    CascadeMux I__4351 (
            .O(N__21887),
            .I(N__21884));
    InMux I__4350 (
            .O(N__21884),
            .I(N__21881));
    LocalMux I__4349 (
            .O(N__21881),
            .I(N__21877));
    InMux I__4348 (
            .O(N__21880),
            .I(N__21873));
    Span4Mux_h I__4347 (
            .O(N__21877),
            .I(N__21870));
    InMux I__4346 (
            .O(N__21876),
            .I(N__21867));
    LocalMux I__4345 (
            .O(N__21873),
            .I(N__21864));
    Odrv4 I__4344 (
            .O(N__21870),
            .I(\eeprom.n2418 ));
    LocalMux I__4343 (
            .O(N__21867),
            .I(\eeprom.n2418 ));
    Odrv4 I__4342 (
            .O(N__21864),
            .I(\eeprom.n2418 ));
    InMux I__4341 (
            .O(N__21857),
            .I(N__21854));
    LocalMux I__4340 (
            .O(N__21854),
            .I(N__21851));
    Odrv4 I__4339 (
            .O(N__21851),
            .I(\eeprom.n2477 ));
    CascadeMux I__4338 (
            .O(N__21848),
            .I(N__21845));
    InMux I__4337 (
            .O(N__21845),
            .I(N__21841));
    InMux I__4336 (
            .O(N__21844),
            .I(N__21838));
    LocalMux I__4335 (
            .O(N__21841),
            .I(N__21834));
    LocalMux I__4334 (
            .O(N__21838),
            .I(N__21831));
    InMux I__4333 (
            .O(N__21837),
            .I(N__21828));
    Odrv4 I__4332 (
            .O(N__21834),
            .I(\eeprom.n2410 ));
    Odrv4 I__4331 (
            .O(N__21831),
            .I(\eeprom.n2410 ));
    LocalMux I__4330 (
            .O(N__21828),
            .I(\eeprom.n2410 ));
    InMux I__4329 (
            .O(N__21821),
            .I(N__21817));
    InMux I__4328 (
            .O(N__21820),
            .I(N__21814));
    LocalMux I__4327 (
            .O(N__21817),
            .I(N__21810));
    LocalMux I__4326 (
            .O(N__21814),
            .I(N__21807));
    InMux I__4325 (
            .O(N__21813),
            .I(N__21804));
    Odrv4 I__4324 (
            .O(N__21810),
            .I(\eeprom.n2408 ));
    Odrv4 I__4323 (
            .O(N__21807),
            .I(\eeprom.n2408 ));
    LocalMux I__4322 (
            .O(N__21804),
            .I(\eeprom.n2408 ));
    InMux I__4321 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__4320 (
            .O(N__21794),
            .I(N__21791));
    Odrv4 I__4319 (
            .O(N__21791),
            .I(\eeprom.n2475 ));
    InMux I__4318 (
            .O(N__21788),
            .I(N__21785));
    LocalMux I__4317 (
            .O(N__21785),
            .I(N__21782));
    Odrv4 I__4316 (
            .O(N__21782),
            .I(\eeprom.n2486 ));
    InMux I__4315 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__4314 (
            .O(N__21776),
            .I(\eeprom.n2484 ));
    InMux I__4313 (
            .O(N__21773),
            .I(N__21769));
    CascadeMux I__4312 (
            .O(N__21772),
            .I(N__21766));
    LocalMux I__4311 (
            .O(N__21769),
            .I(N__21762));
    InMux I__4310 (
            .O(N__21766),
            .I(N__21759));
    CascadeMux I__4309 (
            .O(N__21765),
            .I(N__21756));
    Span4Mux_h I__4308 (
            .O(N__21762),
            .I(N__21753));
    LocalMux I__4307 (
            .O(N__21759),
            .I(N__21750));
    InMux I__4306 (
            .O(N__21756),
            .I(N__21747));
    Odrv4 I__4305 (
            .O(N__21753),
            .I(\eeprom.n2417 ));
    Odrv4 I__4304 (
            .O(N__21750),
            .I(\eeprom.n2417 ));
    LocalMux I__4303 (
            .O(N__21747),
            .I(\eeprom.n2417 ));
    CascadeMux I__4302 (
            .O(N__21740),
            .I(N__21731));
    CascadeMux I__4301 (
            .O(N__21739),
            .I(N__21728));
    CascadeMux I__4300 (
            .O(N__21738),
            .I(N__21724));
    InMux I__4299 (
            .O(N__21737),
            .I(N__21718));
    InMux I__4298 (
            .O(N__21736),
            .I(N__21713));
    InMux I__4297 (
            .O(N__21735),
            .I(N__21713));
    InMux I__4296 (
            .O(N__21734),
            .I(N__21710));
    InMux I__4295 (
            .O(N__21731),
            .I(N__21703));
    InMux I__4294 (
            .O(N__21728),
            .I(N__21703));
    InMux I__4293 (
            .O(N__21727),
            .I(N__21703));
    InMux I__4292 (
            .O(N__21724),
            .I(N__21696));
    InMux I__4291 (
            .O(N__21723),
            .I(N__21696));
    InMux I__4290 (
            .O(N__21722),
            .I(N__21696));
    InMux I__4289 (
            .O(N__21721),
            .I(N__21693));
    LocalMux I__4288 (
            .O(N__21718),
            .I(\eeprom.n2242 ));
    LocalMux I__4287 (
            .O(N__21713),
            .I(\eeprom.n2242 ));
    LocalMux I__4286 (
            .O(N__21710),
            .I(\eeprom.n2242 ));
    LocalMux I__4285 (
            .O(N__21703),
            .I(\eeprom.n2242 ));
    LocalMux I__4284 (
            .O(N__21696),
            .I(\eeprom.n2242 ));
    LocalMux I__4283 (
            .O(N__21693),
            .I(\eeprom.n2242 ));
    InMux I__4282 (
            .O(N__21680),
            .I(N__21677));
    LocalMux I__4281 (
            .O(N__21677),
            .I(\eeprom.n5501 ));
    InMux I__4280 (
            .O(N__21674),
            .I(N__21671));
    LocalMux I__4279 (
            .O(N__21671),
            .I(\eeprom.n2081 ));
    InMux I__4278 (
            .O(N__21668),
            .I(N__21665));
    LocalMux I__4277 (
            .O(N__21665),
            .I(N__21662));
    Odrv4 I__4276 (
            .O(N__21662),
            .I(\eeprom.n2086 ));
    InMux I__4275 (
            .O(N__21659),
            .I(N__21656));
    LocalMux I__4274 (
            .O(N__21656),
            .I(N__21653));
    Odrv4 I__4273 (
            .O(N__21653),
            .I(\eeprom.n5061 ));
    CascadeMux I__4272 (
            .O(N__21650),
            .I(\eeprom.n2118_cascade_ ));
    InMux I__4271 (
            .O(N__21647),
            .I(N__21644));
    LocalMux I__4270 (
            .O(N__21644),
            .I(\eeprom.n4788 ));
    CascadeMux I__4269 (
            .O(N__21641),
            .I(N__21637));
    InMux I__4268 (
            .O(N__21640),
            .I(N__21633));
    InMux I__4267 (
            .O(N__21637),
            .I(N__21630));
    InMux I__4266 (
            .O(N__21636),
            .I(N__21627));
    LocalMux I__4265 (
            .O(N__21633),
            .I(N__21624));
    LocalMux I__4264 (
            .O(N__21630),
            .I(\eeprom.n2212 ));
    LocalMux I__4263 (
            .O(N__21627),
            .I(\eeprom.n2212 ));
    Odrv4 I__4262 (
            .O(N__21624),
            .I(\eeprom.n2212 ));
    InMux I__4261 (
            .O(N__21617),
            .I(N__21612));
    InMux I__4260 (
            .O(N__21616),
            .I(N__21609));
    InMux I__4259 (
            .O(N__21615),
            .I(N__21606));
    LocalMux I__4258 (
            .O(N__21612),
            .I(N__21603));
    LocalMux I__4257 (
            .O(N__21609),
            .I(N__21600));
    LocalMux I__4256 (
            .O(N__21606),
            .I(\eeprom.n2019 ));
    Odrv4 I__4255 (
            .O(N__21603),
            .I(\eeprom.n2019 ));
    Odrv4 I__4254 (
            .O(N__21600),
            .I(\eeprom.n2019 ));
    CascadeMux I__4253 (
            .O(N__21593),
            .I(N__21590));
    InMux I__4252 (
            .O(N__21590),
            .I(N__21587));
    LocalMux I__4251 (
            .O(N__21587),
            .I(N__21584));
    Span4Mux_h I__4250 (
            .O(N__21584),
            .I(N__21581));
    Odrv4 I__4249 (
            .O(N__21581),
            .I(\eeprom.n3721 ));
    InMux I__4248 (
            .O(N__21578),
            .I(N__21573));
    InMux I__4247 (
            .O(N__21577),
            .I(N__21570));
    InMux I__4246 (
            .O(N__21576),
            .I(N__21567));
    LocalMux I__4245 (
            .O(N__21573),
            .I(N__21560));
    LocalMux I__4244 (
            .O(N__21570),
            .I(N__21560));
    LocalMux I__4243 (
            .O(N__21567),
            .I(N__21560));
    Span4Mux_v I__4242 (
            .O(N__21560),
            .I(N__21557));
    Span4Mux_h I__4241 (
            .O(N__21557),
            .I(N__21554));
    Odrv4 I__4240 (
            .O(N__21554),
            .I(\eeprom.n3619 ));
    InMux I__4239 (
            .O(N__21551),
            .I(N__21548));
    LocalMux I__4238 (
            .O(N__21548),
            .I(\eeprom.n2085 ));
    InMux I__4237 (
            .O(N__21545),
            .I(\eeprom.n3980 ));
    InMux I__4236 (
            .O(N__21542),
            .I(N__21538));
    InMux I__4235 (
            .O(N__21541),
            .I(N__21535));
    LocalMux I__4234 (
            .O(N__21538),
            .I(\eeprom.n2084 ));
    LocalMux I__4233 (
            .O(N__21535),
            .I(\eeprom.n2084 ));
    InMux I__4232 (
            .O(N__21530),
            .I(\eeprom.n3981 ));
    InMux I__4231 (
            .O(N__21527),
            .I(\eeprom.n3982 ));
    InMux I__4230 (
            .O(N__21524),
            .I(N__21521));
    LocalMux I__4229 (
            .O(N__21521),
            .I(\eeprom.n2082 ));
    InMux I__4228 (
            .O(N__21518),
            .I(\eeprom.n3983 ));
    InMux I__4227 (
            .O(N__21515),
            .I(\eeprom.n3984 ));
    InMux I__4226 (
            .O(N__21512),
            .I(N__21509));
    LocalMux I__4225 (
            .O(N__21509),
            .I(\eeprom.n2080 ));
    InMux I__4224 (
            .O(N__21506),
            .I(\eeprom.n3985 ));
    InMux I__4223 (
            .O(N__21503),
            .I(\eeprom.n3986 ));
    InMux I__4222 (
            .O(N__21500),
            .I(bfn_23_19_0_));
    InMux I__4221 (
            .O(N__21497),
            .I(N__21493));
    InMux I__4220 (
            .O(N__21496),
            .I(N__21490));
    LocalMux I__4219 (
            .O(N__21493),
            .I(N__21484));
    LocalMux I__4218 (
            .O(N__21490),
            .I(N__21484));
    InMux I__4217 (
            .O(N__21489),
            .I(N__21481));
    Odrv4 I__4216 (
            .O(N__21484),
            .I(\eeprom.n2704 ));
    LocalMux I__4215 (
            .O(N__21481),
            .I(\eeprom.n2704 ));
    CascadeMux I__4214 (
            .O(N__21476),
            .I(N__21466));
    CascadeMux I__4213 (
            .O(N__21475),
            .I(N__21463));
    CascadeMux I__4212 (
            .O(N__21474),
            .I(N__21460));
    CascadeMux I__4211 (
            .O(N__21473),
            .I(N__21457));
    CascadeMux I__4210 (
            .O(N__21472),
            .I(N__21454));
    CascadeMux I__4209 (
            .O(N__21471),
            .I(N__21451));
    CascadeMux I__4208 (
            .O(N__21470),
            .I(N__21448));
    CascadeMux I__4207 (
            .O(N__21469),
            .I(N__21445));
    InMux I__4206 (
            .O(N__21466),
            .I(N__21434));
    InMux I__4205 (
            .O(N__21463),
            .I(N__21434));
    InMux I__4204 (
            .O(N__21460),
            .I(N__21434));
    InMux I__4203 (
            .O(N__21457),
            .I(N__21434));
    InMux I__4202 (
            .O(N__21454),
            .I(N__21425));
    InMux I__4201 (
            .O(N__21451),
            .I(N__21425));
    InMux I__4200 (
            .O(N__21448),
            .I(N__21425));
    InMux I__4199 (
            .O(N__21445),
            .I(N__21425));
    CascadeMux I__4198 (
            .O(N__21444),
            .I(N__21422));
    CascadeMux I__4197 (
            .O(N__21443),
            .I(N__21419));
    LocalMux I__4196 (
            .O(N__21434),
            .I(N__21414));
    LocalMux I__4195 (
            .O(N__21425),
            .I(N__21414));
    InMux I__4194 (
            .O(N__21422),
            .I(N__21409));
    InMux I__4193 (
            .O(N__21419),
            .I(N__21409));
    Odrv4 I__4192 (
            .O(N__21414),
            .I(\eeprom.n2737 ));
    LocalMux I__4191 (
            .O(N__21409),
            .I(\eeprom.n2737 ));
    InMux I__4190 (
            .O(N__21404),
            .I(\eeprom.n4071 ));
    InMux I__4189 (
            .O(N__21401),
            .I(N__21397));
    InMux I__4188 (
            .O(N__21400),
            .I(N__21394));
    LocalMux I__4187 (
            .O(N__21397),
            .I(N__21391));
    LocalMux I__4186 (
            .O(N__21394),
            .I(N__21388));
    Span4Mux_h I__4185 (
            .O(N__21391),
            .I(N__21385));
    Odrv4 I__4184 (
            .O(N__21388),
            .I(\eeprom.n2803 ));
    Odrv4 I__4183 (
            .O(N__21385),
            .I(\eeprom.n2803 ));
    CascadeMux I__4182 (
            .O(N__21380),
            .I(\eeprom.n5005_cascade_ ));
    CascadeMux I__4181 (
            .O(N__21377),
            .I(\eeprom.n5009_cascade_ ));
    CascadeMux I__4180 (
            .O(N__21374),
            .I(\eeprom.n2044_cascade_ ));
    CascadeMux I__4179 (
            .O(N__21371),
            .I(\eeprom.n2116_cascade_ ));
    InMux I__4178 (
            .O(N__21368),
            .I(bfn_23_18_0_));
    InMux I__4177 (
            .O(N__21365),
            .I(N__21361));
    InMux I__4176 (
            .O(N__21364),
            .I(N__21357));
    LocalMux I__4175 (
            .O(N__21361),
            .I(N__21354));
    InMux I__4174 (
            .O(N__21360),
            .I(N__21351));
    LocalMux I__4173 (
            .O(N__21357),
            .I(N__21348));
    Span4Mux_h I__4172 (
            .O(N__21354),
            .I(N__21345));
    LocalMux I__4171 (
            .O(N__21351),
            .I(N__21340));
    Span4Mux_h I__4170 (
            .O(N__21348),
            .I(N__21340));
    Odrv4 I__4169 (
            .O(N__21345),
            .I(\eeprom.n2811 ));
    Odrv4 I__4168 (
            .O(N__21340),
            .I(\eeprom.n2811 ));
    InMux I__4167 (
            .O(N__21335),
            .I(\eeprom.n4063 ));
    InMux I__4166 (
            .O(N__21332),
            .I(N__21328));
    InMux I__4165 (
            .O(N__21331),
            .I(N__21325));
    LocalMux I__4164 (
            .O(N__21328),
            .I(N__21319));
    LocalMux I__4163 (
            .O(N__21325),
            .I(N__21319));
    InMux I__4162 (
            .O(N__21324),
            .I(N__21316));
    Odrv4 I__4161 (
            .O(N__21319),
            .I(\eeprom.n2711 ));
    LocalMux I__4160 (
            .O(N__21316),
            .I(\eeprom.n2711 ));
    InMux I__4159 (
            .O(N__21311),
            .I(N__21305));
    InMux I__4158 (
            .O(N__21310),
            .I(N__21305));
    LocalMux I__4157 (
            .O(N__21305),
            .I(N__21301));
    InMux I__4156 (
            .O(N__21304),
            .I(N__21298));
    Span4Mux_h I__4155 (
            .O(N__21301),
            .I(N__21293));
    LocalMux I__4154 (
            .O(N__21298),
            .I(N__21293));
    Odrv4 I__4153 (
            .O(N__21293),
            .I(\eeprom.n2810 ));
    InMux I__4152 (
            .O(N__21290),
            .I(bfn_22_26_0_));
    InMux I__4151 (
            .O(N__21287),
            .I(N__21283));
    InMux I__4150 (
            .O(N__21286),
            .I(N__21280));
    LocalMux I__4149 (
            .O(N__21283),
            .I(\eeprom.n2710 ));
    LocalMux I__4148 (
            .O(N__21280),
            .I(\eeprom.n2710 ));
    InMux I__4147 (
            .O(N__21275),
            .I(N__21270));
    CascadeMux I__4146 (
            .O(N__21274),
            .I(N__21267));
    InMux I__4145 (
            .O(N__21273),
            .I(N__21264));
    LocalMux I__4144 (
            .O(N__21270),
            .I(N__21261));
    InMux I__4143 (
            .O(N__21267),
            .I(N__21258));
    LocalMux I__4142 (
            .O(N__21264),
            .I(N__21255));
    Span4Mux_h I__4141 (
            .O(N__21261),
            .I(N__21252));
    LocalMux I__4140 (
            .O(N__21258),
            .I(N__21249));
    Span4Mux_h I__4139 (
            .O(N__21255),
            .I(N__21246));
    Odrv4 I__4138 (
            .O(N__21252),
            .I(\eeprom.n2809 ));
    Odrv4 I__4137 (
            .O(N__21249),
            .I(\eeprom.n2809 ));
    Odrv4 I__4136 (
            .O(N__21246),
            .I(\eeprom.n2809 ));
    InMux I__4135 (
            .O(N__21239),
            .I(\eeprom.n4065 ));
    InMux I__4134 (
            .O(N__21236),
            .I(N__21232));
    InMux I__4133 (
            .O(N__21235),
            .I(N__21229));
    LocalMux I__4132 (
            .O(N__21232),
            .I(N__21224));
    LocalMux I__4131 (
            .O(N__21229),
            .I(N__21224));
    Span4Mux_h I__4130 (
            .O(N__21224),
            .I(N__21220));
    InMux I__4129 (
            .O(N__21223),
            .I(N__21217));
    Odrv4 I__4128 (
            .O(N__21220),
            .I(\eeprom.n2709 ));
    LocalMux I__4127 (
            .O(N__21217),
            .I(\eeprom.n2709 ));
    InMux I__4126 (
            .O(N__21212),
            .I(N__21207));
    InMux I__4125 (
            .O(N__21211),
            .I(N__21204));
    InMux I__4124 (
            .O(N__21210),
            .I(N__21201));
    LocalMux I__4123 (
            .O(N__21207),
            .I(N__21194));
    LocalMux I__4122 (
            .O(N__21204),
            .I(N__21194));
    LocalMux I__4121 (
            .O(N__21201),
            .I(N__21194));
    Span4Mux_v I__4120 (
            .O(N__21194),
            .I(N__21191));
    Odrv4 I__4119 (
            .O(N__21191),
            .I(\eeprom.n2808 ));
    InMux I__4118 (
            .O(N__21188),
            .I(\eeprom.n4066 ));
    InMux I__4117 (
            .O(N__21185),
            .I(N__21181));
    InMux I__4116 (
            .O(N__21184),
            .I(N__21178));
    LocalMux I__4115 (
            .O(N__21181),
            .I(N__21172));
    LocalMux I__4114 (
            .O(N__21178),
            .I(N__21172));
    InMux I__4113 (
            .O(N__21177),
            .I(N__21169));
    Odrv12 I__4112 (
            .O(N__21172),
            .I(\eeprom.n2708 ));
    LocalMux I__4111 (
            .O(N__21169),
            .I(\eeprom.n2708 ));
    CascadeMux I__4110 (
            .O(N__21164),
            .I(N__21160));
    InMux I__4109 (
            .O(N__21163),
            .I(N__21156));
    InMux I__4108 (
            .O(N__21160),
            .I(N__21153));
    InMux I__4107 (
            .O(N__21159),
            .I(N__21150));
    LocalMux I__4106 (
            .O(N__21156),
            .I(N__21143));
    LocalMux I__4105 (
            .O(N__21153),
            .I(N__21143));
    LocalMux I__4104 (
            .O(N__21150),
            .I(N__21143));
    Span4Mux_v I__4103 (
            .O(N__21143),
            .I(N__21140));
    Odrv4 I__4102 (
            .O(N__21140),
            .I(\eeprom.n2807 ));
    InMux I__4101 (
            .O(N__21137),
            .I(\eeprom.n4067 ));
    InMux I__4100 (
            .O(N__21134),
            .I(N__21130));
    InMux I__4099 (
            .O(N__21133),
            .I(N__21127));
    LocalMux I__4098 (
            .O(N__21130),
            .I(N__21123));
    LocalMux I__4097 (
            .O(N__21127),
            .I(N__21120));
    InMux I__4096 (
            .O(N__21126),
            .I(N__21117));
    Odrv4 I__4095 (
            .O(N__21123),
            .I(\eeprom.n2707 ));
    Odrv4 I__4094 (
            .O(N__21120),
            .I(\eeprom.n2707 ));
    LocalMux I__4093 (
            .O(N__21117),
            .I(\eeprom.n2707 ));
    CascadeMux I__4092 (
            .O(N__21110),
            .I(N__21106));
    CascadeMux I__4091 (
            .O(N__21109),
            .I(N__21103));
    InMux I__4090 (
            .O(N__21106),
            .I(N__21099));
    InMux I__4089 (
            .O(N__21103),
            .I(N__21096));
    InMux I__4088 (
            .O(N__21102),
            .I(N__21093));
    LocalMux I__4087 (
            .O(N__21099),
            .I(N__21088));
    LocalMux I__4086 (
            .O(N__21096),
            .I(N__21088));
    LocalMux I__4085 (
            .O(N__21093),
            .I(N__21085));
    Span4Mux_h I__4084 (
            .O(N__21088),
            .I(N__21082));
    Odrv4 I__4083 (
            .O(N__21085),
            .I(\eeprom.n2806 ));
    Odrv4 I__4082 (
            .O(N__21082),
            .I(\eeprom.n2806 ));
    InMux I__4081 (
            .O(N__21077),
            .I(\eeprom.n4068 ));
    InMux I__4080 (
            .O(N__21074),
            .I(N__21069));
    InMux I__4079 (
            .O(N__21073),
            .I(N__21066));
    InMux I__4078 (
            .O(N__21072),
            .I(N__21063));
    LocalMux I__4077 (
            .O(N__21069),
            .I(N__21060));
    LocalMux I__4076 (
            .O(N__21066),
            .I(N__21057));
    LocalMux I__4075 (
            .O(N__21063),
            .I(N__21052));
    Span4Mux_h I__4074 (
            .O(N__21060),
            .I(N__21052));
    Odrv4 I__4073 (
            .O(N__21057),
            .I(\eeprom.n2805 ));
    Odrv4 I__4072 (
            .O(N__21052),
            .I(\eeprom.n2805 ));
    InMux I__4071 (
            .O(N__21047),
            .I(\eeprom.n4069 ));
    InMux I__4070 (
            .O(N__21044),
            .I(N__21040));
    InMux I__4069 (
            .O(N__21043),
            .I(N__21037));
    LocalMux I__4068 (
            .O(N__21040),
            .I(N__21032));
    LocalMux I__4067 (
            .O(N__21037),
            .I(N__21032));
    Odrv4 I__4066 (
            .O(N__21032),
            .I(\eeprom.n2705 ));
    CascadeMux I__4065 (
            .O(N__21029),
            .I(N__21025));
    CascadeMux I__4064 (
            .O(N__21028),
            .I(N__21021));
    InMux I__4063 (
            .O(N__21025),
            .I(N__21018));
    InMux I__4062 (
            .O(N__21024),
            .I(N__21015));
    InMux I__4061 (
            .O(N__21021),
            .I(N__21012));
    LocalMux I__4060 (
            .O(N__21018),
            .I(N__21007));
    LocalMux I__4059 (
            .O(N__21015),
            .I(N__21007));
    LocalMux I__4058 (
            .O(N__21012),
            .I(N__21004));
    Span4Mux_h I__4057 (
            .O(N__21007),
            .I(N__21001));
    Odrv4 I__4056 (
            .O(N__21004),
            .I(\eeprom.n2804 ));
    Odrv4 I__4055 (
            .O(N__21001),
            .I(\eeprom.n2804 ));
    InMux I__4054 (
            .O(N__20996),
            .I(\eeprom.n4070 ));
    CascadeMux I__4053 (
            .O(N__20993),
            .I(\eeprom.n2737_cascade_ ));
    InMux I__4052 (
            .O(N__20990),
            .I(N__20987));
    LocalMux I__4051 (
            .O(N__20987),
            .I(N__20983));
    InMux I__4050 (
            .O(N__20986),
            .I(N__20979));
    Span4Mux_v I__4049 (
            .O(N__20983),
            .I(N__20976));
    InMux I__4048 (
            .O(N__20982),
            .I(N__20973));
    LocalMux I__4047 (
            .O(N__20979),
            .I(N__20970));
    Odrv4 I__4046 (
            .O(N__20976),
            .I(\eeprom.n2818 ));
    LocalMux I__4045 (
            .O(N__20973),
            .I(\eeprom.n2818 ));
    Odrv4 I__4044 (
            .O(N__20970),
            .I(\eeprom.n2818 ));
    InMux I__4043 (
            .O(N__20963),
            .I(bfn_22_25_0_));
    InMux I__4042 (
            .O(N__20960),
            .I(N__20955));
    CascadeMux I__4041 (
            .O(N__20959),
            .I(N__20952));
    CascadeMux I__4040 (
            .O(N__20958),
            .I(N__20949));
    LocalMux I__4039 (
            .O(N__20955),
            .I(N__20946));
    InMux I__4038 (
            .O(N__20952),
            .I(N__20943));
    InMux I__4037 (
            .O(N__20949),
            .I(N__20940));
    Span4Mux_h I__4036 (
            .O(N__20946),
            .I(N__20935));
    LocalMux I__4035 (
            .O(N__20943),
            .I(N__20935));
    LocalMux I__4034 (
            .O(N__20940),
            .I(\eeprom.n2817 ));
    Odrv4 I__4033 (
            .O(N__20935),
            .I(\eeprom.n2817 ));
    InMux I__4032 (
            .O(N__20930),
            .I(\eeprom.n4057 ));
    InMux I__4031 (
            .O(N__20927),
            .I(N__20923));
    InMux I__4030 (
            .O(N__20926),
            .I(N__20920));
    LocalMux I__4029 (
            .O(N__20923),
            .I(N__20917));
    LocalMux I__4028 (
            .O(N__20920),
            .I(N__20913));
    Span4Mux_v I__4027 (
            .O(N__20917),
            .I(N__20910));
    InMux I__4026 (
            .O(N__20916),
            .I(N__20907));
    Odrv4 I__4025 (
            .O(N__20913),
            .I(\eeprom.n2717 ));
    Odrv4 I__4024 (
            .O(N__20910),
            .I(\eeprom.n2717 ));
    LocalMux I__4023 (
            .O(N__20907),
            .I(\eeprom.n2717 ));
    InMux I__4022 (
            .O(N__20900),
            .I(N__20897));
    LocalMux I__4021 (
            .O(N__20897),
            .I(N__20893));
    InMux I__4020 (
            .O(N__20896),
            .I(N__20890));
    Span4Mux_h I__4019 (
            .O(N__20893),
            .I(N__20884));
    LocalMux I__4018 (
            .O(N__20890),
            .I(N__20884));
    InMux I__4017 (
            .O(N__20889),
            .I(N__20881));
    Odrv4 I__4016 (
            .O(N__20884),
            .I(\eeprom.n2816 ));
    LocalMux I__4015 (
            .O(N__20881),
            .I(\eeprom.n2816 ));
    InMux I__4014 (
            .O(N__20876),
            .I(\eeprom.n4058 ));
    InMux I__4013 (
            .O(N__20873),
            .I(N__20869));
    InMux I__4012 (
            .O(N__20872),
            .I(N__20866));
    LocalMux I__4011 (
            .O(N__20869),
            .I(N__20861));
    LocalMux I__4010 (
            .O(N__20866),
            .I(N__20861));
    Odrv4 I__4009 (
            .O(N__20861),
            .I(\eeprom.n2716 ));
    InMux I__4008 (
            .O(N__20858),
            .I(N__20855));
    LocalMux I__4007 (
            .O(N__20855),
            .I(N__20851));
    CascadeMux I__4006 (
            .O(N__20854),
            .I(N__20848));
    Span4Mux_h I__4005 (
            .O(N__20851),
            .I(N__20844));
    InMux I__4004 (
            .O(N__20848),
            .I(N__20841));
    CascadeMux I__4003 (
            .O(N__20847),
            .I(N__20838));
    Sp12to4 I__4002 (
            .O(N__20844),
            .I(N__20835));
    LocalMux I__4001 (
            .O(N__20841),
            .I(N__20832));
    InMux I__4000 (
            .O(N__20838),
            .I(N__20829));
    Odrv12 I__3999 (
            .O(N__20835),
            .I(\eeprom.n2815 ));
    Odrv4 I__3998 (
            .O(N__20832),
            .I(\eeprom.n2815 ));
    LocalMux I__3997 (
            .O(N__20829),
            .I(\eeprom.n2815 ));
    InMux I__3996 (
            .O(N__20822),
            .I(\eeprom.n4059 ));
    CascadeMux I__3995 (
            .O(N__20819),
            .I(N__20816));
    InMux I__3994 (
            .O(N__20816),
            .I(N__20812));
    CascadeMux I__3993 (
            .O(N__20815),
            .I(N__20809));
    LocalMux I__3992 (
            .O(N__20812),
            .I(N__20806));
    InMux I__3991 (
            .O(N__20809),
            .I(N__20803));
    Span4Mux_h I__3990 (
            .O(N__20806),
            .I(N__20797));
    LocalMux I__3989 (
            .O(N__20803),
            .I(N__20797));
    InMux I__3988 (
            .O(N__20802),
            .I(N__20794));
    Odrv4 I__3987 (
            .O(N__20797),
            .I(\eeprom.n2814 ));
    LocalMux I__3986 (
            .O(N__20794),
            .I(\eeprom.n2814 ));
    InMux I__3985 (
            .O(N__20789),
            .I(\eeprom.n4060 ));
    CascadeMux I__3984 (
            .O(N__20786),
            .I(N__20782));
    InMux I__3983 (
            .O(N__20785),
            .I(N__20779));
    InMux I__3982 (
            .O(N__20782),
            .I(N__20775));
    LocalMux I__3981 (
            .O(N__20779),
            .I(N__20772));
    InMux I__3980 (
            .O(N__20778),
            .I(N__20769));
    LocalMux I__3979 (
            .O(N__20775),
            .I(\eeprom.n2813 ));
    Odrv4 I__3978 (
            .O(N__20772),
            .I(\eeprom.n2813 ));
    LocalMux I__3977 (
            .O(N__20769),
            .I(\eeprom.n2813 ));
    InMux I__3976 (
            .O(N__20762),
            .I(\eeprom.n4061 ));
    CascadeMux I__3975 (
            .O(N__20759),
            .I(N__20751));
    CascadeMux I__3974 (
            .O(N__20758),
            .I(N__20748));
    CascadeMux I__3973 (
            .O(N__20757),
            .I(N__20745));
    CascadeMux I__3972 (
            .O(N__20756),
            .I(N__20742));
    CascadeMux I__3971 (
            .O(N__20755),
            .I(N__20739));
    CascadeMux I__3970 (
            .O(N__20754),
            .I(N__20736));
    InMux I__3969 (
            .O(N__20751),
            .I(N__20731));
    InMux I__3968 (
            .O(N__20748),
            .I(N__20731));
    InMux I__3967 (
            .O(N__20745),
            .I(N__20722));
    InMux I__3966 (
            .O(N__20742),
            .I(N__20722));
    InMux I__3965 (
            .O(N__20739),
            .I(N__20722));
    InMux I__3964 (
            .O(N__20736),
            .I(N__20722));
    LocalMux I__3963 (
            .O(N__20731),
            .I(\eeprom.n5575 ));
    LocalMux I__3962 (
            .O(N__20722),
            .I(\eeprom.n5575 ));
    CascadeMux I__3961 (
            .O(N__20717),
            .I(N__20714));
    InMux I__3960 (
            .O(N__20714),
            .I(N__20711));
    LocalMux I__3959 (
            .O(N__20711),
            .I(N__20706));
    InMux I__3958 (
            .O(N__20710),
            .I(N__20701));
    InMux I__3957 (
            .O(N__20709),
            .I(N__20701));
    Odrv4 I__3956 (
            .O(N__20706),
            .I(\eeprom.n2812 ));
    LocalMux I__3955 (
            .O(N__20701),
            .I(\eeprom.n2812 ));
    InMux I__3954 (
            .O(N__20696),
            .I(\eeprom.n4062 ));
    InMux I__3953 (
            .O(N__20693),
            .I(N__20688));
    InMux I__3952 (
            .O(N__20692),
            .I(N__20685));
    InMux I__3951 (
            .O(N__20691),
            .I(N__20682));
    LocalMux I__3950 (
            .O(N__20688),
            .I(\eeprom.n2712 ));
    LocalMux I__3949 (
            .O(N__20685),
            .I(\eeprom.n2712 ));
    LocalMux I__3948 (
            .O(N__20682),
            .I(\eeprom.n2712 ));
    CascadeMux I__3947 (
            .O(N__20675),
            .I(\eeprom.n2638_cascade_ ));
    InMux I__3946 (
            .O(N__20672),
            .I(N__20669));
    LocalMux I__3945 (
            .O(N__20669),
            .I(\eeprom.n2684 ));
    CascadeMux I__3944 (
            .O(N__20666),
            .I(\eeprom.n2716_cascade_ ));
    CascadeMux I__3943 (
            .O(N__20663),
            .I(N__20660));
    InMux I__3942 (
            .O(N__20660),
            .I(N__20657));
    LocalMux I__3941 (
            .O(N__20657),
            .I(\eeprom.n2680 ));
    InMux I__3940 (
            .O(N__20654),
            .I(N__20651));
    LocalMux I__3939 (
            .O(N__20651),
            .I(\eeprom.n2679 ));
    CascadeMux I__3938 (
            .O(N__20648),
            .I(N__20645));
    InMux I__3937 (
            .O(N__20645),
            .I(N__20642));
    LocalMux I__3936 (
            .O(N__20642),
            .I(\eeprom.n2676 ));
    InMux I__3935 (
            .O(N__20639),
            .I(N__20636));
    LocalMux I__3934 (
            .O(N__20636),
            .I(\eeprom.n2675 ));
    CascadeMux I__3933 (
            .O(N__20633),
            .I(N__20630));
    InMux I__3932 (
            .O(N__20630),
            .I(N__20627));
    LocalMux I__3931 (
            .O(N__20627),
            .I(\eeprom.n2673 ));
    CascadeMux I__3930 (
            .O(N__20624),
            .I(\eeprom.n2705_cascade_ ));
    InMux I__3929 (
            .O(N__20621),
            .I(N__20618));
    LocalMux I__3928 (
            .O(N__20618),
            .I(\eeprom.n17_adj_339 ));
    CascadeMux I__3927 (
            .O(N__20615),
            .I(\eeprom.n16_adj_338_cascade_ ));
    InMux I__3926 (
            .O(N__20612),
            .I(N__20609));
    LocalMux I__3925 (
            .O(N__20609),
            .I(N__20604));
    InMux I__3924 (
            .O(N__20608),
            .I(N__20599));
    InMux I__3923 (
            .O(N__20607),
            .I(N__20599));
    Odrv4 I__3922 (
            .O(N__20604),
            .I(\eeprom.n2413 ));
    LocalMux I__3921 (
            .O(N__20599),
            .I(\eeprom.n2413 ));
    CascadeMux I__3920 (
            .O(N__20594),
            .I(N__20591));
    InMux I__3919 (
            .O(N__20591),
            .I(N__20588));
    LocalMux I__3918 (
            .O(N__20588),
            .I(\eeprom.n2480 ));
    InMux I__3917 (
            .O(N__20585),
            .I(\eeprom.n4023 ));
    InMux I__3916 (
            .O(N__20582),
            .I(N__20578));
    InMux I__3915 (
            .O(N__20581),
            .I(N__20574));
    LocalMux I__3914 (
            .O(N__20578),
            .I(N__20571));
    InMux I__3913 (
            .O(N__20577),
            .I(N__20568));
    LocalMux I__3912 (
            .O(N__20574),
            .I(N__20565));
    Odrv4 I__3911 (
            .O(N__20571),
            .I(\eeprom.n2412 ));
    LocalMux I__3910 (
            .O(N__20568),
            .I(\eeprom.n2412 ));
    Odrv4 I__3909 (
            .O(N__20565),
            .I(\eeprom.n2412 ));
    CascadeMux I__3908 (
            .O(N__20558),
            .I(N__20555));
    InMux I__3907 (
            .O(N__20555),
            .I(N__20552));
    LocalMux I__3906 (
            .O(N__20552),
            .I(\eeprom.n2479 ));
    InMux I__3905 (
            .O(N__20549),
            .I(\eeprom.n4024 ));
    InMux I__3904 (
            .O(N__20546),
            .I(bfn_22_23_0_));
    InMux I__3903 (
            .O(N__20543),
            .I(\eeprom.n4026 ));
    InMux I__3902 (
            .O(N__20540),
            .I(N__20537));
    LocalMux I__3901 (
            .O(N__20537),
            .I(N__20532));
    InMux I__3900 (
            .O(N__20536),
            .I(N__20527));
    InMux I__3899 (
            .O(N__20535),
            .I(N__20527));
    Odrv4 I__3898 (
            .O(N__20532),
            .I(\eeprom.n2409 ));
    LocalMux I__3897 (
            .O(N__20527),
            .I(\eeprom.n2409 ));
    InMux I__3896 (
            .O(N__20522),
            .I(N__20519));
    LocalMux I__3895 (
            .O(N__20519),
            .I(N__20516));
    Odrv4 I__3894 (
            .O(N__20516),
            .I(\eeprom.n2476 ));
    InMux I__3893 (
            .O(N__20513),
            .I(\eeprom.n4027 ));
    InMux I__3892 (
            .O(N__20510),
            .I(\eeprom.n4028 ));
    CascadeMux I__3891 (
            .O(N__20507),
            .I(N__20504));
    InMux I__3890 (
            .O(N__20504),
            .I(N__20501));
    LocalMux I__3889 (
            .O(N__20501),
            .I(N__20497));
    InMux I__3888 (
            .O(N__20500),
            .I(N__20494));
    Odrv4 I__3887 (
            .O(N__20497),
            .I(\eeprom.n2407 ));
    LocalMux I__3886 (
            .O(N__20494),
            .I(\eeprom.n2407 ));
    InMux I__3885 (
            .O(N__20489),
            .I(\eeprom.n4029 ));
    CascadeMux I__3884 (
            .O(N__20486),
            .I(\eeprom.n2440_cascade_ ));
    InMux I__3883 (
            .O(N__20483),
            .I(N__20480));
    LocalMux I__3882 (
            .O(N__20480),
            .I(\eeprom.n5071 ));
    InMux I__3881 (
            .O(N__20477),
            .I(bfn_22_22_0_));
    InMux I__3880 (
            .O(N__20474),
            .I(\eeprom.n4018 ));
    InMux I__3879 (
            .O(N__20471),
            .I(\eeprom.n4019 ));
    InMux I__3878 (
            .O(N__20468),
            .I(\eeprom.n4020 ));
    InMux I__3877 (
            .O(N__20465),
            .I(\eeprom.n4021 ));
    CascadeMux I__3876 (
            .O(N__20462),
            .I(N__20459));
    InMux I__3875 (
            .O(N__20459),
            .I(N__20456));
    LocalMux I__3874 (
            .O(N__20456),
            .I(N__20451));
    InMux I__3873 (
            .O(N__20455),
            .I(N__20446));
    InMux I__3872 (
            .O(N__20454),
            .I(N__20446));
    Odrv4 I__3871 (
            .O(N__20451),
            .I(\eeprom.n2414 ));
    LocalMux I__3870 (
            .O(N__20446),
            .I(\eeprom.n2414 ));
    InMux I__3869 (
            .O(N__20441),
            .I(N__20438));
    LocalMux I__3868 (
            .O(N__20438),
            .I(\eeprom.n2481 ));
    InMux I__3867 (
            .O(N__20435),
            .I(\eeprom.n4022 ));
    CascadeMux I__3866 (
            .O(N__20432),
            .I(\eeprom.n2309_cascade_ ));
    InMux I__3865 (
            .O(N__20429),
            .I(N__20425));
    InMux I__3864 (
            .O(N__20428),
            .I(N__20422));
    LocalMux I__3863 (
            .O(N__20425),
            .I(N__20416));
    LocalMux I__3862 (
            .O(N__20422),
            .I(N__20416));
    InMux I__3861 (
            .O(N__20421),
            .I(N__20413));
    Span4Mux_h I__3860 (
            .O(N__20416),
            .I(N__20408));
    LocalMux I__3859 (
            .O(N__20413),
            .I(N__20408));
    Odrv4 I__3858 (
            .O(N__20408),
            .I(\eeprom.n2308 ));
    InMux I__3857 (
            .O(N__20405),
            .I(N__20401));
    InMux I__3856 (
            .O(N__20404),
            .I(N__20398));
    LocalMux I__3855 (
            .O(N__20401),
            .I(N__20393));
    LocalMux I__3854 (
            .O(N__20398),
            .I(N__20393));
    Span4Mux_v I__3853 (
            .O(N__20393),
            .I(N__20389));
    InMux I__3852 (
            .O(N__20392),
            .I(N__20386));
    Odrv4 I__3851 (
            .O(N__20389),
            .I(\eeprom.n2312 ));
    LocalMux I__3850 (
            .O(N__20386),
            .I(\eeprom.n2312 ));
    CascadeMux I__3849 (
            .O(N__20381),
            .I(\eeprom.n8_adj_322_cascade_ ));
    InMux I__3848 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__3847 (
            .O(N__20375),
            .I(\eeprom.n7_adj_323 ));
    CascadeMux I__3846 (
            .O(N__20372),
            .I(N__20364));
    CascadeMux I__3845 (
            .O(N__20371),
            .I(N__20361));
    CascadeMux I__3844 (
            .O(N__20370),
            .I(N__20358));
    CascadeMux I__3843 (
            .O(N__20369),
            .I(N__20355));
    CascadeMux I__3842 (
            .O(N__20368),
            .I(N__20352));
    CascadeMux I__3841 (
            .O(N__20367),
            .I(N__20349));
    InMux I__3840 (
            .O(N__20364),
            .I(N__20344));
    InMux I__3839 (
            .O(N__20361),
            .I(N__20344));
    InMux I__3838 (
            .O(N__20358),
            .I(N__20339));
    InMux I__3837 (
            .O(N__20355),
            .I(N__20339));
    InMux I__3836 (
            .O(N__20352),
            .I(N__20334));
    InMux I__3835 (
            .O(N__20349),
            .I(N__20334));
    LocalMux I__3834 (
            .O(N__20344),
            .I(\eeprom.n2341 ));
    LocalMux I__3833 (
            .O(N__20339),
            .I(\eeprom.n2341 ));
    LocalMux I__3832 (
            .O(N__20334),
            .I(\eeprom.n2341 ));
    CascadeMux I__3831 (
            .O(N__20327),
            .I(\eeprom.n2341_cascade_ ));
    CascadeMux I__3830 (
            .O(N__20324),
            .I(N__20316));
    CascadeMux I__3829 (
            .O(N__20323),
            .I(N__20313));
    CascadeMux I__3828 (
            .O(N__20322),
            .I(N__20310));
    CascadeMux I__3827 (
            .O(N__20321),
            .I(N__20307));
    CascadeMux I__3826 (
            .O(N__20320),
            .I(N__20304));
    CascadeMux I__3825 (
            .O(N__20319),
            .I(N__20301));
    InMux I__3824 (
            .O(N__20316),
            .I(N__20296));
    InMux I__3823 (
            .O(N__20313),
            .I(N__20296));
    InMux I__3822 (
            .O(N__20310),
            .I(N__20287));
    InMux I__3821 (
            .O(N__20307),
            .I(N__20287));
    InMux I__3820 (
            .O(N__20304),
            .I(N__20287));
    InMux I__3819 (
            .O(N__20301),
            .I(N__20287));
    LocalMux I__3818 (
            .O(N__20296),
            .I(\eeprom.n5576 ));
    LocalMux I__3817 (
            .O(N__20287),
            .I(\eeprom.n5576 ));
    InMux I__3816 (
            .O(N__20282),
            .I(N__20279));
    LocalMux I__3815 (
            .O(N__20279),
            .I(N__20276));
    Odrv4 I__3814 (
            .O(N__20276),
            .I(\eeprom.n2279 ));
    InMux I__3813 (
            .O(N__20273),
            .I(N__20268));
    InMux I__3812 (
            .O(N__20272),
            .I(N__20265));
    InMux I__3811 (
            .O(N__20271),
            .I(N__20262));
    LocalMux I__3810 (
            .O(N__20268),
            .I(\eeprom.n2311 ));
    LocalMux I__3809 (
            .O(N__20265),
            .I(\eeprom.n2311 ));
    LocalMux I__3808 (
            .O(N__20262),
            .I(\eeprom.n2311 ));
    CascadeMux I__3807 (
            .O(N__20255),
            .I(\eeprom.n5073_cascade_ ));
    CascadeMux I__3806 (
            .O(N__20252),
            .I(\eeprom.n4782_cascade_ ));
    CascadeMux I__3805 (
            .O(N__20249),
            .I(\eeprom.n12_cascade_ ));
    CascadeMux I__3804 (
            .O(N__20246),
            .I(\eeprom.n2242_cascade_ ));
    InMux I__3803 (
            .O(N__20243),
            .I(N__20240));
    LocalMux I__3802 (
            .O(N__20240),
            .I(N__20237));
    Odrv4 I__3801 (
            .O(N__20237),
            .I(\eeprom.n2282 ));
    CascadeMux I__3800 (
            .O(N__20234),
            .I(\eeprom.n5400_cascade_ ));
    CascadeMux I__3799 (
            .O(N__20231),
            .I(N__20227));
    InMux I__3798 (
            .O(N__20230),
            .I(N__20223));
    InMux I__3797 (
            .O(N__20227),
            .I(N__20220));
    InMux I__3796 (
            .O(N__20226),
            .I(N__20217));
    LocalMux I__3795 (
            .O(N__20223),
            .I(\eeprom.n2217 ));
    LocalMux I__3794 (
            .O(N__20220),
            .I(\eeprom.n2217 ));
    LocalMux I__3793 (
            .O(N__20217),
            .I(\eeprom.n2217 ));
    CascadeMux I__3792 (
            .O(N__20210),
            .I(N__20207));
    InMux I__3791 (
            .O(N__20207),
            .I(N__20204));
    LocalMux I__3790 (
            .O(N__20204),
            .I(N__20201));
    Odrv4 I__3789 (
            .O(N__20201),
            .I(\eeprom.n2284 ));
    InMux I__3788 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__3787 (
            .O(N__20195),
            .I(N__20192));
    Odrv4 I__3786 (
            .O(N__20192),
            .I(\eeprom.n2280 ));
    CascadeMux I__3785 (
            .O(N__20189),
            .I(N__20186));
    InMux I__3784 (
            .O(N__20186),
            .I(N__20181));
    InMux I__3783 (
            .O(N__20185),
            .I(N__20176));
    InMux I__3782 (
            .O(N__20184),
            .I(N__20176));
    LocalMux I__3781 (
            .O(N__20181),
            .I(\eeprom.n2213 ));
    LocalMux I__3780 (
            .O(N__20176),
            .I(\eeprom.n2213 ));
    InMux I__3779 (
            .O(N__20171),
            .I(N__20168));
    LocalMux I__3778 (
            .O(N__20168),
            .I(\eeprom.n5405 ));
    InMux I__3777 (
            .O(N__20165),
            .I(N__20160));
    InMux I__3776 (
            .O(N__20164),
            .I(N__20157));
    InMux I__3775 (
            .O(N__20163),
            .I(N__20154));
    LocalMux I__3774 (
            .O(N__20160),
            .I(\eeprom.n2316 ));
    LocalMux I__3773 (
            .O(N__20157),
            .I(\eeprom.n2316 ));
    LocalMux I__3772 (
            .O(N__20154),
            .I(\eeprom.n2316 ));
    InMux I__3771 (
            .O(N__20147),
            .I(N__20142));
    InMux I__3770 (
            .O(N__20146),
            .I(N__20139));
    InMux I__3769 (
            .O(N__20145),
            .I(N__20136));
    LocalMux I__3768 (
            .O(N__20142),
            .I(\eeprom.n2317 ));
    LocalMux I__3767 (
            .O(N__20139),
            .I(\eeprom.n2317 ));
    LocalMux I__3766 (
            .O(N__20136),
            .I(\eeprom.n2317 ));
    CascadeMux I__3765 (
            .O(N__20129),
            .I(N__20124));
    InMux I__3764 (
            .O(N__20128),
            .I(N__20121));
    InMux I__3763 (
            .O(N__20127),
            .I(N__20118));
    InMux I__3762 (
            .O(N__20124),
            .I(N__20115));
    LocalMux I__3761 (
            .O(N__20121),
            .I(\eeprom.n2314 ));
    LocalMux I__3760 (
            .O(N__20118),
            .I(\eeprom.n2314 ));
    LocalMux I__3759 (
            .O(N__20115),
            .I(\eeprom.n2314 ));
    InMux I__3758 (
            .O(N__20108),
            .I(N__20103));
    InMux I__3757 (
            .O(N__20107),
            .I(N__20100));
    InMux I__3756 (
            .O(N__20106),
            .I(N__20097));
    LocalMux I__3755 (
            .O(N__20103),
            .I(\eeprom.n2318 ));
    LocalMux I__3754 (
            .O(N__20100),
            .I(\eeprom.n2318 ));
    LocalMux I__3753 (
            .O(N__20097),
            .I(\eeprom.n2318 ));
    CascadeMux I__3752 (
            .O(N__20090),
            .I(\eeprom.n5085_cascade_ ));
    InMux I__3751 (
            .O(N__20087),
            .I(N__20082));
    InMux I__3750 (
            .O(N__20086),
            .I(N__20079));
    InMux I__3749 (
            .O(N__20085),
            .I(N__20076));
    LocalMux I__3748 (
            .O(N__20082),
            .I(N__20071));
    LocalMux I__3747 (
            .O(N__20079),
            .I(N__20071));
    LocalMux I__3746 (
            .O(N__20076),
            .I(N__20068));
    Odrv12 I__3745 (
            .O(N__20071),
            .I(\eeprom.n2310 ));
    Odrv4 I__3744 (
            .O(N__20068),
            .I(\eeprom.n2310 ));
    CascadeMux I__3743 (
            .O(N__20063),
            .I(N__20058));
    InMux I__3742 (
            .O(N__20062),
            .I(N__20055));
    InMux I__3741 (
            .O(N__20061),
            .I(N__20052));
    InMux I__3740 (
            .O(N__20058),
            .I(N__20049));
    LocalMux I__3739 (
            .O(N__20055),
            .I(\eeprom.n2315 ));
    LocalMux I__3738 (
            .O(N__20052),
            .I(\eeprom.n2315 ));
    LocalMux I__3737 (
            .O(N__20049),
            .I(\eeprom.n2315 ));
    InMux I__3736 (
            .O(N__20042),
            .I(N__20037));
    InMux I__3735 (
            .O(N__20041),
            .I(N__20034));
    InMux I__3734 (
            .O(N__20040),
            .I(N__20031));
    LocalMux I__3733 (
            .O(N__20037),
            .I(\eeprom.n2313 ));
    LocalMux I__3732 (
            .O(N__20034),
            .I(\eeprom.n2313 ));
    LocalMux I__3731 (
            .O(N__20031),
            .I(\eeprom.n2313 ));
    InMux I__3730 (
            .O(N__20024),
            .I(N__20021));
    LocalMux I__3729 (
            .O(N__20021),
            .I(\eeprom.n5081 ));
    InMux I__3728 (
            .O(N__20018),
            .I(N__20015));
    LocalMux I__3727 (
            .O(N__20015),
            .I(N__20012));
    Odrv12 I__3726 (
            .O(N__20012),
            .I(\eeprom.n2277 ));
    InMux I__3725 (
            .O(N__20009),
            .I(N__20005));
    InMux I__3724 (
            .O(N__20008),
            .I(N__20002));
    LocalMux I__3723 (
            .O(N__20005),
            .I(\eeprom.n2309 ));
    LocalMux I__3722 (
            .O(N__20002),
            .I(\eeprom.n2309 ));
    InMux I__3721 (
            .O(N__19997),
            .I(\eeprom.n4005 ));
    InMux I__3720 (
            .O(N__19994),
            .I(\eeprom.n4006 ));
    CascadeMux I__3719 (
            .O(N__19991),
            .I(N__19987));
    CascadeMux I__3718 (
            .O(N__19990),
            .I(N__19984));
    InMux I__3717 (
            .O(N__19987),
            .I(N__19980));
    InMux I__3716 (
            .O(N__19984),
            .I(N__19977));
    InMux I__3715 (
            .O(N__19983),
            .I(N__19974));
    LocalMux I__3714 (
            .O(N__19980),
            .I(\eeprom.n2216 ));
    LocalMux I__3713 (
            .O(N__19977),
            .I(\eeprom.n2216 ));
    LocalMux I__3712 (
            .O(N__19974),
            .I(\eeprom.n2216 ));
    CascadeMux I__3711 (
            .O(N__19967),
            .I(\eeprom.n2143_cascade_ ));
    InMux I__3710 (
            .O(N__19964),
            .I(N__19961));
    LocalMux I__3709 (
            .O(N__19961),
            .I(N__19958));
    Odrv4 I__3708 (
            .O(N__19958),
            .I(\eeprom.n2286 ));
    InMux I__3707 (
            .O(N__19955),
            .I(N__19951));
    CascadeMux I__3706 (
            .O(N__19954),
            .I(N__19947));
    LocalMux I__3705 (
            .O(N__19951),
            .I(N__19944));
    InMux I__3704 (
            .O(N__19950),
            .I(N__19941));
    InMux I__3703 (
            .O(N__19947),
            .I(N__19938));
    Odrv4 I__3702 (
            .O(N__19944),
            .I(\eeprom.n2218 ));
    LocalMux I__3701 (
            .O(N__19941),
            .I(\eeprom.n2218 ));
    LocalMux I__3700 (
            .O(N__19938),
            .I(\eeprom.n2218 ));
    InMux I__3699 (
            .O(N__19931),
            .I(N__19928));
    LocalMux I__3698 (
            .O(N__19928),
            .I(\eeprom.n5045 ));
    CascadeMux I__3697 (
            .O(N__19925),
            .I(N__19922));
    InMux I__3696 (
            .O(N__19922),
            .I(N__19918));
    InMux I__3695 (
            .O(N__19921),
            .I(N__19915));
    LocalMux I__3694 (
            .O(N__19918),
            .I(\eeprom.n2211 ));
    LocalMux I__3693 (
            .O(N__19915),
            .I(\eeprom.n2211 ));
    CascadeMux I__3692 (
            .O(N__19910),
            .I(\eeprom.n4797_cascade_ ));
    InMux I__3691 (
            .O(N__19907),
            .I(N__19904));
    LocalMux I__3690 (
            .O(N__19904),
            .I(N__19901));
    Span4Mux_h I__3689 (
            .O(N__19901),
            .I(N__19898));
    Odrv4 I__3688 (
            .O(N__19898),
            .I(\eeprom.n2285 ));
    InMux I__3687 (
            .O(N__19895),
            .I(\eeprom.n3997 ));
    InMux I__3686 (
            .O(N__19892),
            .I(\eeprom.n3998 ));
    InMux I__3685 (
            .O(N__19889),
            .I(N__19886));
    LocalMux I__3684 (
            .O(N__19886),
            .I(N__19883));
    Odrv4 I__3683 (
            .O(N__19883),
            .I(\eeprom.n2283 ));
    InMux I__3682 (
            .O(N__19880),
            .I(\eeprom.n3999 ));
    CascadeMux I__3681 (
            .O(N__19877),
            .I(N__19874));
    InMux I__3680 (
            .O(N__19874),
            .I(N__19870));
    InMux I__3679 (
            .O(N__19873),
            .I(N__19867));
    LocalMux I__3678 (
            .O(N__19870),
            .I(\eeprom.n2215 ));
    LocalMux I__3677 (
            .O(N__19867),
            .I(\eeprom.n2215 ));
    InMux I__3676 (
            .O(N__19862),
            .I(\eeprom.n4000 ));
    CascadeMux I__3675 (
            .O(N__19859),
            .I(N__19856));
    InMux I__3674 (
            .O(N__19856),
            .I(N__19852));
    InMux I__3673 (
            .O(N__19855),
            .I(N__19849));
    LocalMux I__3672 (
            .O(N__19852),
            .I(N__19846));
    LocalMux I__3671 (
            .O(N__19849),
            .I(\eeprom.n2214 ));
    Odrv4 I__3670 (
            .O(N__19846),
            .I(\eeprom.n2214 ));
    CascadeMux I__3669 (
            .O(N__19841),
            .I(N__19838));
    InMux I__3668 (
            .O(N__19838),
            .I(N__19835));
    LocalMux I__3667 (
            .O(N__19835),
            .I(N__19832));
    Odrv4 I__3666 (
            .O(N__19832),
            .I(\eeprom.n2281 ));
    InMux I__3665 (
            .O(N__19829),
            .I(\eeprom.n4001 ));
    InMux I__3664 (
            .O(N__19826),
            .I(\eeprom.n4002 ));
    InMux I__3663 (
            .O(N__19823),
            .I(\eeprom.n4003 ));
    InMux I__3662 (
            .O(N__19820),
            .I(N__19817));
    LocalMux I__3661 (
            .O(N__19817),
            .I(\eeprom.n2278 ));
    InMux I__3660 (
            .O(N__19814),
            .I(bfn_22_18_0_));
    InMux I__3659 (
            .O(N__19811),
            .I(\eeprom.n4085 ));
    InMux I__3658 (
            .O(N__19808),
            .I(\eeprom.n4086 ));
    InMux I__3657 (
            .O(N__19805),
            .I(bfn_21_29_0_));
    InMux I__3656 (
            .O(N__19802),
            .I(N__19799));
    LocalMux I__3655 (
            .O(N__19799),
            .I(N__19796));
    Odrv4 I__3654 (
            .O(N__19796),
            .I(\eeprom.n2902 ));
    CascadeMux I__3653 (
            .O(N__19793),
            .I(\eeprom.n2902_cascade_ ));
    InMux I__3652 (
            .O(N__19790),
            .I(N__19787));
    LocalMux I__3651 (
            .O(N__19787),
            .I(N__19784));
    Odrv4 I__3650 (
            .O(N__19784),
            .I(\eeprom.n19_adj_327 ));
    InMux I__3649 (
            .O(N__19781),
            .I(N__19778));
    LocalMux I__3648 (
            .O(N__19778),
            .I(\eeprom.n2872 ));
    InMux I__3647 (
            .O(N__19775),
            .I(N__19772));
    LocalMux I__3646 (
            .O(N__19772),
            .I(N__19767));
    InMux I__3645 (
            .O(N__19771),
            .I(N__19764));
    InMux I__3644 (
            .O(N__19770),
            .I(N__19761));
    Odrv4 I__3643 (
            .O(N__19767),
            .I(\eeprom.n2904 ));
    LocalMux I__3642 (
            .O(N__19764),
            .I(\eeprom.n2904 ));
    LocalMux I__3641 (
            .O(N__19761),
            .I(\eeprom.n2904 ));
    InMux I__3640 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__3639 (
            .O(N__19751),
            .I(\eeprom.n2873 ));
    InMux I__3638 (
            .O(N__19748),
            .I(N__19745));
    LocalMux I__3637 (
            .O(N__19745),
            .I(N__19742));
    Span4Mux_s3_v I__3636 (
            .O(N__19742),
            .I(N__19737));
    InMux I__3635 (
            .O(N__19741),
            .I(N__19734));
    InMux I__3634 (
            .O(N__19740),
            .I(N__19731));
    Odrv4 I__3633 (
            .O(N__19737),
            .I(\eeprom.n2905 ));
    LocalMux I__3632 (
            .O(N__19734),
            .I(\eeprom.n2905 ));
    LocalMux I__3631 (
            .O(N__19731),
            .I(\eeprom.n2905 ));
    InMux I__3630 (
            .O(N__19724),
            .I(N__19721));
    LocalMux I__3629 (
            .O(N__19721),
            .I(\eeprom.n2871 ));
    InMux I__3628 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__3627 (
            .O(N__19715),
            .I(N__19711));
    InMux I__3626 (
            .O(N__19714),
            .I(N__19708));
    Span4Mux_v I__3625 (
            .O(N__19711),
            .I(N__19704));
    LocalMux I__3624 (
            .O(N__19708),
            .I(N__19701));
    InMux I__3623 (
            .O(N__19707),
            .I(N__19698));
    Odrv4 I__3622 (
            .O(N__19704),
            .I(\eeprom.n2903 ));
    Odrv4 I__3621 (
            .O(N__19701),
            .I(\eeprom.n2903 ));
    LocalMux I__3620 (
            .O(N__19698),
            .I(\eeprom.n2903 ));
    CascadeMux I__3619 (
            .O(N__19691),
            .I(N__19688));
    InMux I__3618 (
            .O(N__19688),
            .I(N__19685));
    LocalMux I__3617 (
            .O(N__19685),
            .I(\eeprom.n2875 ));
    CascadeMux I__3616 (
            .O(N__19682),
            .I(N__19675));
    InMux I__3615 (
            .O(N__19681),
            .I(N__19667));
    CascadeMux I__3614 (
            .O(N__19680),
            .I(N__19663));
    CascadeMux I__3613 (
            .O(N__19679),
            .I(N__19660));
    CascadeMux I__3612 (
            .O(N__19678),
            .I(N__19657));
    InMux I__3611 (
            .O(N__19675),
            .I(N__19651));
    InMux I__3610 (
            .O(N__19674),
            .I(N__19651));
    CascadeMux I__3609 (
            .O(N__19673),
            .I(N__19648));
    CascadeMux I__3608 (
            .O(N__19672),
            .I(N__19645));
    CascadeMux I__3607 (
            .O(N__19671),
            .I(N__19639));
    InMux I__3606 (
            .O(N__19670),
            .I(N__19635));
    LocalMux I__3605 (
            .O(N__19667),
            .I(N__19632));
    InMux I__3604 (
            .O(N__19666),
            .I(N__19621));
    InMux I__3603 (
            .O(N__19663),
            .I(N__19621));
    InMux I__3602 (
            .O(N__19660),
            .I(N__19621));
    InMux I__3601 (
            .O(N__19657),
            .I(N__19621));
    InMux I__3600 (
            .O(N__19656),
            .I(N__19621));
    LocalMux I__3599 (
            .O(N__19651),
            .I(N__19618));
    InMux I__3598 (
            .O(N__19648),
            .I(N__19609));
    InMux I__3597 (
            .O(N__19645),
            .I(N__19609));
    InMux I__3596 (
            .O(N__19644),
            .I(N__19609));
    InMux I__3595 (
            .O(N__19643),
            .I(N__19609));
    InMux I__3594 (
            .O(N__19642),
            .I(N__19602));
    InMux I__3593 (
            .O(N__19639),
            .I(N__19602));
    InMux I__3592 (
            .O(N__19638),
            .I(N__19602));
    LocalMux I__3591 (
            .O(N__19635),
            .I(\eeprom.n2836 ));
    Odrv4 I__3590 (
            .O(N__19632),
            .I(\eeprom.n2836 ));
    LocalMux I__3589 (
            .O(N__19621),
            .I(\eeprom.n2836 ));
    Odrv4 I__3588 (
            .O(N__19618),
            .I(\eeprom.n2836 ));
    LocalMux I__3587 (
            .O(N__19609),
            .I(\eeprom.n2836 ));
    LocalMux I__3586 (
            .O(N__19602),
            .I(\eeprom.n2836 ));
    InMux I__3585 (
            .O(N__19589),
            .I(N__19585));
    InMux I__3584 (
            .O(N__19588),
            .I(N__19582));
    LocalMux I__3583 (
            .O(N__19585),
            .I(N__19579));
    LocalMux I__3582 (
            .O(N__19582),
            .I(N__19575));
    Span4Mux_h I__3581 (
            .O(N__19579),
            .I(N__19572));
    InMux I__3580 (
            .O(N__19578),
            .I(N__19569));
    Span4Mux_h I__3579 (
            .O(N__19575),
            .I(N__19566));
    Odrv4 I__3578 (
            .O(N__19572),
            .I(\eeprom.n2907 ));
    LocalMux I__3577 (
            .O(N__19569),
            .I(\eeprom.n2907 ));
    Odrv4 I__3576 (
            .O(N__19566),
            .I(\eeprom.n2907 ));
    InMux I__3575 (
            .O(N__19559),
            .I(bfn_22_17_0_));
    InMux I__3574 (
            .O(N__19556),
            .I(N__19553));
    LocalMux I__3573 (
            .O(N__19553),
            .I(N__19550));
    Odrv4 I__3572 (
            .O(N__19550),
            .I(\eeprom.n2880 ));
    InMux I__3571 (
            .O(N__19547),
            .I(\eeprom.n4077 ));
    InMux I__3570 (
            .O(N__19544),
            .I(N__19541));
    LocalMux I__3569 (
            .O(N__19541),
            .I(\eeprom.n2879 ));
    InMux I__3568 (
            .O(N__19538),
            .I(\eeprom.n4078 ));
    InMux I__3567 (
            .O(N__19535),
            .I(N__19532));
    LocalMux I__3566 (
            .O(N__19532),
            .I(\eeprom.n2878 ));
    InMux I__3565 (
            .O(N__19529),
            .I(bfn_21_28_0_));
    CascadeMux I__3564 (
            .O(N__19526),
            .I(N__19523));
    InMux I__3563 (
            .O(N__19523),
            .I(N__19520));
    LocalMux I__3562 (
            .O(N__19520),
            .I(\eeprom.n2877 ));
    InMux I__3561 (
            .O(N__19517),
            .I(\eeprom.n4080 ));
    InMux I__3560 (
            .O(N__19514),
            .I(N__19511));
    LocalMux I__3559 (
            .O(N__19511),
            .I(N__19508));
    Odrv4 I__3558 (
            .O(N__19508),
            .I(\eeprom.n2876 ));
    InMux I__3557 (
            .O(N__19505),
            .I(\eeprom.n4081 ));
    InMux I__3556 (
            .O(N__19502),
            .I(\eeprom.n4082 ));
    CascadeMux I__3555 (
            .O(N__19499),
            .I(N__19496));
    InMux I__3554 (
            .O(N__19496),
            .I(N__19493));
    LocalMux I__3553 (
            .O(N__19493),
            .I(\eeprom.n2874 ));
    InMux I__3552 (
            .O(N__19490),
            .I(\eeprom.n4083 ));
    InMux I__3551 (
            .O(N__19487),
            .I(\eeprom.n4084 ));
    InMux I__3550 (
            .O(N__19484),
            .I(N__19481));
    LocalMux I__3549 (
            .O(N__19481),
            .I(\eeprom.n5153 ));
    CascadeMux I__3548 (
            .O(N__19478),
            .I(N__19475));
    InMux I__3547 (
            .O(N__19475),
            .I(N__19470));
    CascadeMux I__3546 (
            .O(N__19474),
            .I(N__19467));
    InMux I__3545 (
            .O(N__19473),
            .I(N__19464));
    LocalMux I__3544 (
            .O(N__19470),
            .I(N__19461));
    InMux I__3543 (
            .O(N__19467),
            .I(N__19458));
    LocalMux I__3542 (
            .O(N__19464),
            .I(N__19455));
    Odrv12 I__3541 (
            .O(N__19461),
            .I(\eeprom.n2918 ));
    LocalMux I__3540 (
            .O(N__19458),
            .I(\eeprom.n2918 ));
    Odrv4 I__3539 (
            .O(N__19455),
            .I(\eeprom.n2918 ));
    InMux I__3538 (
            .O(N__19448),
            .I(N__19444));
    InMux I__3537 (
            .O(N__19447),
            .I(N__19441));
    LocalMux I__3536 (
            .O(N__19444),
            .I(N__19438));
    LocalMux I__3535 (
            .O(N__19441),
            .I(N__19435));
    Span4Mux_h I__3534 (
            .O(N__19438),
            .I(N__19429));
    Span4Mux_s3_v I__3533 (
            .O(N__19435),
            .I(N__19429));
    InMux I__3532 (
            .O(N__19434),
            .I(N__19426));
    Odrv4 I__3531 (
            .O(N__19429),
            .I(\eeprom.n2911 ));
    LocalMux I__3530 (
            .O(N__19426),
            .I(\eeprom.n2911 ));
    CascadeMux I__3529 (
            .O(N__19421),
            .I(N__19418));
    InMux I__3528 (
            .O(N__19418),
            .I(N__19415));
    LocalMux I__3527 (
            .O(N__19415),
            .I(\eeprom.n2886 ));
    InMux I__3526 (
            .O(N__19412),
            .I(bfn_21_27_0_));
    InMux I__3525 (
            .O(N__19409),
            .I(N__19406));
    LocalMux I__3524 (
            .O(N__19406),
            .I(\eeprom.n2885 ));
    InMux I__3523 (
            .O(N__19403),
            .I(\eeprom.n4072 ));
    CascadeMux I__3522 (
            .O(N__19400),
            .I(N__19397));
    InMux I__3521 (
            .O(N__19397),
            .I(N__19394));
    LocalMux I__3520 (
            .O(N__19394),
            .I(\eeprom.n2884 ));
    InMux I__3519 (
            .O(N__19391),
            .I(\eeprom.n4073 ));
    InMux I__3518 (
            .O(N__19388),
            .I(N__19385));
    LocalMux I__3517 (
            .O(N__19385),
            .I(\eeprom.n2883 ));
    InMux I__3516 (
            .O(N__19382),
            .I(\eeprom.n4074 ));
    CascadeMux I__3515 (
            .O(N__19379),
            .I(N__19376));
    InMux I__3514 (
            .O(N__19376),
            .I(N__19373));
    LocalMux I__3513 (
            .O(N__19373),
            .I(N__19370));
    Odrv4 I__3512 (
            .O(N__19370),
            .I(\eeprom.n2882 ));
    InMux I__3511 (
            .O(N__19367),
            .I(\eeprom.n4075 ));
    InMux I__3510 (
            .O(N__19364),
            .I(N__19361));
    LocalMux I__3509 (
            .O(N__19361),
            .I(\eeprom.n2881 ));
    InMux I__3508 (
            .O(N__19358),
            .I(\eeprom.n4076 ));
    InMux I__3507 (
            .O(N__19355),
            .I(\eeprom.n4055 ));
    InMux I__3506 (
            .O(N__19352),
            .I(\eeprom.n4056 ));
    InMux I__3505 (
            .O(N__19349),
            .I(N__19346));
    LocalMux I__3504 (
            .O(N__19346),
            .I(\eeprom.n2677 ));
    InMux I__3503 (
            .O(N__19343),
            .I(N__19340));
    LocalMux I__3502 (
            .O(N__19340),
            .I(\eeprom.n2678 ));
    CascadeMux I__3501 (
            .O(N__19337),
            .I(\eeprom.n2710_cascade_ ));
    InMux I__3500 (
            .O(N__19334),
            .I(N__19331));
    LocalMux I__3499 (
            .O(N__19331),
            .I(N__19328));
    Odrv4 I__3498 (
            .O(N__19328),
            .I(\eeprom.n2686 ));
    CascadeMux I__3497 (
            .O(N__19325),
            .I(N__19322));
    InMux I__3496 (
            .O(N__19322),
            .I(N__19319));
    LocalMux I__3495 (
            .O(N__19319),
            .I(N__19314));
    InMux I__3494 (
            .O(N__19318),
            .I(N__19309));
    InMux I__3493 (
            .O(N__19317),
            .I(N__19309));
    Span4Mux_v I__3492 (
            .O(N__19314),
            .I(N__19306));
    LocalMux I__3491 (
            .O(N__19309),
            .I(\eeprom.n2912 ));
    Odrv4 I__3490 (
            .O(N__19306),
            .I(\eeprom.n2912 ));
    CascadeMux I__3489 (
            .O(N__19301),
            .I(\eeprom.n5157_cascade_ ));
    InMux I__3488 (
            .O(N__19298),
            .I(N__19295));
    LocalMux I__3487 (
            .O(N__19295),
            .I(N__19292));
    Odrv4 I__3486 (
            .O(N__19292),
            .I(\eeprom.n16 ));
    InMux I__3485 (
            .O(N__19289),
            .I(\eeprom.n4046 ));
    InMux I__3484 (
            .O(N__19286),
            .I(\eeprom.n4047 ));
    InMux I__3483 (
            .O(N__19283),
            .I(\eeprom.n4048 ));
    InMux I__3482 (
            .O(N__19280),
            .I(\eeprom.n4049 ));
    InMux I__3481 (
            .O(N__19277),
            .I(bfn_21_24_0_));
    InMux I__3480 (
            .O(N__19274),
            .I(\eeprom.n4051 ));
    InMux I__3479 (
            .O(N__19271),
            .I(\eeprom.n4052 ));
    InMux I__3478 (
            .O(N__19268),
            .I(\eeprom.n4053 ));
    InMux I__3477 (
            .O(N__19265),
            .I(\eeprom.n4054 ));
    CascadeMux I__3476 (
            .O(N__19262),
            .I(N__19259));
    InMux I__3475 (
            .O(N__19259),
            .I(N__19255));
    InMux I__3474 (
            .O(N__19258),
            .I(N__19251));
    LocalMux I__3473 (
            .O(N__19255),
            .I(N__19248));
    InMux I__3472 (
            .O(N__19254),
            .I(N__19245));
    LocalMux I__3471 (
            .O(N__19251),
            .I(\eeprom.n3403 ));
    Odrv4 I__3470 (
            .O(N__19248),
            .I(\eeprom.n3403 ));
    LocalMux I__3469 (
            .O(N__19245),
            .I(\eeprom.n3403 ));
    CascadeMux I__3468 (
            .O(N__19238),
            .I(N__19235));
    InMux I__3467 (
            .O(N__19235),
            .I(N__19232));
    LocalMux I__3466 (
            .O(N__19232),
            .I(N__19229));
    Span4Mux_v I__3465 (
            .O(N__19229),
            .I(N__19226));
    Odrv4 I__3464 (
            .O(N__19226),
            .I(\eeprom.n3470 ));
    CascadeMux I__3463 (
            .O(N__19223),
            .I(N__19216));
    CascadeMux I__3462 (
            .O(N__19222),
            .I(N__19211));
    InMux I__3461 (
            .O(N__19221),
            .I(N__19208));
    CascadeMux I__3460 (
            .O(N__19220),
            .I(N__19200));
    CascadeMux I__3459 (
            .O(N__19219),
            .I(N__19197));
    InMux I__3458 (
            .O(N__19216),
            .I(N__19191));
    CascadeMux I__3457 (
            .O(N__19215),
            .I(N__19185));
    InMux I__3456 (
            .O(N__19214),
            .I(N__19180));
    InMux I__3455 (
            .O(N__19211),
            .I(N__19180));
    LocalMux I__3454 (
            .O(N__19208),
            .I(N__19177));
    InMux I__3453 (
            .O(N__19207),
            .I(N__19174));
    CascadeMux I__3452 (
            .O(N__19206),
            .I(N__19169));
    CascadeMux I__3451 (
            .O(N__19205),
            .I(N__19165));
    CascadeMux I__3450 (
            .O(N__19204),
            .I(N__19162));
    CascadeMux I__3449 (
            .O(N__19203),
            .I(N__19158));
    InMux I__3448 (
            .O(N__19200),
            .I(N__19151));
    InMux I__3447 (
            .O(N__19197),
            .I(N__19151));
    InMux I__3446 (
            .O(N__19196),
            .I(N__19151));
    InMux I__3445 (
            .O(N__19195),
            .I(N__19146));
    InMux I__3444 (
            .O(N__19194),
            .I(N__19146));
    LocalMux I__3443 (
            .O(N__19191),
            .I(N__19143));
    InMux I__3442 (
            .O(N__19190),
            .I(N__19140));
    InMux I__3441 (
            .O(N__19189),
            .I(N__19133));
    InMux I__3440 (
            .O(N__19188),
            .I(N__19133));
    InMux I__3439 (
            .O(N__19185),
            .I(N__19133));
    LocalMux I__3438 (
            .O(N__19180),
            .I(N__19126));
    Span4Mux_v I__3437 (
            .O(N__19177),
            .I(N__19126));
    LocalMux I__3436 (
            .O(N__19174),
            .I(N__19126));
    InMux I__3435 (
            .O(N__19173),
            .I(N__19115));
    InMux I__3434 (
            .O(N__19172),
            .I(N__19115));
    InMux I__3433 (
            .O(N__19169),
            .I(N__19115));
    InMux I__3432 (
            .O(N__19168),
            .I(N__19115));
    InMux I__3431 (
            .O(N__19165),
            .I(N__19115));
    InMux I__3430 (
            .O(N__19162),
            .I(N__19108));
    InMux I__3429 (
            .O(N__19161),
            .I(N__19108));
    InMux I__3428 (
            .O(N__19158),
            .I(N__19108));
    LocalMux I__3427 (
            .O(N__19151),
            .I(N__19101));
    LocalMux I__3426 (
            .O(N__19146),
            .I(N__19101));
    Span4Mux_h I__3425 (
            .O(N__19143),
            .I(N__19101));
    LocalMux I__3424 (
            .O(N__19140),
            .I(\eeprom.n3430 ));
    LocalMux I__3423 (
            .O(N__19133),
            .I(\eeprom.n3430 ));
    Odrv4 I__3422 (
            .O(N__19126),
            .I(\eeprom.n3430 ));
    LocalMux I__3421 (
            .O(N__19115),
            .I(\eeprom.n3430 ));
    LocalMux I__3420 (
            .O(N__19108),
            .I(\eeprom.n3430 ));
    Odrv4 I__3419 (
            .O(N__19101),
            .I(\eeprom.n3430 ));
    CascadeMux I__3418 (
            .O(N__19088),
            .I(N__19085));
    InMux I__3417 (
            .O(N__19085),
            .I(N__19081));
    InMux I__3416 (
            .O(N__19084),
            .I(N__19078));
    LocalMux I__3415 (
            .O(N__19081),
            .I(N__19075));
    LocalMux I__3414 (
            .O(N__19078),
            .I(N__19071));
    Span4Mux_h I__3413 (
            .O(N__19075),
            .I(N__19068));
    InMux I__3412 (
            .O(N__19074),
            .I(N__19065));
    Span4Mux_h I__3411 (
            .O(N__19071),
            .I(N__19062));
    Odrv4 I__3410 (
            .O(N__19068),
            .I(\eeprom.n3502 ));
    LocalMux I__3409 (
            .O(N__19065),
            .I(\eeprom.n3502 ));
    Odrv4 I__3408 (
            .O(N__19062),
            .I(\eeprom.n3502 ));
    CascadeMux I__3407 (
            .O(N__19055),
            .I(\eeprom.n2511_cascade_ ));
    CascadeMux I__3406 (
            .O(N__19052),
            .I(\eeprom.n2618_cascade_ ));
    InMux I__3405 (
            .O(N__19049),
            .I(bfn_21_23_0_));
    InMux I__3404 (
            .O(N__19046),
            .I(N__19043));
    LocalMux I__3403 (
            .O(N__19043),
            .I(\eeprom.n2685 ));
    InMux I__3402 (
            .O(N__19040),
            .I(\eeprom.n4043 ));
    InMux I__3401 (
            .O(N__19037),
            .I(\eeprom.n4044 ));
    InMux I__3400 (
            .O(N__19034),
            .I(\eeprom.n4045 ));
    InMux I__3399 (
            .O(N__19031),
            .I(\eeprom.n4009 ));
    InMux I__3398 (
            .O(N__19028),
            .I(\eeprom.n4010 ));
    InMux I__3397 (
            .O(N__19025),
            .I(\eeprom.n4011 ));
    InMux I__3396 (
            .O(N__19022),
            .I(\eeprom.n4012 ));
    InMux I__3395 (
            .O(N__19019),
            .I(\eeprom.n4013 ));
    InMux I__3394 (
            .O(N__19016),
            .I(bfn_21_21_0_));
    InMux I__3393 (
            .O(N__19013),
            .I(\eeprom.n4015 ));
    InMux I__3392 (
            .O(N__19010),
            .I(\eeprom.n4016 ));
    InMux I__3391 (
            .O(N__19007),
            .I(\eeprom.n4017 ));
    CascadeMux I__3390 (
            .O(N__19004),
            .I(\eeprom.n2214_cascade_ ));
    InMux I__3389 (
            .O(N__19001),
            .I(N__18998));
    LocalMux I__3388 (
            .O(N__18998),
            .I(N__18995));
    Odrv4 I__3387 (
            .O(N__18995),
            .I(\eeprom.n3720 ));
    InMux I__3386 (
            .O(N__18992),
            .I(bfn_21_20_0_));
    InMux I__3385 (
            .O(N__18989),
            .I(\eeprom.n4007 ));
    InMux I__3384 (
            .O(N__18986),
            .I(\eeprom.n4008 ));
    CascadeMux I__3383 (
            .O(N__18983),
            .I(\eeprom.n4847_cascade_ ));
    InMux I__3382 (
            .O(N__18980),
            .I(N__18977));
    LocalMux I__3381 (
            .O(N__18977),
            .I(\eeprom.enable_N_60_5 ));
    InMux I__3380 (
            .O(N__18974),
            .I(N__18971));
    LocalMux I__3379 (
            .O(N__18971),
            .I(\eeprom.enable_N_60_7 ));
    InMux I__3378 (
            .O(N__18968),
            .I(N__18965));
    LocalMux I__3377 (
            .O(N__18965),
            .I(\eeprom.enable_N_60_6 ));
    CascadeMux I__3376 (
            .O(N__18962),
            .I(\eeprom.n4853_cascade_ ));
    InMux I__3375 (
            .O(N__18959),
            .I(N__18956));
    LocalMux I__3374 (
            .O(N__18956),
            .I(\eeprom.enable_N_60_8 ));
    InMux I__3373 (
            .O(N__18953),
            .I(N__18950));
    LocalMux I__3372 (
            .O(N__18950),
            .I(\eeprom.enable_N_60_10 ));
    InMux I__3371 (
            .O(N__18947),
            .I(N__18944));
    LocalMux I__3370 (
            .O(N__18944),
            .I(\eeprom.enable_N_60_9 ));
    CascadeMux I__3369 (
            .O(N__18941),
            .I(\eeprom.n4859_cascade_ ));
    InMux I__3368 (
            .O(N__18938),
            .I(N__18935));
    LocalMux I__3367 (
            .O(N__18935),
            .I(\eeprom.enable_N_60_11 ));
    CascadeMux I__3366 (
            .O(N__18932),
            .I(\eeprom.n4865_cascade_ ));
    CascadeMux I__3365 (
            .O(N__18929),
            .I(\eeprom.enable_N_59_cascade_ ));
    InMux I__3364 (
            .O(N__18926),
            .I(N__18920));
    InMux I__3363 (
            .O(N__18925),
            .I(N__18920));
    LocalMux I__3362 (
            .O(N__18920),
            .I(\eeprom.enable_N_60_12 ));
    InMux I__3361 (
            .O(N__18917),
            .I(N__18911));
    InMux I__3360 (
            .O(N__18916),
            .I(N__18911));
    LocalMux I__3359 (
            .O(N__18911),
            .I(\eeprom.enable_N_60_14 ));
    CascadeMux I__3358 (
            .O(N__18908),
            .I(N__18905));
    InMux I__3357 (
            .O(N__18905),
            .I(N__18901));
    InMux I__3356 (
            .O(N__18904),
            .I(N__18898));
    LocalMux I__3355 (
            .O(N__18901),
            .I(\eeprom.enable_N_60_13 ));
    LocalMux I__3354 (
            .O(N__18898),
            .I(\eeprom.enable_N_60_13 ));
    InMux I__3353 (
            .O(N__18893),
            .I(N__18890));
    LocalMux I__3352 (
            .O(N__18890),
            .I(\eeprom.n4865 ));
    CascadeMux I__3351 (
            .O(N__18887),
            .I(\eeprom.n2211_cascade_ ));
    InMux I__3350 (
            .O(N__18884),
            .I(N__18881));
    LocalMux I__3349 (
            .O(N__18881),
            .I(N__18878));
    Odrv4 I__3348 (
            .O(N__18878),
            .I(\eeprom.n2975 ));
    InMux I__3347 (
            .O(N__18875),
            .I(\eeprom.n4098 ));
    InMux I__3346 (
            .O(N__18872),
            .I(N__18869));
    LocalMux I__3345 (
            .O(N__18869),
            .I(N__18866));
    Odrv4 I__3344 (
            .O(N__18866),
            .I(\eeprom.n2974 ));
    InMux I__3343 (
            .O(N__18863),
            .I(\eeprom.n4099 ));
    CascadeMux I__3342 (
            .O(N__18860),
            .I(N__18857));
    InMux I__3341 (
            .O(N__18857),
            .I(N__18853));
    InMux I__3340 (
            .O(N__18856),
            .I(N__18850));
    LocalMux I__3339 (
            .O(N__18853),
            .I(N__18844));
    LocalMux I__3338 (
            .O(N__18850),
            .I(N__18844));
    InMux I__3337 (
            .O(N__18849),
            .I(N__18841));
    Odrv4 I__3336 (
            .O(N__18844),
            .I(\eeprom.n2906 ));
    LocalMux I__3335 (
            .O(N__18841),
            .I(\eeprom.n2906 ));
    InMux I__3334 (
            .O(N__18836),
            .I(N__18833));
    LocalMux I__3333 (
            .O(N__18833),
            .I(N__18830));
    Odrv4 I__3332 (
            .O(N__18830),
            .I(\eeprom.n2973 ));
    InMux I__3331 (
            .O(N__18827),
            .I(\eeprom.n4100 ));
    CascadeMux I__3330 (
            .O(N__18824),
            .I(N__18821));
    InMux I__3329 (
            .O(N__18821),
            .I(N__18818));
    LocalMux I__3328 (
            .O(N__18818),
            .I(N__18815));
    Odrv4 I__3327 (
            .O(N__18815),
            .I(\eeprom.n2972 ));
    InMux I__3326 (
            .O(N__18812),
            .I(\eeprom.n4101 ));
    InMux I__3325 (
            .O(N__18809),
            .I(N__18806));
    LocalMux I__3324 (
            .O(N__18806),
            .I(\eeprom.n2971 ));
    InMux I__3323 (
            .O(N__18803),
            .I(\eeprom.n4102 ));
    InMux I__3322 (
            .O(N__18800),
            .I(N__18797));
    LocalMux I__3321 (
            .O(N__18797),
            .I(N__18794));
    Span4Mux_v I__3320 (
            .O(N__18794),
            .I(N__18791));
    Odrv4 I__3319 (
            .O(N__18791),
            .I(\eeprom.n2970 ));
    InMux I__3318 (
            .O(N__18788),
            .I(bfn_20_31_0_));
    CascadeMux I__3317 (
            .O(N__18785),
            .I(N__18780));
    CascadeMux I__3316 (
            .O(N__18784),
            .I(N__18771));
    CascadeMux I__3315 (
            .O(N__18783),
            .I(N__18767));
    InMux I__3314 (
            .O(N__18780),
            .I(N__18764));
    InMux I__3313 (
            .O(N__18779),
            .I(N__18761));
    CascadeMux I__3312 (
            .O(N__18778),
            .I(N__18757));
    CascadeMux I__3311 (
            .O(N__18777),
            .I(N__18754));
    CascadeMux I__3310 (
            .O(N__18776),
            .I(N__18750));
    CascadeMux I__3309 (
            .O(N__18775),
            .I(N__18747));
    CascadeMux I__3308 (
            .O(N__18774),
            .I(N__18742));
    InMux I__3307 (
            .O(N__18771),
            .I(N__18733));
    InMux I__3306 (
            .O(N__18770),
            .I(N__18733));
    InMux I__3305 (
            .O(N__18767),
            .I(N__18733));
    LocalMux I__3304 (
            .O(N__18764),
            .I(N__18730));
    LocalMux I__3303 (
            .O(N__18761),
            .I(N__18727));
    CascadeMux I__3302 (
            .O(N__18760),
            .I(N__18724));
    InMux I__3301 (
            .O(N__18757),
            .I(N__18714));
    InMux I__3300 (
            .O(N__18754),
            .I(N__18714));
    InMux I__3299 (
            .O(N__18753),
            .I(N__18714));
    InMux I__3298 (
            .O(N__18750),
            .I(N__18714));
    InMux I__3297 (
            .O(N__18747),
            .I(N__18707));
    InMux I__3296 (
            .O(N__18746),
            .I(N__18707));
    InMux I__3295 (
            .O(N__18745),
            .I(N__18707));
    InMux I__3294 (
            .O(N__18742),
            .I(N__18700));
    InMux I__3293 (
            .O(N__18741),
            .I(N__18700));
    InMux I__3292 (
            .O(N__18740),
            .I(N__18700));
    LocalMux I__3291 (
            .O(N__18733),
            .I(N__18693));
    Span4Mux_s2_v I__3290 (
            .O(N__18730),
            .I(N__18693));
    Span4Mux_h I__3289 (
            .O(N__18727),
            .I(N__18693));
    InMux I__3288 (
            .O(N__18724),
            .I(N__18688));
    InMux I__3287 (
            .O(N__18723),
            .I(N__18688));
    LocalMux I__3286 (
            .O(N__18714),
            .I(\eeprom.n2935 ));
    LocalMux I__3285 (
            .O(N__18707),
            .I(\eeprom.n2935 ));
    LocalMux I__3284 (
            .O(N__18700),
            .I(\eeprom.n2935 ));
    Odrv4 I__3283 (
            .O(N__18693),
            .I(\eeprom.n2935 ));
    LocalMux I__3282 (
            .O(N__18688),
            .I(\eeprom.n2935 ));
    InMux I__3281 (
            .O(N__18677),
            .I(\eeprom.n4104 ));
    InMux I__3280 (
            .O(N__18674),
            .I(N__18670));
    InMux I__3279 (
            .O(N__18673),
            .I(N__18667));
    LocalMux I__3278 (
            .O(N__18670),
            .I(N__18664));
    LocalMux I__3277 (
            .O(N__18667),
            .I(N__18661));
    Span4Mux_v I__3276 (
            .O(N__18664),
            .I(N__18658));
    Odrv4 I__3275 (
            .O(N__18661),
            .I(\eeprom.n3001 ));
    Odrv4 I__3274 (
            .O(N__18658),
            .I(\eeprom.n3001 ));
    InMux I__3273 (
            .O(N__18653),
            .I(N__18650));
    LocalMux I__3272 (
            .O(N__18650),
            .I(\eeprom.enable_N_60_0 ));
    InMux I__3271 (
            .O(N__18647),
            .I(N__18644));
    LocalMux I__3270 (
            .O(N__18644),
            .I(\eeprom.enable_N_60_1 ));
    InMux I__3269 (
            .O(N__18641),
            .I(N__18638));
    LocalMux I__3268 (
            .O(N__18638),
            .I(\eeprom.enable_N_60_2 ));
    InMux I__3267 (
            .O(N__18635),
            .I(N__18632));
    LocalMux I__3266 (
            .O(N__18632),
            .I(N__18629));
    Odrv4 I__3265 (
            .O(N__18629),
            .I(\eeprom.enable_N_60_3 ));
    InMux I__3264 (
            .O(N__18626),
            .I(N__18623));
    LocalMux I__3263 (
            .O(N__18623),
            .I(\eeprom.enable_N_60_4 ));
    InMux I__3262 (
            .O(N__18620),
            .I(\eeprom.n4090 ));
    CascadeMux I__3261 (
            .O(N__18617),
            .I(N__18613));
    CascadeMux I__3260 (
            .O(N__18616),
            .I(N__18610));
    InMux I__3259 (
            .O(N__18613),
            .I(N__18606));
    InMux I__3258 (
            .O(N__18610),
            .I(N__18603));
    InMux I__3257 (
            .O(N__18609),
            .I(N__18600));
    LocalMux I__3256 (
            .O(N__18606),
            .I(\eeprom.n2915 ));
    LocalMux I__3255 (
            .O(N__18603),
            .I(\eeprom.n2915 ));
    LocalMux I__3254 (
            .O(N__18600),
            .I(\eeprom.n2915 ));
    InMux I__3253 (
            .O(N__18593),
            .I(N__18590));
    LocalMux I__3252 (
            .O(N__18590),
            .I(N__18587));
    Span4Mux_h I__3251 (
            .O(N__18587),
            .I(N__18584));
    Odrv4 I__3250 (
            .O(N__18584),
            .I(\eeprom.n2982 ));
    InMux I__3249 (
            .O(N__18581),
            .I(\eeprom.n4091 ));
    CascadeMux I__3248 (
            .O(N__18578),
            .I(N__18575));
    InMux I__3247 (
            .O(N__18575),
            .I(N__18571));
    InMux I__3246 (
            .O(N__18574),
            .I(N__18568));
    LocalMux I__3245 (
            .O(N__18571),
            .I(N__18565));
    LocalMux I__3244 (
            .O(N__18568),
            .I(\eeprom.n2914 ));
    Odrv4 I__3243 (
            .O(N__18565),
            .I(\eeprom.n2914 ));
    CascadeMux I__3242 (
            .O(N__18560),
            .I(N__18557));
    InMux I__3241 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__3240 (
            .O(N__18554),
            .I(N__18551));
    Odrv4 I__3239 (
            .O(N__18551),
            .I(\eeprom.n2981 ));
    InMux I__3238 (
            .O(N__18548),
            .I(\eeprom.n4092 ));
    InMux I__3237 (
            .O(N__18545),
            .I(N__18541));
    InMux I__3236 (
            .O(N__18544),
            .I(N__18538));
    LocalMux I__3235 (
            .O(N__18541),
            .I(\eeprom.n2913 ));
    LocalMux I__3234 (
            .O(N__18538),
            .I(\eeprom.n2913 ));
    CascadeMux I__3233 (
            .O(N__18533),
            .I(N__18530));
    InMux I__3232 (
            .O(N__18530),
            .I(N__18527));
    LocalMux I__3231 (
            .O(N__18527),
            .I(N__18524));
    Odrv4 I__3230 (
            .O(N__18524),
            .I(\eeprom.n2980 ));
    InMux I__3229 (
            .O(N__18521),
            .I(\eeprom.n4093 ));
    InMux I__3228 (
            .O(N__18518),
            .I(N__18515));
    LocalMux I__3227 (
            .O(N__18515),
            .I(N__18512));
    Span4Mux_v I__3226 (
            .O(N__18512),
            .I(N__18509));
    Odrv4 I__3225 (
            .O(N__18509),
            .I(\eeprom.n2979 ));
    InMux I__3224 (
            .O(N__18506),
            .I(\eeprom.n4094 ));
    InMux I__3223 (
            .O(N__18503),
            .I(N__18500));
    LocalMux I__3222 (
            .O(N__18500),
            .I(\eeprom.n2978 ));
    InMux I__3221 (
            .O(N__18497),
            .I(bfn_20_30_0_));
    CascadeMux I__3220 (
            .O(N__18494),
            .I(N__18490));
    InMux I__3219 (
            .O(N__18493),
            .I(N__18487));
    InMux I__3218 (
            .O(N__18490),
            .I(N__18484));
    LocalMux I__3217 (
            .O(N__18487),
            .I(N__18481));
    LocalMux I__3216 (
            .O(N__18484),
            .I(\eeprom.n2910 ));
    Odrv12 I__3215 (
            .O(N__18481),
            .I(\eeprom.n2910 ));
    InMux I__3214 (
            .O(N__18476),
            .I(N__18473));
    LocalMux I__3213 (
            .O(N__18473),
            .I(N__18470));
    Span4Mux_v I__3212 (
            .O(N__18470),
            .I(N__18467));
    Odrv4 I__3211 (
            .O(N__18467),
            .I(\eeprom.n2977 ));
    InMux I__3210 (
            .O(N__18464),
            .I(\eeprom.n4096 ));
    InMux I__3209 (
            .O(N__18461),
            .I(N__18456));
    InMux I__3208 (
            .O(N__18460),
            .I(N__18453));
    InMux I__3207 (
            .O(N__18459),
            .I(N__18450));
    LocalMux I__3206 (
            .O(N__18456),
            .I(N__18445));
    LocalMux I__3205 (
            .O(N__18453),
            .I(N__18445));
    LocalMux I__3204 (
            .O(N__18450),
            .I(\eeprom.n2909 ));
    Odrv4 I__3203 (
            .O(N__18445),
            .I(\eeprom.n2909 ));
    InMux I__3202 (
            .O(N__18440),
            .I(N__18437));
    LocalMux I__3201 (
            .O(N__18437),
            .I(N__18434));
    Odrv4 I__3200 (
            .O(N__18434),
            .I(\eeprom.n2976 ));
    InMux I__3199 (
            .O(N__18431),
            .I(\eeprom.n4097 ));
    InMux I__3198 (
            .O(N__18428),
            .I(N__18423));
    InMux I__3197 (
            .O(N__18427),
            .I(N__18420));
    InMux I__3196 (
            .O(N__18426),
            .I(N__18417));
    LocalMux I__3195 (
            .O(N__18423),
            .I(N__18414));
    LocalMux I__3194 (
            .O(N__18420),
            .I(\eeprom.n2908 ));
    LocalMux I__3193 (
            .O(N__18417),
            .I(\eeprom.n2908 ));
    Odrv4 I__3192 (
            .O(N__18414),
            .I(\eeprom.n2908 ));
    CascadeMux I__3191 (
            .O(N__18407),
            .I(\eeprom.n2836_cascade_ ));
    CascadeMux I__3190 (
            .O(N__18404),
            .I(\eeprom.n2913_cascade_ ));
    InMux I__3189 (
            .O(N__18401),
            .I(N__18398));
    LocalMux I__3188 (
            .O(N__18398),
            .I(\eeprom.n5297 ));
    InMux I__3187 (
            .O(N__18395),
            .I(N__18392));
    LocalMux I__3186 (
            .O(N__18392),
            .I(N__18389));
    Span4Mux_h I__3185 (
            .O(N__18389),
            .I(N__18386));
    Odrv4 I__3184 (
            .O(N__18386),
            .I(\eeprom.n2986 ));
    InMux I__3183 (
            .O(N__18383),
            .I(bfn_20_29_0_));
    InMux I__3182 (
            .O(N__18380),
            .I(N__18377));
    LocalMux I__3181 (
            .O(N__18377),
            .I(N__18374));
    Odrv4 I__3180 (
            .O(N__18374),
            .I(\eeprom.n2985 ));
    InMux I__3179 (
            .O(N__18371),
            .I(\eeprom.n4088 ));
    CascadeMux I__3178 (
            .O(N__18368),
            .I(N__18365));
    InMux I__3177 (
            .O(N__18365),
            .I(N__18360));
    InMux I__3176 (
            .O(N__18364),
            .I(N__18355));
    InMux I__3175 (
            .O(N__18363),
            .I(N__18355));
    LocalMux I__3174 (
            .O(N__18360),
            .I(\eeprom.n2917 ));
    LocalMux I__3173 (
            .O(N__18355),
            .I(\eeprom.n2917 ));
    CascadeMux I__3172 (
            .O(N__18350),
            .I(N__18347));
    InMux I__3171 (
            .O(N__18347),
            .I(N__18344));
    LocalMux I__3170 (
            .O(N__18344),
            .I(N__18341));
    Odrv4 I__3169 (
            .O(N__18341),
            .I(\eeprom.n2984 ));
    InMux I__3168 (
            .O(N__18338),
            .I(\eeprom.n4089 ));
    CascadeMux I__3167 (
            .O(N__18335),
            .I(N__18332));
    InMux I__3166 (
            .O(N__18332),
            .I(N__18328));
    InMux I__3165 (
            .O(N__18331),
            .I(N__18324));
    LocalMux I__3164 (
            .O(N__18328),
            .I(N__18321));
    InMux I__3163 (
            .O(N__18327),
            .I(N__18318));
    LocalMux I__3162 (
            .O(N__18324),
            .I(\eeprom.n2916 ));
    Odrv4 I__3161 (
            .O(N__18321),
            .I(\eeprom.n2916 ));
    LocalMux I__3160 (
            .O(N__18318),
            .I(\eeprom.n2916 ));
    InMux I__3159 (
            .O(N__18311),
            .I(N__18308));
    LocalMux I__3158 (
            .O(N__18308),
            .I(N__18305));
    Odrv4 I__3157 (
            .O(N__18305),
            .I(\eeprom.n2983 ));
    CascadeMux I__3156 (
            .O(N__18302),
            .I(\eeprom.n2910_cascade_ ));
    InMux I__3155 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__3154 (
            .O(N__18296),
            .I(\eeprom.n15_adj_300 ));
    CascadeMux I__3153 (
            .O(N__18293),
            .I(\eeprom.n22_adj_331_cascade_ ));
    InMux I__3152 (
            .O(N__18290),
            .I(N__18287));
    LocalMux I__3151 (
            .O(N__18287),
            .I(\eeprom.n18_adj_330 ));
    CascadeMux I__3150 (
            .O(N__18284),
            .I(\eeprom.n2935_cascade_ ));
    CascadeMux I__3149 (
            .O(N__18281),
            .I(N__18278));
    InMux I__3148 (
            .O(N__18278),
            .I(N__18274));
    InMux I__3147 (
            .O(N__18277),
            .I(N__18271));
    LocalMux I__3146 (
            .O(N__18274),
            .I(N__18268));
    LocalMux I__3145 (
            .O(N__18271),
            .I(N__18263));
    Span4Mux_h I__3144 (
            .O(N__18268),
            .I(N__18263));
    Odrv4 I__3143 (
            .O(N__18263),
            .I(\eeprom.n3015 ));
    CascadeMux I__3142 (
            .O(N__18260),
            .I(N__18257));
    InMux I__3141 (
            .O(N__18257),
            .I(N__18254));
    LocalMux I__3140 (
            .O(N__18254),
            .I(N__18251));
    Span4Mux_v I__3139 (
            .O(N__18251),
            .I(N__18247));
    InMux I__3138 (
            .O(N__18250),
            .I(N__18244));
    Odrv4 I__3137 (
            .O(N__18247),
            .I(\eeprom.n3013 ));
    LocalMux I__3136 (
            .O(N__18244),
            .I(\eeprom.n3013 ));
    CascadeMux I__3135 (
            .O(N__18239),
            .I(\eeprom.n3015_cascade_ ));
    InMux I__3134 (
            .O(N__18236),
            .I(N__18233));
    LocalMux I__3133 (
            .O(N__18233),
            .I(\eeprom.n5143 ));
    CascadeMux I__3132 (
            .O(N__18230),
            .I(\eeprom.n18_adj_290_cascade_ ));
    CascadeMux I__3131 (
            .O(N__18227),
            .I(\eeprom.n20_adj_291_cascade_ ));
    InMux I__3130 (
            .O(N__18224),
            .I(N__18220));
    InMux I__3129 (
            .O(N__18223),
            .I(N__18217));
    LocalMux I__3128 (
            .O(N__18220),
            .I(N__18213));
    LocalMux I__3127 (
            .O(N__18217),
            .I(N__18210));
    InMux I__3126 (
            .O(N__18216),
            .I(N__18207));
    Span4Mux_h I__3125 (
            .O(N__18213),
            .I(N__18204));
    Odrv4 I__3124 (
            .O(N__18210),
            .I(\eeprom.n3211 ));
    LocalMux I__3123 (
            .O(N__18207),
            .I(\eeprom.n3211 ));
    Odrv4 I__3122 (
            .O(N__18204),
            .I(\eeprom.n3211 ));
    CascadeMux I__3121 (
            .O(N__18197),
            .I(\eeprom.n3208_cascade_ ));
    CascadeMux I__3120 (
            .O(N__18194),
            .I(N__18190));
    InMux I__3119 (
            .O(N__18193),
            .I(N__18187));
    InMux I__3118 (
            .O(N__18190),
            .I(N__18183));
    LocalMux I__3117 (
            .O(N__18187),
            .I(N__18180));
    InMux I__3116 (
            .O(N__18186),
            .I(N__18177));
    LocalMux I__3115 (
            .O(N__18183),
            .I(N__18172));
    Span4Mux_h I__3114 (
            .O(N__18180),
            .I(N__18172));
    LocalMux I__3113 (
            .O(N__18177),
            .I(\eeprom.n3210 ));
    Odrv4 I__3112 (
            .O(N__18172),
            .I(\eeprom.n3210 ));
    InMux I__3111 (
            .O(N__18167),
            .I(N__18164));
    LocalMux I__3110 (
            .O(N__18164),
            .I(\eeprom.n26_adj_302 ));
    InMux I__3109 (
            .O(N__18161),
            .I(N__18158));
    LocalMux I__3108 (
            .O(N__18158),
            .I(N__18155));
    Span4Mux_h I__3107 (
            .O(N__18155),
            .I(N__18152));
    Odrv4 I__3106 (
            .O(N__18152),
            .I(\eeprom.n3080 ));
    CascadeMux I__3105 (
            .O(N__18149),
            .I(\eeprom.n3013_cascade_ ));
    InMux I__3104 (
            .O(N__18146),
            .I(N__18139));
    CascadeMux I__3103 (
            .O(N__18145),
            .I(N__18135));
    InMux I__3102 (
            .O(N__18144),
            .I(N__18130));
    CascadeMux I__3101 (
            .O(N__18143),
            .I(N__18125));
    CascadeMux I__3100 (
            .O(N__18142),
            .I(N__18121));
    LocalMux I__3099 (
            .O(N__18139),
            .I(N__18116));
    InMux I__3098 (
            .O(N__18138),
            .I(N__18111));
    InMux I__3097 (
            .O(N__18135),
            .I(N__18111));
    CascadeMux I__3096 (
            .O(N__18134),
            .I(N__18105));
    CascadeMux I__3095 (
            .O(N__18133),
            .I(N__18102));
    LocalMux I__3094 (
            .O(N__18130),
            .I(N__18097));
    InMux I__3093 (
            .O(N__18129),
            .I(N__18092));
    InMux I__3092 (
            .O(N__18128),
            .I(N__18092));
    InMux I__3091 (
            .O(N__18125),
            .I(N__18089));
    InMux I__3090 (
            .O(N__18124),
            .I(N__18080));
    InMux I__3089 (
            .O(N__18121),
            .I(N__18080));
    InMux I__3088 (
            .O(N__18120),
            .I(N__18080));
    InMux I__3087 (
            .O(N__18119),
            .I(N__18080));
    Span4Mux_v I__3086 (
            .O(N__18116),
            .I(N__18075));
    LocalMux I__3085 (
            .O(N__18111),
            .I(N__18075));
    InMux I__3084 (
            .O(N__18110),
            .I(N__18068));
    InMux I__3083 (
            .O(N__18109),
            .I(N__18068));
    InMux I__3082 (
            .O(N__18108),
            .I(N__18068));
    InMux I__3081 (
            .O(N__18105),
            .I(N__18059));
    InMux I__3080 (
            .O(N__18102),
            .I(N__18059));
    InMux I__3079 (
            .O(N__18101),
            .I(N__18059));
    InMux I__3078 (
            .O(N__18100),
            .I(N__18059));
    Span4Mux_h I__3077 (
            .O(N__18097),
            .I(N__18056));
    LocalMux I__3076 (
            .O(N__18092),
            .I(\eeprom.n3034 ));
    LocalMux I__3075 (
            .O(N__18089),
            .I(\eeprom.n3034 ));
    LocalMux I__3074 (
            .O(N__18080),
            .I(\eeprom.n3034 ));
    Odrv4 I__3073 (
            .O(N__18075),
            .I(\eeprom.n3034 ));
    LocalMux I__3072 (
            .O(N__18068),
            .I(\eeprom.n3034 ));
    LocalMux I__3071 (
            .O(N__18059),
            .I(\eeprom.n3034 ));
    Odrv4 I__3070 (
            .O(N__18056),
            .I(\eeprom.n3034 ));
    CascadeMux I__3069 (
            .O(N__18041),
            .I(N__18038));
    InMux I__3068 (
            .O(N__18038),
            .I(N__18035));
    LocalMux I__3067 (
            .O(N__18035),
            .I(N__18030));
    InMux I__3066 (
            .O(N__18034),
            .I(N__18025));
    InMux I__3065 (
            .O(N__18033),
            .I(N__18025));
    Span4Mux_v I__3064 (
            .O(N__18030),
            .I(N__18022));
    LocalMux I__3063 (
            .O(N__18025),
            .I(\eeprom.n3112 ));
    Odrv4 I__3062 (
            .O(N__18022),
            .I(\eeprom.n3112 ));
    CascadeMux I__3061 (
            .O(N__18017),
            .I(N__18014));
    InMux I__3060 (
            .O(N__18014),
            .I(N__18010));
    InMux I__3059 (
            .O(N__18013),
            .I(N__18006));
    LocalMux I__3058 (
            .O(N__18010),
            .I(N__18003));
    InMux I__3057 (
            .O(N__18009),
            .I(N__18000));
    LocalMux I__3056 (
            .O(N__18006),
            .I(N__17995));
    Span4Mux_v I__3055 (
            .O(N__18003),
            .I(N__17995));
    LocalMux I__3054 (
            .O(N__18000),
            .I(\eeprom.n3011 ));
    Odrv4 I__3053 (
            .O(N__17995),
            .I(\eeprom.n3011 ));
    InMux I__3052 (
            .O(N__17990),
            .I(N__17987));
    LocalMux I__3051 (
            .O(N__17987),
            .I(\eeprom.n5301 ));
    InMux I__3050 (
            .O(N__17984),
            .I(N__17980));
    InMux I__3049 (
            .O(N__17983),
            .I(N__17976));
    LocalMux I__3048 (
            .O(N__17980),
            .I(N__17973));
    InMux I__3047 (
            .O(N__17979),
            .I(N__17970));
    LocalMux I__3046 (
            .O(N__17976),
            .I(N__17967));
    Span4Mux_s3_v I__3045 (
            .O(N__17973),
            .I(N__17964));
    LocalMux I__3044 (
            .O(N__17970),
            .I(\eeprom.n3110 ));
    Odrv4 I__3043 (
            .O(N__17967),
            .I(\eeprom.n3110 ));
    Odrv4 I__3042 (
            .O(N__17964),
            .I(\eeprom.n3110 ));
    CascadeMux I__3041 (
            .O(N__17957),
            .I(N__17949));
    CascadeMux I__3040 (
            .O(N__17956),
            .I(N__17942));
    CascadeMux I__3039 (
            .O(N__17955),
            .I(N__17938));
    InMux I__3038 (
            .O(N__17954),
            .I(N__17935));
    CascadeMux I__3037 (
            .O(N__17953),
            .I(N__17930));
    CascadeMux I__3036 (
            .O(N__17952),
            .I(N__17927));
    InMux I__3035 (
            .O(N__17949),
            .I(N__17923));
    CascadeMux I__3034 (
            .O(N__17948),
            .I(N__17916));
    InMux I__3033 (
            .O(N__17947),
            .I(N__17912));
    InMux I__3032 (
            .O(N__17946),
            .I(N__17907));
    InMux I__3031 (
            .O(N__17945),
            .I(N__17907));
    InMux I__3030 (
            .O(N__17942),
            .I(N__17902));
    InMux I__3029 (
            .O(N__17941),
            .I(N__17902));
    InMux I__3028 (
            .O(N__17938),
            .I(N__17899));
    LocalMux I__3027 (
            .O(N__17935),
            .I(N__17896));
    InMux I__3026 (
            .O(N__17934),
            .I(N__17885));
    InMux I__3025 (
            .O(N__17933),
            .I(N__17885));
    InMux I__3024 (
            .O(N__17930),
            .I(N__17885));
    InMux I__3023 (
            .O(N__17927),
            .I(N__17885));
    InMux I__3022 (
            .O(N__17926),
            .I(N__17885));
    LocalMux I__3021 (
            .O(N__17923),
            .I(N__17882));
    InMux I__3020 (
            .O(N__17922),
            .I(N__17879));
    InMux I__3019 (
            .O(N__17921),
            .I(N__17868));
    InMux I__3018 (
            .O(N__17920),
            .I(N__17868));
    InMux I__3017 (
            .O(N__17919),
            .I(N__17868));
    InMux I__3016 (
            .O(N__17916),
            .I(N__17868));
    InMux I__3015 (
            .O(N__17915),
            .I(N__17868));
    LocalMux I__3014 (
            .O(N__17912),
            .I(\eeprom.n3133 ));
    LocalMux I__3013 (
            .O(N__17907),
            .I(\eeprom.n3133 ));
    LocalMux I__3012 (
            .O(N__17902),
            .I(\eeprom.n3133 ));
    LocalMux I__3011 (
            .O(N__17899),
            .I(\eeprom.n3133 ));
    Odrv4 I__3010 (
            .O(N__17896),
            .I(\eeprom.n3133 ));
    LocalMux I__3009 (
            .O(N__17885),
            .I(\eeprom.n3133 ));
    Odrv12 I__3008 (
            .O(N__17882),
            .I(\eeprom.n3133 ));
    LocalMux I__3007 (
            .O(N__17879),
            .I(\eeprom.n3133 ));
    LocalMux I__3006 (
            .O(N__17868),
            .I(\eeprom.n3133 ));
    InMux I__3005 (
            .O(N__17849),
            .I(N__17846));
    LocalMux I__3004 (
            .O(N__17846),
            .I(N__17843));
    Span4Mux_v I__3003 (
            .O(N__17843),
            .I(N__17840));
    Odrv4 I__3002 (
            .O(N__17840),
            .I(\eeprom.n3177 ));
    InMux I__3001 (
            .O(N__17837),
            .I(N__17833));
    CascadeMux I__3000 (
            .O(N__17836),
            .I(N__17830));
    LocalMux I__2999 (
            .O(N__17833),
            .I(N__17827));
    InMux I__2998 (
            .O(N__17830),
            .I(N__17824));
    Span4Mux_h I__2997 (
            .O(N__17827),
            .I(N__17821));
    LocalMux I__2996 (
            .O(N__17824),
            .I(N__17817));
    Span4Mux_h I__2995 (
            .O(N__17821),
            .I(N__17814));
    InMux I__2994 (
            .O(N__17820),
            .I(N__17811));
    Span4Mux_h I__2993 (
            .O(N__17817),
            .I(N__17808));
    Odrv4 I__2992 (
            .O(N__17814),
            .I(\eeprom.n3209 ));
    LocalMux I__2991 (
            .O(N__17811),
            .I(\eeprom.n3209 ));
    Odrv4 I__2990 (
            .O(N__17808),
            .I(\eeprom.n3209 ));
    CascadeMux I__2989 (
            .O(N__17801),
            .I(N__17798));
    InMux I__2988 (
            .O(N__17798),
            .I(N__17795));
    LocalMux I__2987 (
            .O(N__17795),
            .I(N__17792));
    Span4Mux_h I__2986 (
            .O(N__17792),
            .I(N__17789));
    Odrv4 I__2985 (
            .O(N__17789),
            .I(\eeprom.n3283 ));
    CascadeMux I__2984 (
            .O(N__17786),
            .I(N__17783));
    InMux I__2983 (
            .O(N__17783),
            .I(N__17779));
    InMux I__2982 (
            .O(N__17782),
            .I(N__17768));
    LocalMux I__2981 (
            .O(N__17779),
            .I(N__17765));
    CascadeMux I__2980 (
            .O(N__17778),
            .I(N__17759));
    CascadeMux I__2979 (
            .O(N__17777),
            .I(N__17755));
    CascadeMux I__2978 (
            .O(N__17776),
            .I(N__17751));
    CascadeMux I__2977 (
            .O(N__17775),
            .I(N__17748));
    CascadeMux I__2976 (
            .O(N__17774),
            .I(N__17745));
    CascadeMux I__2975 (
            .O(N__17773),
            .I(N__17741));
    InMux I__2974 (
            .O(N__17772),
            .I(N__17737));
    CascadeMux I__2973 (
            .O(N__17771),
            .I(N__17732));
    LocalMux I__2972 (
            .O(N__17768),
            .I(N__17726));
    Span4Mux_v I__2971 (
            .O(N__17765),
            .I(N__17726));
    InMux I__2970 (
            .O(N__17764),
            .I(N__17721));
    InMux I__2969 (
            .O(N__17763),
            .I(N__17721));
    InMux I__2968 (
            .O(N__17762),
            .I(N__17716));
    InMux I__2967 (
            .O(N__17759),
            .I(N__17716));
    InMux I__2966 (
            .O(N__17758),
            .I(N__17709));
    InMux I__2965 (
            .O(N__17755),
            .I(N__17709));
    InMux I__2964 (
            .O(N__17754),
            .I(N__17709));
    InMux I__2963 (
            .O(N__17751),
            .I(N__17700));
    InMux I__2962 (
            .O(N__17748),
            .I(N__17700));
    InMux I__2961 (
            .O(N__17745),
            .I(N__17700));
    InMux I__2960 (
            .O(N__17744),
            .I(N__17700));
    InMux I__2959 (
            .O(N__17741),
            .I(N__17695));
    InMux I__2958 (
            .O(N__17740),
            .I(N__17695));
    LocalMux I__2957 (
            .O(N__17737),
            .I(N__17692));
    InMux I__2956 (
            .O(N__17736),
            .I(N__17689));
    InMux I__2955 (
            .O(N__17735),
            .I(N__17682));
    InMux I__2954 (
            .O(N__17732),
            .I(N__17682));
    InMux I__2953 (
            .O(N__17731),
            .I(N__17682));
    Span4Mux_v I__2952 (
            .O(N__17726),
            .I(N__17679));
    LocalMux I__2951 (
            .O(N__17721),
            .I(\eeprom.n3232 ));
    LocalMux I__2950 (
            .O(N__17716),
            .I(\eeprom.n3232 ));
    LocalMux I__2949 (
            .O(N__17709),
            .I(\eeprom.n3232 ));
    LocalMux I__2948 (
            .O(N__17700),
            .I(\eeprom.n3232 ));
    LocalMux I__2947 (
            .O(N__17695),
            .I(\eeprom.n3232 ));
    Odrv4 I__2946 (
            .O(N__17692),
            .I(\eeprom.n3232 ));
    LocalMux I__2945 (
            .O(N__17689),
            .I(\eeprom.n3232 ));
    LocalMux I__2944 (
            .O(N__17682),
            .I(\eeprom.n3232 ));
    Odrv4 I__2943 (
            .O(N__17679),
            .I(\eeprom.n3232 ));
    CascadeMux I__2942 (
            .O(N__17660),
            .I(N__17656));
    InMux I__2941 (
            .O(N__17659),
            .I(N__17652));
    InMux I__2940 (
            .O(N__17656),
            .I(N__17649));
    CascadeMux I__2939 (
            .O(N__17655),
            .I(N__17646));
    LocalMux I__2938 (
            .O(N__17652),
            .I(N__17643));
    LocalMux I__2937 (
            .O(N__17649),
            .I(N__17640));
    InMux I__2936 (
            .O(N__17646),
            .I(N__17637));
    Odrv4 I__2935 (
            .O(N__17643),
            .I(\eeprom.n3315 ));
    Odrv4 I__2934 (
            .O(N__17640),
            .I(\eeprom.n3315 ));
    LocalMux I__2933 (
            .O(N__17637),
            .I(\eeprom.n3315 ));
    InMux I__2932 (
            .O(N__17630),
            .I(N__17626));
    CascadeMux I__2931 (
            .O(N__17629),
            .I(N__17623));
    LocalMux I__2930 (
            .O(N__17626),
            .I(N__17620));
    InMux I__2929 (
            .O(N__17623),
            .I(N__17617));
    Span4Mux_v I__2928 (
            .O(N__17620),
            .I(N__17613));
    LocalMux I__2927 (
            .O(N__17617),
            .I(N__17610));
    InMux I__2926 (
            .O(N__17616),
            .I(N__17607));
    Odrv4 I__2925 (
            .O(N__17613),
            .I(\eeprom.n3114 ));
    Odrv4 I__2924 (
            .O(N__17610),
            .I(\eeprom.n3114 ));
    LocalMux I__2923 (
            .O(N__17607),
            .I(\eeprom.n3114 ));
    CascadeMux I__2922 (
            .O(N__17600),
            .I(N__17597));
    InMux I__2921 (
            .O(N__17597),
            .I(N__17594));
    LocalMux I__2920 (
            .O(N__17594),
            .I(N__17591));
    Span4Mux_v I__2919 (
            .O(N__17591),
            .I(N__17588));
    Odrv4 I__2918 (
            .O(N__17588),
            .I(\eeprom.n3181 ));
    InMux I__2917 (
            .O(N__17585),
            .I(N__17581));
    InMux I__2916 (
            .O(N__17584),
            .I(N__17578));
    LocalMux I__2915 (
            .O(N__17581),
            .I(N__17575));
    LocalMux I__2914 (
            .O(N__17578),
            .I(N__17572));
    Span4Mux_v I__2913 (
            .O(N__17575),
            .I(N__17569));
    Span4Mux_h I__2912 (
            .O(N__17572),
            .I(N__17566));
    Odrv4 I__2911 (
            .O(N__17569),
            .I(\eeprom.n3213 ));
    Odrv4 I__2910 (
            .O(N__17566),
            .I(\eeprom.n3213 ));
    CascadeMux I__2909 (
            .O(N__17561),
            .I(\eeprom.n3213_cascade_ ));
    InMux I__2908 (
            .O(N__17558),
            .I(N__17555));
    LocalMux I__2907 (
            .O(N__17555),
            .I(N__17552));
    Span4Mux_v I__2906 (
            .O(N__17552),
            .I(N__17549));
    Odrv4 I__2905 (
            .O(N__17549),
            .I(\eeprom.n3182 ));
    CascadeMux I__2904 (
            .O(N__17546),
            .I(N__17543));
    InMux I__2903 (
            .O(N__17543),
            .I(N__17539));
    CascadeMux I__2902 (
            .O(N__17542),
            .I(N__17536));
    LocalMux I__2901 (
            .O(N__17539),
            .I(N__17533));
    InMux I__2900 (
            .O(N__17536),
            .I(N__17530));
    Span4Mux_h I__2899 (
            .O(N__17533),
            .I(N__17526));
    LocalMux I__2898 (
            .O(N__17530),
            .I(N__17523));
    InMux I__2897 (
            .O(N__17529),
            .I(N__17520));
    Odrv4 I__2896 (
            .O(N__17526),
            .I(\eeprom.n3115 ));
    Odrv4 I__2895 (
            .O(N__17523),
            .I(\eeprom.n3115 ));
    LocalMux I__2894 (
            .O(N__17520),
            .I(\eeprom.n3115 ));
    InMux I__2893 (
            .O(N__17513),
            .I(N__17510));
    LocalMux I__2892 (
            .O(N__17510),
            .I(N__17506));
    InMux I__2891 (
            .O(N__17509),
            .I(N__17503));
    Span4Mux_v I__2890 (
            .O(N__17506),
            .I(N__17500));
    LocalMux I__2889 (
            .O(N__17503),
            .I(\eeprom.n3214 ));
    Odrv4 I__2888 (
            .O(N__17500),
            .I(\eeprom.n3214 ));
    CascadeMux I__2887 (
            .O(N__17495),
            .I(N__17492));
    InMux I__2886 (
            .O(N__17492),
            .I(N__17488));
    InMux I__2885 (
            .O(N__17491),
            .I(N__17485));
    LocalMux I__2884 (
            .O(N__17488),
            .I(N__17481));
    LocalMux I__2883 (
            .O(N__17485),
            .I(N__17478));
    InMux I__2882 (
            .O(N__17484),
            .I(N__17475));
    Span4Mux_h I__2881 (
            .O(N__17481),
            .I(N__17472));
    Odrv4 I__2880 (
            .O(N__17478),
            .I(\eeprom.n3216 ));
    LocalMux I__2879 (
            .O(N__17475),
            .I(\eeprom.n3216 ));
    Odrv4 I__2878 (
            .O(N__17472),
            .I(\eeprom.n3216 ));
    CascadeMux I__2877 (
            .O(N__17465),
            .I(\eeprom.n3214_cascade_ ));
    InMux I__2876 (
            .O(N__17462),
            .I(N__17459));
    LocalMux I__2875 (
            .O(N__17459),
            .I(\eeprom.n5205 ));
    CascadeMux I__2874 (
            .O(N__17456),
            .I(N__17453));
    InMux I__2873 (
            .O(N__17453),
            .I(N__17450));
    LocalMux I__2872 (
            .O(N__17450),
            .I(\eeprom.n5209 ));
    InMux I__2871 (
            .O(N__17447),
            .I(N__17443));
    CascadeMux I__2870 (
            .O(N__17446),
            .I(N__17440));
    LocalMux I__2869 (
            .O(N__17443),
            .I(N__17437));
    InMux I__2868 (
            .O(N__17440),
            .I(N__17434));
    Span4Mux_v I__2867 (
            .O(N__17437),
            .I(N__17430));
    LocalMux I__2866 (
            .O(N__17434),
            .I(N__17427));
    InMux I__2865 (
            .O(N__17433),
            .I(N__17424));
    Odrv4 I__2864 (
            .O(N__17430),
            .I(\eeprom.n3116 ));
    Odrv4 I__2863 (
            .O(N__17427),
            .I(\eeprom.n3116 ));
    LocalMux I__2862 (
            .O(N__17424),
            .I(\eeprom.n3116 ));
    CascadeMux I__2861 (
            .O(N__17417),
            .I(N__17414));
    InMux I__2860 (
            .O(N__17414),
            .I(N__17411));
    LocalMux I__2859 (
            .O(N__17411),
            .I(N__17408));
    Span4Mux_v I__2858 (
            .O(N__17408),
            .I(N__17405));
    Odrv4 I__2857 (
            .O(N__17405),
            .I(\eeprom.n3183 ));
    CascadeMux I__2856 (
            .O(N__17402),
            .I(N__17399));
    InMux I__2855 (
            .O(N__17399),
            .I(N__17395));
    InMux I__2854 (
            .O(N__17398),
            .I(N__17392));
    LocalMux I__2853 (
            .O(N__17395),
            .I(N__17389));
    LocalMux I__2852 (
            .O(N__17392),
            .I(N__17385));
    Span4Mux_h I__2851 (
            .O(N__17389),
            .I(N__17382));
    InMux I__2850 (
            .O(N__17388),
            .I(N__17379));
    Odrv4 I__2849 (
            .O(N__17385),
            .I(\eeprom.n3215 ));
    Odrv4 I__2848 (
            .O(N__17382),
            .I(\eeprom.n3215 ));
    LocalMux I__2847 (
            .O(N__17379),
            .I(\eeprom.n3215 ));
    InMux I__2846 (
            .O(N__17372),
            .I(N__17369));
    LocalMux I__2845 (
            .O(N__17369),
            .I(N__17366));
    Span4Mux_v I__2844 (
            .O(N__17366),
            .I(N__17363));
    Odrv4 I__2843 (
            .O(N__17363),
            .I(\eeprom.n3185 ));
    InMux I__2842 (
            .O(N__17360),
            .I(N__17356));
    CascadeMux I__2841 (
            .O(N__17359),
            .I(N__17353));
    LocalMux I__2840 (
            .O(N__17356),
            .I(N__17349));
    InMux I__2839 (
            .O(N__17353),
            .I(N__17346));
    CascadeMux I__2838 (
            .O(N__17352),
            .I(N__17343));
    Span4Mux_v I__2837 (
            .O(N__17349),
            .I(N__17340));
    LocalMux I__2836 (
            .O(N__17346),
            .I(N__17337));
    InMux I__2835 (
            .O(N__17343),
            .I(N__17334));
    Odrv4 I__2834 (
            .O(N__17340),
            .I(\eeprom.n3118 ));
    Odrv12 I__2833 (
            .O(N__17337),
            .I(\eeprom.n3118 ));
    LocalMux I__2832 (
            .O(N__17334),
            .I(\eeprom.n3118 ));
    CascadeMux I__2831 (
            .O(N__17327),
            .I(N__17324));
    InMux I__2830 (
            .O(N__17324),
            .I(N__17321));
    LocalMux I__2829 (
            .O(N__17321),
            .I(N__17316));
    InMux I__2828 (
            .O(N__17320),
            .I(N__17313));
    InMux I__2827 (
            .O(N__17319),
            .I(N__17310));
    Span4Mux_h I__2826 (
            .O(N__17316),
            .I(N__17307));
    LocalMux I__2825 (
            .O(N__17313),
            .I(\eeprom.n3217 ));
    LocalMux I__2824 (
            .O(N__17310),
            .I(\eeprom.n3217 ));
    Odrv4 I__2823 (
            .O(N__17307),
            .I(\eeprom.n3217 ));
    InMux I__2822 (
            .O(N__17300),
            .I(N__17296));
    InMux I__2821 (
            .O(N__17299),
            .I(N__17293));
    LocalMux I__2820 (
            .O(N__17296),
            .I(N__17289));
    LocalMux I__2819 (
            .O(N__17293),
            .I(N__17286));
    InMux I__2818 (
            .O(N__17292),
            .I(N__17283));
    Span4Mux_h I__2817 (
            .O(N__17289),
            .I(N__17280));
    Span4Mux_s2_v I__2816 (
            .O(N__17286),
            .I(N__17277));
    LocalMux I__2815 (
            .O(N__17283),
            .I(N__17274));
    Odrv4 I__2814 (
            .O(N__17280),
            .I(\eeprom.n3109 ));
    Odrv4 I__2813 (
            .O(N__17277),
            .I(\eeprom.n3109 ));
    Odrv4 I__2812 (
            .O(N__17274),
            .I(\eeprom.n3109 ));
    CascadeMux I__2811 (
            .O(N__17267),
            .I(N__17264));
    InMux I__2810 (
            .O(N__17264),
            .I(N__17261));
    LocalMux I__2809 (
            .O(N__17261),
            .I(N__17258));
    Span4Mux_v I__2808 (
            .O(N__17258),
            .I(N__17255));
    Odrv4 I__2807 (
            .O(N__17255),
            .I(\eeprom.n3176 ));
    InMux I__2806 (
            .O(N__17252),
            .I(N__17248));
    InMux I__2805 (
            .O(N__17251),
            .I(N__17245));
    LocalMux I__2804 (
            .O(N__17248),
            .I(N__17242));
    LocalMux I__2803 (
            .O(N__17245),
            .I(N__17239));
    Span4Mux_h I__2802 (
            .O(N__17242),
            .I(N__17234));
    Span4Mux_h I__2801 (
            .O(N__17239),
            .I(N__17234));
    Odrv4 I__2800 (
            .O(N__17234),
            .I(\eeprom.n3208 ));
    CascadeMux I__2799 (
            .O(N__17231),
            .I(\eeprom.n3413_cascade_ ));
    CascadeMux I__2798 (
            .O(N__17228),
            .I(N__17224));
    InMux I__2797 (
            .O(N__17227),
            .I(N__17221));
    InMux I__2796 (
            .O(N__17224),
            .I(N__17218));
    LocalMux I__2795 (
            .O(N__17221),
            .I(N__17212));
    LocalMux I__2794 (
            .O(N__17218),
            .I(N__17212));
    InMux I__2793 (
            .O(N__17217),
            .I(N__17209));
    Span4Mux_h I__2792 (
            .O(N__17212),
            .I(N__17206));
    LocalMux I__2791 (
            .O(N__17209),
            .I(\eeprom.n3415 ));
    Odrv4 I__2790 (
            .O(N__17206),
            .I(\eeprom.n3415 ));
    InMux I__2789 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__2788 (
            .O(N__17198),
            .I(\eeprom.n5289 ));
    InMux I__2787 (
            .O(N__17195),
            .I(N__17192));
    LocalMux I__2786 (
            .O(N__17192),
            .I(N__17189));
    Span4Mux_v I__2785 (
            .O(N__17189),
            .I(N__17186));
    Span4Mux_h I__2784 (
            .O(N__17186),
            .I(N__17183));
    Odrv4 I__2783 (
            .O(N__17183),
            .I(\eeprom.n3278 ));
    CascadeMux I__2782 (
            .O(N__17180),
            .I(N__17177));
    InMux I__2781 (
            .O(N__17177),
            .I(N__17174));
    LocalMux I__2780 (
            .O(N__17174),
            .I(N__17171));
    Span4Mux_h I__2779 (
            .O(N__17171),
            .I(N__17167));
    InMux I__2778 (
            .O(N__17170),
            .I(N__17164));
    Odrv4 I__2777 (
            .O(N__17167),
            .I(\eeprom.n3310 ));
    LocalMux I__2776 (
            .O(N__17164),
            .I(\eeprom.n3310 ));
    InMux I__2775 (
            .O(N__17159),
            .I(N__17152));
    CascadeMux I__2774 (
            .O(N__17158),
            .I(N__17142));
    CascadeMux I__2773 (
            .O(N__17157),
            .I(N__17137));
    CascadeMux I__2772 (
            .O(N__17156),
            .I(N__17133));
    InMux I__2771 (
            .O(N__17155),
            .I(N__17129));
    LocalMux I__2770 (
            .O(N__17152),
            .I(N__17126));
    CascadeMux I__2769 (
            .O(N__17151),
            .I(N__17120));
    CascadeMux I__2768 (
            .O(N__17150),
            .I(N__17116));
    InMux I__2767 (
            .O(N__17149),
            .I(N__17112));
    InMux I__2766 (
            .O(N__17148),
            .I(N__17107));
    InMux I__2765 (
            .O(N__17147),
            .I(N__17107));
    InMux I__2764 (
            .O(N__17146),
            .I(N__17096));
    InMux I__2763 (
            .O(N__17145),
            .I(N__17096));
    InMux I__2762 (
            .O(N__17142),
            .I(N__17096));
    InMux I__2761 (
            .O(N__17141),
            .I(N__17096));
    InMux I__2760 (
            .O(N__17140),
            .I(N__17096));
    InMux I__2759 (
            .O(N__17137),
            .I(N__17087));
    InMux I__2758 (
            .O(N__17136),
            .I(N__17087));
    InMux I__2757 (
            .O(N__17133),
            .I(N__17087));
    InMux I__2756 (
            .O(N__17132),
            .I(N__17087));
    LocalMux I__2755 (
            .O(N__17129),
            .I(N__17084));
    Span4Mux_h I__2754 (
            .O(N__17126),
            .I(N__17081));
    InMux I__2753 (
            .O(N__17125),
            .I(N__17074));
    InMux I__2752 (
            .O(N__17124),
            .I(N__17074));
    InMux I__2751 (
            .O(N__17123),
            .I(N__17074));
    InMux I__2750 (
            .O(N__17120),
            .I(N__17065));
    InMux I__2749 (
            .O(N__17119),
            .I(N__17065));
    InMux I__2748 (
            .O(N__17116),
            .I(N__17065));
    InMux I__2747 (
            .O(N__17115),
            .I(N__17065));
    LocalMux I__2746 (
            .O(N__17112),
            .I(\eeprom.n3331 ));
    LocalMux I__2745 (
            .O(N__17107),
            .I(\eeprom.n3331 ));
    LocalMux I__2744 (
            .O(N__17096),
            .I(\eeprom.n3331 ));
    LocalMux I__2743 (
            .O(N__17087),
            .I(\eeprom.n3331 ));
    Odrv4 I__2742 (
            .O(N__17084),
            .I(\eeprom.n3331 ));
    Odrv4 I__2741 (
            .O(N__17081),
            .I(\eeprom.n3331 ));
    LocalMux I__2740 (
            .O(N__17074),
            .I(\eeprom.n3331 ));
    LocalMux I__2739 (
            .O(N__17065),
            .I(\eeprom.n3331 ));
    CascadeMux I__2738 (
            .O(N__17048),
            .I(\eeprom.n3310_cascade_ ));
    InMux I__2737 (
            .O(N__17045),
            .I(N__17042));
    LocalMux I__2736 (
            .O(N__17042),
            .I(N__17039));
    Span4Mux_v I__2735 (
            .O(N__17039),
            .I(N__17036));
    Odrv4 I__2734 (
            .O(N__17036),
            .I(\eeprom.n3377 ));
    CascadeMux I__2733 (
            .O(N__17033),
            .I(N__17030));
    InMux I__2732 (
            .O(N__17030),
            .I(N__17026));
    CascadeMux I__2731 (
            .O(N__17029),
            .I(N__17023));
    LocalMux I__2730 (
            .O(N__17026),
            .I(N__17019));
    InMux I__2729 (
            .O(N__17023),
            .I(N__17014));
    InMux I__2728 (
            .O(N__17022),
            .I(N__17014));
    Span4Mux_h I__2727 (
            .O(N__17019),
            .I(N__17011));
    LocalMux I__2726 (
            .O(N__17014),
            .I(\eeprom.n3409 ));
    Odrv4 I__2725 (
            .O(N__17011),
            .I(\eeprom.n3409 ));
    InMux I__2724 (
            .O(N__17006),
            .I(N__17003));
    LocalMux I__2723 (
            .O(N__17003),
            .I(N__17000));
    Span4Mux_h I__2722 (
            .O(N__17000),
            .I(N__16997));
    Odrv4 I__2721 (
            .O(N__16997),
            .I(\eeprom.n3284 ));
    InMux I__2720 (
            .O(N__16994),
            .I(N__16991));
    LocalMux I__2719 (
            .O(N__16991),
            .I(N__16986));
    InMux I__2718 (
            .O(N__16990),
            .I(N__16983));
    CascadeMux I__2717 (
            .O(N__16989),
            .I(N__16980));
    Span4Mux_v I__2716 (
            .O(N__16986),
            .I(N__16977));
    LocalMux I__2715 (
            .O(N__16983),
            .I(N__16974));
    InMux I__2714 (
            .O(N__16980),
            .I(N__16971));
    Odrv4 I__2713 (
            .O(N__16977),
            .I(\eeprom.n3218 ));
    Odrv4 I__2712 (
            .O(N__16974),
            .I(\eeprom.n3218 ));
    LocalMux I__2711 (
            .O(N__16971),
            .I(\eeprom.n3218 ));
    InMux I__2710 (
            .O(N__16964),
            .I(N__16961));
    LocalMux I__2709 (
            .O(N__16961),
            .I(N__16958));
    Span4Mux_h I__2708 (
            .O(N__16958),
            .I(N__16955));
    Odrv4 I__2707 (
            .O(N__16955),
            .I(\eeprom.n3285 ));
    InMux I__2706 (
            .O(N__16952),
            .I(N__16948));
    InMux I__2705 (
            .O(N__16951),
            .I(N__16945));
    LocalMux I__2704 (
            .O(N__16948),
            .I(N__16942));
    LocalMux I__2703 (
            .O(N__16945),
            .I(N__16939));
    Odrv4 I__2702 (
            .O(N__16942),
            .I(\eeprom.n3317 ));
    Odrv4 I__2701 (
            .O(N__16939),
            .I(\eeprom.n3317 ));
    CascadeMux I__2700 (
            .O(N__16934),
            .I(N__16931));
    InMux I__2699 (
            .O(N__16931),
            .I(N__16928));
    LocalMux I__2698 (
            .O(N__16928),
            .I(N__16925));
    Span4Mux_h I__2697 (
            .O(N__16925),
            .I(N__16921));
    InMux I__2696 (
            .O(N__16924),
            .I(N__16918));
    Odrv4 I__2695 (
            .O(N__16921),
            .I(\eeprom.n3314 ));
    LocalMux I__2694 (
            .O(N__16918),
            .I(\eeprom.n3314 ));
    CascadeMux I__2693 (
            .O(N__16913),
            .I(\eeprom.n3317_cascade_ ));
    CascadeMux I__2692 (
            .O(N__16910),
            .I(N__16907));
    InMux I__2691 (
            .O(N__16907),
            .I(N__16902));
    InMux I__2690 (
            .O(N__16906),
            .I(N__16899));
    InMux I__2689 (
            .O(N__16905),
            .I(N__16896));
    LocalMux I__2688 (
            .O(N__16902),
            .I(N__16893));
    LocalMux I__2687 (
            .O(N__16899),
            .I(N__16890));
    LocalMux I__2686 (
            .O(N__16896),
            .I(N__16885));
    Span4Mux_h I__2685 (
            .O(N__16893),
            .I(N__16885));
    Odrv4 I__2684 (
            .O(N__16890),
            .I(\eeprom.n3316 ));
    Odrv4 I__2683 (
            .O(N__16885),
            .I(\eeprom.n3316 ));
    CascadeMux I__2682 (
            .O(N__16880),
            .I(N__16875));
    InMux I__2681 (
            .O(N__16879),
            .I(N__16872));
    InMux I__2680 (
            .O(N__16878),
            .I(N__16869));
    InMux I__2679 (
            .O(N__16875),
            .I(N__16866));
    LocalMux I__2678 (
            .O(N__16872),
            .I(N__16863));
    LocalMux I__2677 (
            .O(N__16869),
            .I(\eeprom.n3318 ));
    LocalMux I__2676 (
            .O(N__16866),
            .I(\eeprom.n3318 ));
    Odrv4 I__2675 (
            .O(N__16863),
            .I(\eeprom.n3318 ));
    CascadeMux I__2674 (
            .O(N__16856),
            .I(\eeprom.n5315_cascade_ ));
    InMux I__2673 (
            .O(N__16853),
            .I(N__16850));
    LocalMux I__2672 (
            .O(N__16850),
            .I(\eeprom.n5313 ));
    CascadeMux I__2671 (
            .O(N__16847),
            .I(N__16844));
    InMux I__2670 (
            .O(N__16844),
            .I(N__16841));
    LocalMux I__2669 (
            .O(N__16841),
            .I(N__16837));
    InMux I__2668 (
            .O(N__16840),
            .I(N__16833));
    Span4Mux_h I__2667 (
            .O(N__16837),
            .I(N__16830));
    InMux I__2666 (
            .O(N__16836),
            .I(N__16827));
    LocalMux I__2665 (
            .O(N__16833),
            .I(\eeprom.n3303 ));
    Odrv4 I__2664 (
            .O(N__16830),
            .I(\eeprom.n3303 ));
    LocalMux I__2663 (
            .O(N__16827),
            .I(\eeprom.n3303 ));
    CascadeMux I__2662 (
            .O(N__16820),
            .I(N__16816));
    InMux I__2661 (
            .O(N__16819),
            .I(N__16813));
    InMux I__2660 (
            .O(N__16816),
            .I(N__16810));
    LocalMux I__2659 (
            .O(N__16813),
            .I(N__16806));
    LocalMux I__2658 (
            .O(N__16810),
            .I(N__16803));
    InMux I__2657 (
            .O(N__16809),
            .I(N__16800));
    Odrv4 I__2656 (
            .O(N__16806),
            .I(\eeprom.n3304 ));
    Odrv4 I__2655 (
            .O(N__16803),
            .I(\eeprom.n3304 ));
    LocalMux I__2654 (
            .O(N__16800),
            .I(\eeprom.n3304 ));
    CascadeMux I__2653 (
            .O(N__16793),
            .I(\eeprom.n4820_cascade_ ));
    InMux I__2652 (
            .O(N__16790),
            .I(N__16786));
    InMux I__2651 (
            .O(N__16789),
            .I(N__16782));
    LocalMux I__2650 (
            .O(N__16786),
            .I(N__16779));
    CascadeMux I__2649 (
            .O(N__16785),
            .I(N__16776));
    LocalMux I__2648 (
            .O(N__16782),
            .I(N__16773));
    Span4Mux_h I__2647 (
            .O(N__16779),
            .I(N__16770));
    InMux I__2646 (
            .O(N__16776),
            .I(N__16767));
    Span4Mux_h I__2645 (
            .O(N__16773),
            .I(N__16764));
    Odrv4 I__2644 (
            .O(N__16770),
            .I(\eeprom.n3302 ));
    LocalMux I__2643 (
            .O(N__16767),
            .I(\eeprom.n3302 ));
    Odrv4 I__2642 (
            .O(N__16764),
            .I(\eeprom.n3302 ));
    InMux I__2641 (
            .O(N__16757),
            .I(N__16754));
    LocalMux I__2640 (
            .O(N__16754),
            .I(\eeprom.n26 ));
    CascadeMux I__2639 (
            .O(N__16751),
            .I(N__16747));
    CascadeMux I__2638 (
            .O(N__16750),
            .I(N__16744));
    InMux I__2637 (
            .O(N__16747),
            .I(N__16741));
    InMux I__2636 (
            .O(N__16744),
            .I(N__16738));
    LocalMux I__2635 (
            .O(N__16741),
            .I(N__16734));
    LocalMux I__2634 (
            .O(N__16738),
            .I(N__16731));
    InMux I__2633 (
            .O(N__16737),
            .I(N__16728));
    Span4Mux_v I__2632 (
            .O(N__16734),
            .I(N__16725));
    Odrv4 I__2631 (
            .O(N__16731),
            .I(\eeprom.n3405 ));
    LocalMux I__2630 (
            .O(N__16728),
            .I(\eeprom.n3405 ));
    Odrv4 I__2629 (
            .O(N__16725),
            .I(\eeprom.n3405 ));
    CascadeMux I__2628 (
            .O(N__16718),
            .I(\eeprom.n4824_cascade_ ));
    InMux I__2627 (
            .O(N__16715),
            .I(N__16711));
    InMux I__2626 (
            .O(N__16714),
            .I(N__16707));
    LocalMux I__2625 (
            .O(N__16711),
            .I(N__16704));
    CascadeMux I__2624 (
            .O(N__16710),
            .I(N__16701));
    LocalMux I__2623 (
            .O(N__16707),
            .I(N__16698));
    Span4Mux_v I__2622 (
            .O(N__16704),
            .I(N__16695));
    InMux I__2621 (
            .O(N__16701),
            .I(N__16692));
    Span4Mux_h I__2620 (
            .O(N__16698),
            .I(N__16689));
    Odrv4 I__2619 (
            .O(N__16695),
            .I(\eeprom.n3404 ));
    LocalMux I__2618 (
            .O(N__16692),
            .I(\eeprom.n3404 ));
    Odrv4 I__2617 (
            .O(N__16689),
            .I(\eeprom.n3404 ));
    InMux I__2616 (
            .O(N__16682),
            .I(N__16679));
    LocalMux I__2615 (
            .O(N__16679),
            .I(\eeprom.n28_adj_261 ));
    InMux I__2614 (
            .O(N__16676),
            .I(N__16673));
    LocalMux I__2613 (
            .O(N__16673),
            .I(N__16670));
    Span4Mux_h I__2612 (
            .O(N__16670),
            .I(N__16667));
    Odrv4 I__2611 (
            .O(N__16667),
            .I(\eeprom.n3386 ));
    CascadeMux I__2610 (
            .O(N__16664),
            .I(N__16661));
    InMux I__2609 (
            .O(N__16661),
            .I(N__16658));
    LocalMux I__2608 (
            .O(N__16658),
            .I(N__16653));
    InMux I__2607 (
            .O(N__16657),
            .I(N__16650));
    InMux I__2606 (
            .O(N__16656),
            .I(N__16647));
    Span4Mux_h I__2605 (
            .O(N__16653),
            .I(N__16644));
    LocalMux I__2604 (
            .O(N__16650),
            .I(\eeprom.n3418 ));
    LocalMux I__2603 (
            .O(N__16647),
            .I(\eeprom.n3418 ));
    Odrv4 I__2602 (
            .O(N__16644),
            .I(\eeprom.n3418 ));
    InMux I__2601 (
            .O(N__16637),
            .I(N__16634));
    LocalMux I__2600 (
            .O(N__16634),
            .I(N__16631));
    Span4Mux_v I__2599 (
            .O(N__16631),
            .I(N__16628));
    Odrv4 I__2598 (
            .O(N__16628),
            .I(\eeprom.n3384 ));
    CascadeMux I__2597 (
            .O(N__16625),
            .I(N__16622));
    InMux I__2596 (
            .O(N__16622),
            .I(N__16619));
    LocalMux I__2595 (
            .O(N__16619),
            .I(N__16614));
    InMux I__2594 (
            .O(N__16618),
            .I(N__16611));
    InMux I__2593 (
            .O(N__16617),
            .I(N__16608));
    Span4Mux_h I__2592 (
            .O(N__16614),
            .I(N__16605));
    LocalMux I__2591 (
            .O(N__16611),
            .I(\eeprom.n3416 ));
    LocalMux I__2590 (
            .O(N__16608),
            .I(\eeprom.n3416 ));
    Odrv4 I__2589 (
            .O(N__16605),
            .I(\eeprom.n3416 ));
    CascadeMux I__2588 (
            .O(N__16598),
            .I(N__16595));
    InMux I__2587 (
            .O(N__16595),
            .I(N__16592));
    LocalMux I__2586 (
            .O(N__16592),
            .I(N__16589));
    Span4Mux_v I__2585 (
            .O(N__16589),
            .I(N__16586));
    Odrv4 I__2584 (
            .O(N__16586),
            .I(\eeprom.n3383 ));
    CascadeMux I__2583 (
            .O(N__16583),
            .I(N__16579));
    InMux I__2582 (
            .O(N__16582),
            .I(N__16576));
    InMux I__2581 (
            .O(N__16579),
            .I(N__16573));
    LocalMux I__2580 (
            .O(N__16576),
            .I(N__16569));
    LocalMux I__2579 (
            .O(N__16573),
            .I(N__16566));
    InMux I__2578 (
            .O(N__16572),
            .I(N__16563));
    Odrv4 I__2577 (
            .O(N__16569),
            .I(\eeprom.n3313 ));
    Odrv4 I__2576 (
            .O(N__16566),
            .I(\eeprom.n3313 ));
    LocalMux I__2575 (
            .O(N__16563),
            .I(\eeprom.n3313 ));
    CascadeMux I__2574 (
            .O(N__16556),
            .I(N__16553));
    InMux I__2573 (
            .O(N__16553),
            .I(N__16550));
    LocalMux I__2572 (
            .O(N__16550),
            .I(N__16547));
    Span4Mux_h I__2571 (
            .O(N__16547),
            .I(N__16544));
    Odrv4 I__2570 (
            .O(N__16544),
            .I(\eeprom.n3371 ));
    CascadeMux I__2569 (
            .O(N__16541),
            .I(N__16538));
    InMux I__2568 (
            .O(N__16538),
            .I(N__16535));
    LocalMux I__2567 (
            .O(N__16535),
            .I(N__16532));
    Span4Mux_h I__2566 (
            .O(N__16532),
            .I(N__16529));
    Odrv4 I__2565 (
            .O(N__16529),
            .I(\eeprom.n3282 ));
    InMux I__2564 (
            .O(N__16526),
            .I(N__16523));
    LocalMux I__2563 (
            .O(N__16523),
            .I(N__16520));
    Span4Mux_h I__2562 (
            .O(N__16520),
            .I(N__16517));
    Odrv4 I__2561 (
            .O(N__16517),
            .I(\eeprom.n3381 ));
    CascadeMux I__2560 (
            .O(N__16514),
            .I(\eeprom.n3314_cascade_ ));
    CascadeMux I__2559 (
            .O(N__16511),
            .I(N__16507));
    InMux I__2558 (
            .O(N__16510),
            .I(N__16504));
    InMux I__2557 (
            .O(N__16507),
            .I(N__16501));
    LocalMux I__2556 (
            .O(N__16504),
            .I(N__16496));
    LocalMux I__2555 (
            .O(N__16501),
            .I(N__16496));
    Span4Mux_h I__2554 (
            .O(N__16496),
            .I(N__16493));
    Odrv4 I__2553 (
            .O(N__16493),
            .I(\eeprom.n3413 ));
    InMux I__2552 (
            .O(N__16490),
            .I(\eeprom.n4222 ));
    CascadeMux I__2551 (
            .O(N__16487),
            .I(N__16482));
    InMux I__2550 (
            .O(N__16486),
            .I(N__16479));
    InMux I__2549 (
            .O(N__16485),
            .I(N__16476));
    InMux I__2548 (
            .O(N__16482),
            .I(N__16473));
    LocalMux I__2547 (
            .O(N__16479),
            .I(\eeprom.n3500 ));
    LocalMux I__2546 (
            .O(N__16476),
            .I(\eeprom.n3500 ));
    LocalMux I__2545 (
            .O(N__16473),
            .I(\eeprom.n3500 ));
    InMux I__2544 (
            .O(N__16466),
            .I(N__16463));
    LocalMux I__2543 (
            .O(N__16463),
            .I(N__16460));
    Odrv4 I__2542 (
            .O(N__16460),
            .I(\eeprom.n3567 ));
    InMux I__2541 (
            .O(N__16457),
            .I(\eeprom.n4223 ));
    CascadeMux I__2540 (
            .O(N__16454),
            .I(N__16450));
    InMux I__2539 (
            .O(N__16453),
            .I(N__16446));
    InMux I__2538 (
            .O(N__16450),
            .I(N__16443));
    InMux I__2537 (
            .O(N__16449),
            .I(N__16440));
    LocalMux I__2536 (
            .O(N__16446),
            .I(\eeprom.n3499 ));
    LocalMux I__2535 (
            .O(N__16443),
            .I(\eeprom.n3499 ));
    LocalMux I__2534 (
            .O(N__16440),
            .I(\eeprom.n3499 ));
    InMux I__2533 (
            .O(N__16433),
            .I(N__16430));
    LocalMux I__2532 (
            .O(N__16430),
            .I(\eeprom.n3566 ));
    InMux I__2531 (
            .O(N__16427),
            .I(\eeprom.n4224 ));
    InMux I__2530 (
            .O(N__16424),
            .I(N__16421));
    LocalMux I__2529 (
            .O(N__16421),
            .I(N__16417));
    CascadeMux I__2528 (
            .O(N__16420),
            .I(N__16414));
    Span4Mux_h I__2527 (
            .O(N__16417),
            .I(N__16411));
    InMux I__2526 (
            .O(N__16414),
            .I(N__16408));
    Odrv4 I__2525 (
            .O(N__16411),
            .I(\eeprom.n3498 ));
    LocalMux I__2524 (
            .O(N__16408),
            .I(\eeprom.n3498 ));
    InMux I__2523 (
            .O(N__16403),
            .I(N__16400));
    LocalMux I__2522 (
            .O(N__16400),
            .I(N__16397));
    Odrv4 I__2521 (
            .O(N__16397),
            .I(\eeprom.n3565 ));
    InMux I__2520 (
            .O(N__16394),
            .I(\eeprom.n4225 ));
    InMux I__2519 (
            .O(N__16391),
            .I(N__16387));
    InMux I__2518 (
            .O(N__16390),
            .I(N__16384));
    LocalMux I__2517 (
            .O(N__16387),
            .I(N__16381));
    LocalMux I__2516 (
            .O(N__16384),
            .I(N__16377));
    Span4Mux_h I__2515 (
            .O(N__16381),
            .I(N__16374));
    InMux I__2514 (
            .O(N__16380),
            .I(N__16371));
    Odrv4 I__2513 (
            .O(N__16377),
            .I(\eeprom.n3497 ));
    Odrv4 I__2512 (
            .O(N__16374),
            .I(\eeprom.n3497 ));
    LocalMux I__2511 (
            .O(N__16371),
            .I(\eeprom.n3497 ));
    InMux I__2510 (
            .O(N__16364),
            .I(N__16361));
    LocalMux I__2509 (
            .O(N__16361),
            .I(\eeprom.n3564 ));
    InMux I__2508 (
            .O(N__16358),
            .I(\eeprom.n4226 ));
    InMux I__2507 (
            .O(N__16355),
            .I(N__16352));
    LocalMux I__2506 (
            .O(N__16352),
            .I(N__16348));
    InMux I__2505 (
            .O(N__16351),
            .I(N__16345));
    Span4Mux_v I__2504 (
            .O(N__16348),
            .I(N__16340));
    LocalMux I__2503 (
            .O(N__16345),
            .I(N__16340));
    Span4Mux_h I__2502 (
            .O(N__16340),
            .I(N__16337));
    Odrv4 I__2501 (
            .O(N__16337),
            .I(\eeprom.n3496 ));
    CascadeMux I__2500 (
            .O(N__16334),
            .I(N__16331));
    InMux I__2499 (
            .O(N__16331),
            .I(N__16325));
    InMux I__2498 (
            .O(N__16330),
            .I(N__16314));
    InMux I__2497 (
            .O(N__16329),
            .I(N__16314));
    InMux I__2496 (
            .O(N__16328),
            .I(N__16311));
    LocalMux I__2495 (
            .O(N__16325),
            .I(N__16308));
    CascadeMux I__2494 (
            .O(N__16324),
            .I(N__16305));
    CascadeMux I__2493 (
            .O(N__16323),
            .I(N__16302));
    CascadeMux I__2492 (
            .O(N__16322),
            .I(N__16294));
    CascadeMux I__2491 (
            .O(N__16321),
            .I(N__16291));
    CascadeMux I__2490 (
            .O(N__16320),
            .I(N__16286));
    CascadeMux I__2489 (
            .O(N__16319),
            .I(N__16280));
    LocalMux I__2488 (
            .O(N__16314),
            .I(N__16274));
    LocalMux I__2487 (
            .O(N__16311),
            .I(N__16269));
    Span4Mux_h I__2486 (
            .O(N__16308),
            .I(N__16269));
    InMux I__2485 (
            .O(N__16305),
            .I(N__16260));
    InMux I__2484 (
            .O(N__16302),
            .I(N__16260));
    InMux I__2483 (
            .O(N__16301),
            .I(N__16260));
    InMux I__2482 (
            .O(N__16300),
            .I(N__16260));
    InMux I__2481 (
            .O(N__16299),
            .I(N__16247));
    InMux I__2480 (
            .O(N__16298),
            .I(N__16247));
    InMux I__2479 (
            .O(N__16297),
            .I(N__16247));
    InMux I__2478 (
            .O(N__16294),
            .I(N__16247));
    InMux I__2477 (
            .O(N__16291),
            .I(N__16247));
    InMux I__2476 (
            .O(N__16290),
            .I(N__16247));
    InMux I__2475 (
            .O(N__16289),
            .I(N__16236));
    InMux I__2474 (
            .O(N__16286),
            .I(N__16236));
    InMux I__2473 (
            .O(N__16285),
            .I(N__16236));
    InMux I__2472 (
            .O(N__16284),
            .I(N__16236));
    InMux I__2471 (
            .O(N__16283),
            .I(N__16236));
    InMux I__2470 (
            .O(N__16280),
            .I(N__16227));
    InMux I__2469 (
            .O(N__16279),
            .I(N__16227));
    InMux I__2468 (
            .O(N__16278),
            .I(N__16227));
    InMux I__2467 (
            .O(N__16277),
            .I(N__16227));
    Odrv4 I__2466 (
            .O(N__16274),
            .I(\eeprom.n3529 ));
    Odrv4 I__2465 (
            .O(N__16269),
            .I(\eeprom.n3529 ));
    LocalMux I__2464 (
            .O(N__16260),
            .I(\eeprom.n3529 ));
    LocalMux I__2463 (
            .O(N__16247),
            .I(\eeprom.n3529 ));
    LocalMux I__2462 (
            .O(N__16236),
            .I(\eeprom.n3529 ));
    LocalMux I__2461 (
            .O(N__16227),
            .I(\eeprom.n3529 ));
    InMux I__2460 (
            .O(N__16214),
            .I(\eeprom.n4227 ));
    InMux I__2459 (
            .O(N__16211),
            .I(N__16208));
    LocalMux I__2458 (
            .O(N__16208),
            .I(N__16205));
    Span4Mux_h I__2457 (
            .O(N__16205),
            .I(N__16202));
    Odrv4 I__2456 (
            .O(N__16202),
            .I(\eeprom.n5355 ));
    InMux I__2455 (
            .O(N__16199),
            .I(N__16196));
    LocalMux I__2454 (
            .O(N__16196),
            .I(N__16193));
    Span4Mux_h I__2453 (
            .O(N__16193),
            .I(N__16190));
    Odrv4 I__2452 (
            .O(N__16190),
            .I(\eeprom.n3382 ));
    CascadeMux I__2451 (
            .O(N__16187),
            .I(N__16184));
    InMux I__2450 (
            .O(N__16184),
            .I(N__16180));
    InMux I__2449 (
            .O(N__16183),
            .I(N__16177));
    LocalMux I__2448 (
            .O(N__16180),
            .I(N__16172));
    LocalMux I__2447 (
            .O(N__16177),
            .I(N__16172));
    Span4Mux_v I__2446 (
            .O(N__16172),
            .I(N__16169));
    Odrv4 I__2445 (
            .O(N__16169),
            .I(\eeprom.n3414 ));
    CascadeMux I__2444 (
            .O(N__16166),
            .I(N__16162));
    InMux I__2443 (
            .O(N__16165),
            .I(N__16159));
    InMux I__2442 (
            .O(N__16162),
            .I(N__16156));
    LocalMux I__2441 (
            .O(N__16159),
            .I(N__16152));
    LocalMux I__2440 (
            .O(N__16156),
            .I(N__16149));
    InMux I__2439 (
            .O(N__16155),
            .I(N__16146));
    Span4Mux_h I__2438 (
            .O(N__16152),
            .I(N__16141));
    Span4Mux_h I__2437 (
            .O(N__16149),
            .I(N__16141));
    LocalMux I__2436 (
            .O(N__16146),
            .I(\eeprom.n3417 ));
    Odrv4 I__2435 (
            .O(N__16141),
            .I(\eeprom.n3417 ));
    CascadeMux I__2434 (
            .O(N__16136),
            .I(\eeprom.n3414_cascade_ ));
    CascadeMux I__2433 (
            .O(N__16133),
            .I(\eeprom.n5291_cascade_ ));
    InMux I__2432 (
            .O(N__16130),
            .I(N__16125));
    InMux I__2431 (
            .O(N__16129),
            .I(N__16122));
    InMux I__2430 (
            .O(N__16128),
            .I(N__16119));
    LocalMux I__2429 (
            .O(N__16125),
            .I(N__16116));
    LocalMux I__2428 (
            .O(N__16122),
            .I(N__16113));
    LocalMux I__2427 (
            .O(N__16119),
            .I(N__16110));
    Span4Mux_h I__2426 (
            .O(N__16116),
            .I(N__16105));
    Span4Mux_h I__2425 (
            .O(N__16113),
            .I(N__16105));
    Odrv4 I__2424 (
            .O(N__16110),
            .I(\eeprom.n3508 ));
    Odrv4 I__2423 (
            .O(N__16105),
            .I(\eeprom.n3508 ));
    InMux I__2422 (
            .O(N__16100),
            .I(N__16097));
    LocalMux I__2421 (
            .O(N__16097),
            .I(\eeprom.n3575 ));
    InMux I__2420 (
            .O(N__16094),
            .I(\eeprom.n4215 ));
    InMux I__2419 (
            .O(N__16091),
            .I(N__16087));
    InMux I__2418 (
            .O(N__16090),
            .I(N__16084));
    LocalMux I__2417 (
            .O(N__16087),
            .I(N__16079));
    LocalMux I__2416 (
            .O(N__16084),
            .I(N__16079));
    Span4Mux_h I__2415 (
            .O(N__16079),
            .I(N__16076));
    Odrv4 I__2414 (
            .O(N__16076),
            .I(\eeprom.n3507 ));
    InMux I__2413 (
            .O(N__16073),
            .I(N__16070));
    LocalMux I__2412 (
            .O(N__16070),
            .I(\eeprom.n3574 ));
    InMux I__2411 (
            .O(N__16067),
            .I(\eeprom.n4216 ));
    InMux I__2410 (
            .O(N__16064),
            .I(N__16059));
    InMux I__2409 (
            .O(N__16063),
            .I(N__16056));
    InMux I__2408 (
            .O(N__16062),
            .I(N__16053));
    LocalMux I__2407 (
            .O(N__16059),
            .I(\eeprom.n3506 ));
    LocalMux I__2406 (
            .O(N__16056),
            .I(\eeprom.n3506 ));
    LocalMux I__2405 (
            .O(N__16053),
            .I(\eeprom.n3506 ));
    InMux I__2404 (
            .O(N__16046),
            .I(N__16043));
    LocalMux I__2403 (
            .O(N__16043),
            .I(N__16040));
    Span4Mux_h I__2402 (
            .O(N__16040),
            .I(N__16037));
    Odrv4 I__2401 (
            .O(N__16037),
            .I(\eeprom.n3573 ));
    InMux I__2400 (
            .O(N__16034),
            .I(\eeprom.n4217 ));
    InMux I__2399 (
            .O(N__16031),
            .I(N__16027));
    InMux I__2398 (
            .O(N__16030),
            .I(N__16024));
    LocalMux I__2397 (
            .O(N__16027),
            .I(N__16021));
    LocalMux I__2396 (
            .O(N__16024),
            .I(N__16018));
    Odrv4 I__2395 (
            .O(N__16021),
            .I(\eeprom.n3505 ));
    Odrv4 I__2394 (
            .O(N__16018),
            .I(\eeprom.n3505 ));
    InMux I__2393 (
            .O(N__16013),
            .I(N__16010));
    LocalMux I__2392 (
            .O(N__16010),
            .I(\eeprom.n3572 ));
    InMux I__2391 (
            .O(N__16007),
            .I(\eeprom.n4218 ));
    InMux I__2390 (
            .O(N__16004),
            .I(N__16000));
    InMux I__2389 (
            .O(N__16003),
            .I(N__15997));
    LocalMux I__2388 (
            .O(N__16000),
            .I(N__15994));
    LocalMux I__2387 (
            .O(N__15997),
            .I(N__15990));
    Span4Mux_v I__2386 (
            .O(N__15994),
            .I(N__15987));
    InMux I__2385 (
            .O(N__15993),
            .I(N__15984));
    Odrv4 I__2384 (
            .O(N__15990),
            .I(\eeprom.n3504 ));
    Odrv4 I__2383 (
            .O(N__15987),
            .I(\eeprom.n3504 ));
    LocalMux I__2382 (
            .O(N__15984),
            .I(\eeprom.n3504 ));
    InMux I__2381 (
            .O(N__15977),
            .I(N__15974));
    LocalMux I__2380 (
            .O(N__15974),
            .I(\eeprom.n3571 ));
    InMux I__2379 (
            .O(N__15971),
            .I(\eeprom.n4219 ));
    InMux I__2378 (
            .O(N__15968),
            .I(N__15965));
    LocalMux I__2377 (
            .O(N__15965),
            .I(N__15962));
    Span4Mux_h I__2376 (
            .O(N__15962),
            .I(N__15957));
    InMux I__2375 (
            .O(N__15961),
            .I(N__15952));
    InMux I__2374 (
            .O(N__15960),
            .I(N__15952));
    Odrv4 I__2373 (
            .O(N__15957),
            .I(\eeprom.n3503 ));
    LocalMux I__2372 (
            .O(N__15952),
            .I(\eeprom.n3503 ));
    InMux I__2371 (
            .O(N__15947),
            .I(N__15944));
    LocalMux I__2370 (
            .O(N__15944),
            .I(N__15941));
    Odrv4 I__2369 (
            .O(N__15941),
            .I(\eeprom.n3570 ));
    InMux I__2368 (
            .O(N__15938),
            .I(bfn_20_21_0_));
    InMux I__2367 (
            .O(N__15935),
            .I(N__15932));
    LocalMux I__2366 (
            .O(N__15932),
            .I(N__15929));
    Span4Mux_h I__2365 (
            .O(N__15929),
            .I(N__15926));
    Odrv4 I__2364 (
            .O(N__15926),
            .I(\eeprom.n3569 ));
    InMux I__2363 (
            .O(N__15923),
            .I(\eeprom.n4221 ));
    InMux I__2362 (
            .O(N__15920),
            .I(N__15917));
    LocalMux I__2361 (
            .O(N__15917),
            .I(N__15912));
    InMux I__2360 (
            .O(N__15916),
            .I(N__15909));
    InMux I__2359 (
            .O(N__15915),
            .I(N__15906));
    Span4Mux_v I__2358 (
            .O(N__15912),
            .I(N__15901));
    LocalMux I__2357 (
            .O(N__15909),
            .I(N__15901));
    LocalMux I__2356 (
            .O(N__15906),
            .I(N__15898));
    Odrv4 I__2355 (
            .O(N__15901),
            .I(\eeprom.n3501 ));
    Odrv12 I__2354 (
            .O(N__15898),
            .I(\eeprom.n3501 ));
    InMux I__2353 (
            .O(N__15893),
            .I(N__15890));
    LocalMux I__2352 (
            .O(N__15890),
            .I(N__15887));
    Odrv4 I__2351 (
            .O(N__15887),
            .I(\eeprom.n3568 ));
    CascadeMux I__2350 (
            .O(N__15884),
            .I(N__15881));
    InMux I__2349 (
            .O(N__15881),
            .I(N__15877));
    InMux I__2348 (
            .O(N__15880),
            .I(N__15874));
    LocalMux I__2347 (
            .O(N__15877),
            .I(N__15871));
    LocalMux I__2346 (
            .O(N__15874),
            .I(N__15867));
    Span4Mux_v I__2345 (
            .O(N__15871),
            .I(N__15864));
    InMux I__2344 (
            .O(N__15870),
            .I(N__15861));
    Odrv4 I__2343 (
            .O(N__15867),
            .I(\eeprom.n3516 ));
    Odrv4 I__2342 (
            .O(N__15864),
            .I(\eeprom.n3516 ));
    LocalMux I__2341 (
            .O(N__15861),
            .I(\eeprom.n3516 ));
    InMux I__2340 (
            .O(N__15854),
            .I(N__15851));
    LocalMux I__2339 (
            .O(N__15851),
            .I(N__15848));
    Odrv4 I__2338 (
            .O(N__15848),
            .I(\eeprom.n3583 ));
    InMux I__2337 (
            .O(N__15845),
            .I(\eeprom.n4207 ));
    CascadeMux I__2336 (
            .O(N__15842),
            .I(N__15838));
    InMux I__2335 (
            .O(N__15841),
            .I(N__15835));
    InMux I__2334 (
            .O(N__15838),
            .I(N__15832));
    LocalMux I__2333 (
            .O(N__15835),
            .I(N__15828));
    LocalMux I__2332 (
            .O(N__15832),
            .I(N__15825));
    InMux I__2331 (
            .O(N__15831),
            .I(N__15822));
    Odrv4 I__2330 (
            .O(N__15828),
            .I(\eeprom.n3515 ));
    Odrv4 I__2329 (
            .O(N__15825),
            .I(\eeprom.n3515 ));
    LocalMux I__2328 (
            .O(N__15822),
            .I(\eeprom.n3515 ));
    CascadeMux I__2327 (
            .O(N__15815),
            .I(N__15812));
    InMux I__2326 (
            .O(N__15812),
            .I(N__15809));
    LocalMux I__2325 (
            .O(N__15809),
            .I(N__15806));
    Odrv4 I__2324 (
            .O(N__15806),
            .I(\eeprom.n3582 ));
    InMux I__2323 (
            .O(N__15803),
            .I(\eeprom.n4208 ));
    CascadeMux I__2322 (
            .O(N__15800),
            .I(N__15797));
    InMux I__2321 (
            .O(N__15797),
            .I(N__15794));
    LocalMux I__2320 (
            .O(N__15794),
            .I(N__15790));
    InMux I__2319 (
            .O(N__15793),
            .I(N__15787));
    Span4Mux_h I__2318 (
            .O(N__15790),
            .I(N__15784));
    LocalMux I__2317 (
            .O(N__15787),
            .I(\eeprom.n3514 ));
    Odrv4 I__2316 (
            .O(N__15784),
            .I(\eeprom.n3514 ));
    InMux I__2315 (
            .O(N__15779),
            .I(N__15776));
    LocalMux I__2314 (
            .O(N__15776),
            .I(N__15773));
    Span4Mux_v I__2313 (
            .O(N__15773),
            .I(N__15770));
    Odrv4 I__2312 (
            .O(N__15770),
            .I(\eeprom.n3581_adj_292 ));
    InMux I__2311 (
            .O(N__15767),
            .I(\eeprom.n4209 ));
    CascadeMux I__2310 (
            .O(N__15764),
            .I(N__15761));
    InMux I__2309 (
            .O(N__15761),
            .I(N__15758));
    LocalMux I__2308 (
            .O(N__15758),
            .I(N__15754));
    InMux I__2307 (
            .O(N__15757),
            .I(N__15751));
    Span4Mux_h I__2306 (
            .O(N__15754),
            .I(N__15748));
    LocalMux I__2305 (
            .O(N__15751),
            .I(\eeprom.n3513 ));
    Odrv4 I__2304 (
            .O(N__15748),
            .I(\eeprom.n3513 ));
    InMux I__2303 (
            .O(N__15743),
            .I(N__15740));
    LocalMux I__2302 (
            .O(N__15740),
            .I(N__15737));
    Odrv4 I__2301 (
            .O(N__15737),
            .I(\eeprom.n3580 ));
    InMux I__2300 (
            .O(N__15734),
            .I(\eeprom.n4210 ));
    CascadeMux I__2299 (
            .O(N__15731),
            .I(N__15728));
    InMux I__2298 (
            .O(N__15728),
            .I(N__15724));
    InMux I__2297 (
            .O(N__15727),
            .I(N__15721));
    LocalMux I__2296 (
            .O(N__15724),
            .I(N__15718));
    LocalMux I__2295 (
            .O(N__15721),
            .I(\eeprom.n3512 ));
    Odrv4 I__2294 (
            .O(N__15718),
            .I(\eeprom.n3512 ));
    InMux I__2293 (
            .O(N__15713),
            .I(N__15710));
    LocalMux I__2292 (
            .O(N__15710),
            .I(N__15707));
    Span4Mux_h I__2291 (
            .O(N__15707),
            .I(N__15704));
    Odrv4 I__2290 (
            .O(N__15704),
            .I(\eeprom.n3579 ));
    InMux I__2289 (
            .O(N__15701),
            .I(\eeprom.n4211 ));
    CascadeMux I__2288 (
            .O(N__15698),
            .I(N__15695));
    InMux I__2287 (
            .O(N__15695),
            .I(N__15692));
    LocalMux I__2286 (
            .O(N__15692),
            .I(N__15687));
    InMux I__2285 (
            .O(N__15691),
            .I(N__15684));
    InMux I__2284 (
            .O(N__15690),
            .I(N__15681));
    Span4Mux_v I__2283 (
            .O(N__15687),
            .I(N__15678));
    LocalMux I__2282 (
            .O(N__15684),
            .I(\eeprom.n3511 ));
    LocalMux I__2281 (
            .O(N__15681),
            .I(\eeprom.n3511 ));
    Odrv4 I__2280 (
            .O(N__15678),
            .I(\eeprom.n3511 ));
    InMux I__2279 (
            .O(N__15671),
            .I(N__15668));
    LocalMux I__2278 (
            .O(N__15668),
            .I(\eeprom.n3578 ));
    InMux I__2277 (
            .O(N__15665),
            .I(bfn_20_20_0_));
    CascadeMux I__2276 (
            .O(N__15662),
            .I(N__15659));
    InMux I__2275 (
            .O(N__15659),
            .I(N__15656));
    LocalMux I__2274 (
            .O(N__15656),
            .I(N__15651));
    InMux I__2273 (
            .O(N__15655),
            .I(N__15648));
    InMux I__2272 (
            .O(N__15654),
            .I(N__15645));
    Span4Mux_v I__2271 (
            .O(N__15651),
            .I(N__15642));
    LocalMux I__2270 (
            .O(N__15648),
            .I(\eeprom.n3510 ));
    LocalMux I__2269 (
            .O(N__15645),
            .I(\eeprom.n3510 ));
    Odrv4 I__2268 (
            .O(N__15642),
            .I(\eeprom.n3510 ));
    CascadeMux I__2267 (
            .O(N__15635),
            .I(N__15632));
    InMux I__2266 (
            .O(N__15632),
            .I(N__15629));
    LocalMux I__2265 (
            .O(N__15629),
            .I(\eeprom.n3577 ));
    InMux I__2264 (
            .O(N__15626),
            .I(\eeprom.n4213 ));
    CascadeMux I__2263 (
            .O(N__15623),
            .I(N__15620));
    InMux I__2262 (
            .O(N__15620),
            .I(N__15616));
    CascadeMux I__2261 (
            .O(N__15619),
            .I(N__15613));
    LocalMux I__2260 (
            .O(N__15616),
            .I(N__15610));
    InMux I__2259 (
            .O(N__15613),
            .I(N__15606));
    Span4Mux_h I__2258 (
            .O(N__15610),
            .I(N__15603));
    InMux I__2257 (
            .O(N__15609),
            .I(N__15600));
    LocalMux I__2256 (
            .O(N__15606),
            .I(\eeprom.n3509 ));
    Odrv4 I__2255 (
            .O(N__15603),
            .I(\eeprom.n3509 ));
    LocalMux I__2254 (
            .O(N__15600),
            .I(\eeprom.n3509 ));
    InMux I__2253 (
            .O(N__15593),
            .I(N__15590));
    LocalMux I__2252 (
            .O(N__15590),
            .I(\eeprom.n3576 ));
    InMux I__2251 (
            .O(N__15587),
            .I(\eeprom.n4214 ));
    InMux I__2250 (
            .O(N__15584),
            .I(N__15581));
    LocalMux I__2249 (
            .O(N__15581),
            .I(\eeprom.n5559 ));
    CascadeMux I__2248 (
            .O(N__15578),
            .I(N__15575));
    InMux I__2247 (
            .O(N__15575),
            .I(N__15572));
    LocalMux I__2246 (
            .O(N__15572),
            .I(\eeprom.n3714 ));
    InMux I__2245 (
            .O(N__15569),
            .I(\eeprom.n4238 ));
    InMux I__2244 (
            .O(N__15566),
            .I(N__15563));
    LocalMux I__2243 (
            .O(N__15563),
            .I(N__15560));
    Odrv4 I__2242 (
            .O(N__15560),
            .I(\eeprom.n5562 ));
    CascadeMux I__2241 (
            .O(N__15557),
            .I(N__15554));
    InMux I__2240 (
            .O(N__15554),
            .I(N__15551));
    LocalMux I__2239 (
            .O(N__15551),
            .I(N__15548));
    Odrv4 I__2238 (
            .O(N__15548),
            .I(\eeprom.n3713 ));
    InMux I__2237 (
            .O(N__15545),
            .I(\eeprom.n4239 ));
    InMux I__2236 (
            .O(N__15542),
            .I(N__15539));
    LocalMux I__2235 (
            .O(N__15539),
            .I(\eeprom.n5565 ));
    CascadeMux I__2234 (
            .O(N__15536),
            .I(N__15533));
    InMux I__2233 (
            .O(N__15533),
            .I(N__15530));
    LocalMux I__2232 (
            .O(N__15530),
            .I(\eeprom.n3712 ));
    InMux I__2231 (
            .O(N__15527),
            .I(\eeprom.n4240 ));
    InMux I__2230 (
            .O(N__15524),
            .I(N__15521));
    LocalMux I__2229 (
            .O(N__15521),
            .I(\eeprom.n3711 ));
    CascadeMux I__2228 (
            .O(N__15518),
            .I(N__15515));
    InMux I__2227 (
            .O(N__15515),
            .I(N__15512));
    LocalMux I__2226 (
            .O(N__15512),
            .I(N__15509));
    Span4Mux_h I__2225 (
            .O(N__15509),
            .I(N__15506));
    Odrv4 I__2224 (
            .O(N__15506),
            .I(\eeprom.n5568 ));
    InMux I__2223 (
            .O(N__15503),
            .I(\eeprom.n4241 ));
    InMux I__2222 (
            .O(N__15500),
            .I(N__15494));
    InMux I__2221 (
            .O(N__15499),
            .I(N__15494));
    LocalMux I__2220 (
            .O(N__15494),
            .I(\eeprom.n3716 ));
    InMux I__2219 (
            .O(N__15491),
            .I(N__15488));
    LocalMux I__2218 (
            .O(N__15488),
            .I(\eeprom.n5553 ));
    InMux I__2217 (
            .O(N__15485),
            .I(N__15482));
    LocalMux I__2216 (
            .O(N__15482),
            .I(N__15479));
    Span4Mux_v I__2215 (
            .O(N__15479),
            .I(N__15476));
    Odrv4 I__2214 (
            .O(N__15476),
            .I(\eeprom.n3586 ));
    InMux I__2213 (
            .O(N__15473),
            .I(bfn_20_19_0_));
    CascadeMux I__2212 (
            .O(N__15470),
            .I(N__15466));
    InMux I__2211 (
            .O(N__15469),
            .I(N__15462));
    InMux I__2210 (
            .O(N__15466),
            .I(N__15459));
    InMux I__2209 (
            .O(N__15465),
            .I(N__15456));
    LocalMux I__2208 (
            .O(N__15462),
            .I(\eeprom.n3518 ));
    LocalMux I__2207 (
            .O(N__15459),
            .I(\eeprom.n3518 ));
    LocalMux I__2206 (
            .O(N__15456),
            .I(\eeprom.n3518 ));
    CascadeMux I__2205 (
            .O(N__15449),
            .I(N__15446));
    InMux I__2204 (
            .O(N__15446),
            .I(N__15443));
    LocalMux I__2203 (
            .O(N__15443),
            .I(\eeprom.n3585_adj_296 ));
    InMux I__2202 (
            .O(N__15440),
            .I(\eeprom.n4205 ));
    CascadeMux I__2201 (
            .O(N__15437),
            .I(N__15433));
    InMux I__2200 (
            .O(N__15436),
            .I(N__15430));
    InMux I__2199 (
            .O(N__15433),
            .I(N__15427));
    LocalMux I__2198 (
            .O(N__15430),
            .I(N__15423));
    LocalMux I__2197 (
            .O(N__15427),
            .I(N__15420));
    InMux I__2196 (
            .O(N__15426),
            .I(N__15417));
    Odrv4 I__2195 (
            .O(N__15423),
            .I(\eeprom.n3517 ));
    Odrv4 I__2194 (
            .O(N__15420),
            .I(\eeprom.n3517 ));
    LocalMux I__2193 (
            .O(N__15417),
            .I(\eeprom.n3517 ));
    CascadeMux I__2192 (
            .O(N__15410),
            .I(N__15407));
    InMux I__2191 (
            .O(N__15407),
            .I(N__15404));
    LocalMux I__2190 (
            .O(N__15404),
            .I(N__15401));
    Odrv4 I__2189 (
            .O(N__15401),
            .I(\eeprom.n3584 ));
    InMux I__2188 (
            .O(N__15398),
            .I(\eeprom.n4206 ));
    InMux I__2187 (
            .O(N__15395),
            .I(\eeprom.n4229 ));
    InMux I__2186 (
            .O(N__15392),
            .I(\eeprom.n4230 ));
    InMux I__2185 (
            .O(N__15389),
            .I(\eeprom.n4231 ));
    InMux I__2184 (
            .O(N__15386),
            .I(\eeprom.n4232 ));
    InMux I__2183 (
            .O(N__15383),
            .I(\eeprom.n4233 ));
    InMux I__2182 (
            .O(N__15380),
            .I(N__15377));
    LocalMux I__2181 (
            .O(N__15377),
            .I(\eeprom.n5547 ));
    CascadeMux I__2180 (
            .O(N__15374),
            .I(N__15371));
    InMux I__2179 (
            .O(N__15371),
            .I(N__15368));
    LocalMux I__2178 (
            .O(N__15368),
            .I(\eeprom.n5362 ));
    InMux I__2177 (
            .O(N__15365),
            .I(\eeprom.n4234 ));
    InMux I__2176 (
            .O(N__15362),
            .I(N__15359));
    LocalMux I__2175 (
            .O(N__15359),
            .I(\eeprom.n5550 ));
    CascadeMux I__2174 (
            .O(N__15356),
            .I(N__15353));
    InMux I__2173 (
            .O(N__15353),
            .I(N__15350));
    LocalMux I__2172 (
            .O(N__15350),
            .I(\eeprom.n3717 ));
    InMux I__2171 (
            .O(N__15347),
            .I(bfn_20_18_0_));
    InMux I__2170 (
            .O(N__15344),
            .I(\eeprom.n4236 ));
    InMux I__2169 (
            .O(N__15341),
            .I(N__15338));
    LocalMux I__2168 (
            .O(N__15338),
            .I(\eeprom.n5556 ));
    CascadeMux I__2167 (
            .O(N__15335),
            .I(N__15332));
    InMux I__2166 (
            .O(N__15332),
            .I(N__15329));
    LocalMux I__2165 (
            .O(N__15329),
            .I(\eeprom.n3715 ));
    InMux I__2164 (
            .O(N__15326),
            .I(\eeprom.n4237 ));
    CascadeMux I__2163 (
            .O(N__15323),
            .I(N__15320));
    InMux I__2162 (
            .O(N__15320),
            .I(N__15316));
    CascadeMux I__2161 (
            .O(N__15319),
            .I(N__15313));
    LocalMux I__2160 (
            .O(N__15316),
            .I(N__15309));
    InMux I__2159 (
            .O(N__15313),
            .I(N__15306));
    InMux I__2158 (
            .O(N__15312),
            .I(N__15303));
    Span4Mux_h I__2157 (
            .O(N__15309),
            .I(N__15300));
    LocalMux I__2156 (
            .O(N__15306),
            .I(N__15295));
    LocalMux I__2155 (
            .O(N__15303),
            .I(N__15295));
    Odrv4 I__2154 (
            .O(N__15300),
            .I(\eeprom.n3105 ));
    Odrv12 I__2153 (
            .O(N__15295),
            .I(\eeprom.n3105 ));
    InMux I__2152 (
            .O(N__15290),
            .I(N__15287));
    LocalMux I__2151 (
            .O(N__15287),
            .I(N__15284));
    Sp12to4 I__2150 (
            .O(N__15284),
            .I(N__15281));
    Odrv12 I__2149 (
            .O(N__15281),
            .I(\eeprom.n3172 ));
    InMux I__2148 (
            .O(N__15278),
            .I(\eeprom.n4136 ));
    InMux I__2147 (
            .O(N__15275),
            .I(N__15272));
    LocalMux I__2146 (
            .O(N__15272),
            .I(N__15267));
    InMux I__2145 (
            .O(N__15271),
            .I(N__15264));
    InMux I__2144 (
            .O(N__15270),
            .I(N__15261));
    Span4Mux_h I__2143 (
            .O(N__15267),
            .I(N__15258));
    LocalMux I__2142 (
            .O(N__15264),
            .I(N__15255));
    LocalMux I__2141 (
            .O(N__15261),
            .I(N__15252));
    Odrv4 I__2140 (
            .O(N__15258),
            .I(\eeprom.n3104 ));
    Odrv4 I__2139 (
            .O(N__15255),
            .I(\eeprom.n3104 ));
    Odrv12 I__2138 (
            .O(N__15252),
            .I(\eeprom.n3104 ));
    InMux I__2137 (
            .O(N__15245),
            .I(N__15242));
    LocalMux I__2136 (
            .O(N__15242),
            .I(N__15239));
    Span4Mux_v I__2135 (
            .O(N__15239),
            .I(N__15236));
    Odrv4 I__2134 (
            .O(N__15236),
            .I(\eeprom.n3171 ));
    InMux I__2133 (
            .O(N__15233),
            .I(\eeprom.n4137 ));
    CascadeMux I__2132 (
            .O(N__15230),
            .I(N__15227));
    InMux I__2131 (
            .O(N__15227),
            .I(N__15222));
    InMux I__2130 (
            .O(N__15226),
            .I(N__15219));
    InMux I__2129 (
            .O(N__15225),
            .I(N__15216));
    LocalMux I__2128 (
            .O(N__15222),
            .I(N__15211));
    LocalMux I__2127 (
            .O(N__15219),
            .I(N__15211));
    LocalMux I__2126 (
            .O(N__15216),
            .I(\eeprom.n3103 ));
    Odrv12 I__2125 (
            .O(N__15211),
            .I(\eeprom.n3103 ));
    InMux I__2124 (
            .O(N__15206),
            .I(N__15203));
    LocalMux I__2123 (
            .O(N__15203),
            .I(N__15200));
    Span4Mux_v I__2122 (
            .O(N__15200),
            .I(N__15197));
    Odrv4 I__2121 (
            .O(N__15197),
            .I(\eeprom.n3170 ));
    InMux I__2120 (
            .O(N__15194),
            .I(bfn_19_32_0_));
    InMux I__2119 (
            .O(N__15191),
            .I(N__15188));
    LocalMux I__2118 (
            .O(N__15188),
            .I(N__15185));
    Span4Mux_s2_v I__2117 (
            .O(N__15185),
            .I(N__15180));
    InMux I__2116 (
            .O(N__15184),
            .I(N__15175));
    InMux I__2115 (
            .O(N__15183),
            .I(N__15175));
    Odrv4 I__2114 (
            .O(N__15180),
            .I(\eeprom.n3102 ));
    LocalMux I__2113 (
            .O(N__15175),
            .I(\eeprom.n3102 ));
    CascadeMux I__2112 (
            .O(N__15170),
            .I(N__15167));
    InMux I__2111 (
            .O(N__15167),
            .I(N__15164));
    LocalMux I__2110 (
            .O(N__15164),
            .I(N__15161));
    Span4Mux_v I__2109 (
            .O(N__15161),
            .I(N__15158));
    Odrv4 I__2108 (
            .O(N__15158),
            .I(\eeprom.n3169 ));
    InMux I__2107 (
            .O(N__15155),
            .I(\eeprom.n4139 ));
    InMux I__2106 (
            .O(N__15152),
            .I(N__15148));
    InMux I__2105 (
            .O(N__15151),
            .I(N__15145));
    LocalMux I__2104 (
            .O(N__15148),
            .I(N__15142));
    LocalMux I__2103 (
            .O(N__15145),
            .I(N__15138));
    Span4Mux_s3_v I__2102 (
            .O(N__15142),
            .I(N__15135));
    InMux I__2101 (
            .O(N__15141),
            .I(N__15132));
    Odrv4 I__2100 (
            .O(N__15138),
            .I(\eeprom.n3101 ));
    Odrv4 I__2099 (
            .O(N__15135),
            .I(\eeprom.n3101 ));
    LocalMux I__2098 (
            .O(N__15132),
            .I(\eeprom.n3101 ));
    CascadeMux I__2097 (
            .O(N__15125),
            .I(N__15122));
    InMux I__2096 (
            .O(N__15122),
            .I(N__15119));
    LocalMux I__2095 (
            .O(N__15119),
            .I(N__15116));
    Span4Mux_h I__2094 (
            .O(N__15116),
            .I(N__15113));
    Span4Mux_v I__2093 (
            .O(N__15113),
            .I(N__15110));
    Odrv4 I__2092 (
            .O(N__15110),
            .I(\eeprom.n3168 ));
    InMux I__2091 (
            .O(N__15107),
            .I(\eeprom.n4140 ));
    CascadeMux I__2090 (
            .O(N__15104),
            .I(N__15101));
    InMux I__2089 (
            .O(N__15101),
            .I(N__15097));
    InMux I__2088 (
            .O(N__15100),
            .I(N__15094));
    LocalMux I__2087 (
            .O(N__15097),
            .I(N__15091));
    LocalMux I__2086 (
            .O(N__15094),
            .I(\eeprom.n3100 ));
    Odrv12 I__2085 (
            .O(N__15091),
            .I(\eeprom.n3100 ));
    InMux I__2084 (
            .O(N__15086),
            .I(\eeprom.n4141 ));
    InMux I__2083 (
            .O(N__15083),
            .I(N__15079));
    InMux I__2082 (
            .O(N__15082),
            .I(N__15076));
    LocalMux I__2081 (
            .O(N__15079),
            .I(N__15073));
    LocalMux I__2080 (
            .O(N__15076),
            .I(N__15070));
    Span4Mux_h I__2079 (
            .O(N__15073),
            .I(N__15067));
    Span4Mux_h I__2078 (
            .O(N__15070),
            .I(N__15064));
    Span4Mux_v I__2077 (
            .O(N__15067),
            .I(N__15061));
    Odrv4 I__2076 (
            .O(N__15064),
            .I(\eeprom.n3199 ));
    Odrv4 I__2075 (
            .O(N__15061),
            .I(\eeprom.n3199 ));
    InMux I__2074 (
            .O(N__15056),
            .I(bfn_20_17_0_));
    InMux I__2073 (
            .O(N__15053),
            .I(\eeprom.n4228 ));
    InMux I__2072 (
            .O(N__15050),
            .I(N__15046));
    InMux I__2071 (
            .O(N__15049),
            .I(N__15043));
    LocalMux I__2070 (
            .O(N__15046),
            .I(N__15040));
    LocalMux I__2069 (
            .O(N__15043),
            .I(\eeprom.n3113 ));
    Odrv4 I__2068 (
            .O(N__15040),
            .I(\eeprom.n3113 ));
    CascadeMux I__2067 (
            .O(N__15035),
            .I(N__15032));
    InMux I__2066 (
            .O(N__15032),
            .I(N__15029));
    LocalMux I__2065 (
            .O(N__15029),
            .I(N__15026));
    Span4Mux_h I__2064 (
            .O(N__15026),
            .I(N__15023));
    Odrv4 I__2063 (
            .O(N__15023),
            .I(\eeprom.n3180 ));
    InMux I__2062 (
            .O(N__15020),
            .I(\eeprom.n4128 ));
    InMux I__2061 (
            .O(N__15017),
            .I(N__15014));
    LocalMux I__2060 (
            .O(N__15014),
            .I(N__15011));
    Span4Mux_v I__2059 (
            .O(N__15011),
            .I(N__15008));
    Odrv4 I__2058 (
            .O(N__15008),
            .I(\eeprom.n3179 ));
    InMux I__2057 (
            .O(N__15005),
            .I(\eeprom.n4129 ));
    InMux I__2056 (
            .O(N__15002),
            .I(N__14999));
    LocalMux I__2055 (
            .O(N__14999),
            .I(N__14994));
    InMux I__2054 (
            .O(N__14998),
            .I(N__14991));
    InMux I__2053 (
            .O(N__14997),
            .I(N__14988));
    Span4Mux_s3_v I__2052 (
            .O(N__14994),
            .I(N__14985));
    LocalMux I__2051 (
            .O(N__14991),
            .I(N__14980));
    LocalMux I__2050 (
            .O(N__14988),
            .I(N__14980));
    Odrv4 I__2049 (
            .O(N__14985),
            .I(\eeprom.n3111 ));
    Odrv4 I__2048 (
            .O(N__14980),
            .I(\eeprom.n3111 ));
    InMux I__2047 (
            .O(N__14975),
            .I(N__14972));
    LocalMux I__2046 (
            .O(N__14972),
            .I(N__14969));
    Span4Mux_v I__2045 (
            .O(N__14969),
            .I(N__14966));
    Odrv4 I__2044 (
            .O(N__14966),
            .I(\eeprom.n3178 ));
    InMux I__2043 (
            .O(N__14963),
            .I(bfn_19_31_0_));
    InMux I__2042 (
            .O(N__14960),
            .I(\eeprom.n4131 ));
    InMux I__2041 (
            .O(N__14957),
            .I(\eeprom.n4132 ));
    CascadeMux I__2040 (
            .O(N__14954),
            .I(N__14951));
    InMux I__2039 (
            .O(N__14951),
            .I(N__14947));
    CascadeMux I__2038 (
            .O(N__14950),
            .I(N__14944));
    LocalMux I__2037 (
            .O(N__14947),
            .I(N__14941));
    InMux I__2036 (
            .O(N__14944),
            .I(N__14938));
    Span4Mux_v I__2035 (
            .O(N__14941),
            .I(N__14935));
    LocalMux I__2034 (
            .O(N__14938),
            .I(\eeprom.n3108 ));
    Odrv4 I__2033 (
            .O(N__14935),
            .I(\eeprom.n3108 ));
    InMux I__2032 (
            .O(N__14930),
            .I(N__14927));
    LocalMux I__2031 (
            .O(N__14927),
            .I(N__14924));
    Span4Mux_v I__2030 (
            .O(N__14924),
            .I(N__14921));
    Odrv4 I__2029 (
            .O(N__14921),
            .I(\eeprom.n3175 ));
    InMux I__2028 (
            .O(N__14918),
            .I(\eeprom.n4133 ));
    CascadeMux I__2027 (
            .O(N__14915),
            .I(N__14911));
    InMux I__2026 (
            .O(N__14914),
            .I(N__14907));
    InMux I__2025 (
            .O(N__14911),
            .I(N__14902));
    InMux I__2024 (
            .O(N__14910),
            .I(N__14902));
    LocalMux I__2023 (
            .O(N__14907),
            .I(N__14899));
    LocalMux I__2022 (
            .O(N__14902),
            .I(N__14896));
    Odrv4 I__2021 (
            .O(N__14899),
            .I(\eeprom.n3107 ));
    Odrv4 I__2020 (
            .O(N__14896),
            .I(\eeprom.n3107 ));
    InMux I__2019 (
            .O(N__14891),
            .I(N__14888));
    LocalMux I__2018 (
            .O(N__14888),
            .I(N__14885));
    Span4Mux_v I__2017 (
            .O(N__14885),
            .I(N__14882));
    Odrv4 I__2016 (
            .O(N__14882),
            .I(\eeprom.n3174 ));
    InMux I__2015 (
            .O(N__14879),
            .I(\eeprom.n4134 ));
    InMux I__2014 (
            .O(N__14876),
            .I(N__14871));
    InMux I__2013 (
            .O(N__14875),
            .I(N__14866));
    InMux I__2012 (
            .O(N__14874),
            .I(N__14866));
    LocalMux I__2011 (
            .O(N__14871),
            .I(N__14863));
    LocalMux I__2010 (
            .O(N__14866),
            .I(N__14860));
    Odrv12 I__2009 (
            .O(N__14863),
            .I(\eeprom.n3106 ));
    Odrv4 I__2008 (
            .O(N__14860),
            .I(\eeprom.n3106 ));
    InMux I__2007 (
            .O(N__14855),
            .I(N__14852));
    LocalMux I__2006 (
            .O(N__14852),
            .I(N__14849));
    Odrv12 I__2005 (
            .O(N__14849),
            .I(\eeprom.n3173 ));
    InMux I__2004 (
            .O(N__14846),
            .I(\eeprom.n4135 ));
    InMux I__2003 (
            .O(N__14843),
            .I(N__14836));
    InMux I__2002 (
            .O(N__14842),
            .I(N__14836));
    InMux I__2001 (
            .O(N__14841),
            .I(N__14833));
    LocalMux I__2000 (
            .O(N__14836),
            .I(\eeprom.n3012 ));
    LocalMux I__1999 (
            .O(N__14833),
            .I(\eeprom.n3012 ));
    InMux I__1998 (
            .O(N__14828),
            .I(N__14824));
    InMux I__1997 (
            .O(N__14827),
            .I(N__14821));
    LocalMux I__1996 (
            .O(N__14824),
            .I(N__14818));
    LocalMux I__1995 (
            .O(N__14821),
            .I(N__14814));
    Span4Mux_h I__1994 (
            .O(N__14818),
            .I(N__14811));
    InMux I__1993 (
            .O(N__14817),
            .I(N__14808));
    Odrv4 I__1992 (
            .O(N__14814),
            .I(\eeprom.n3003 ));
    Odrv4 I__1991 (
            .O(N__14811),
            .I(\eeprom.n3003 ));
    LocalMux I__1990 (
            .O(N__14808),
            .I(\eeprom.n3003 ));
    InMux I__1989 (
            .O(N__14801),
            .I(N__14798));
    LocalMux I__1988 (
            .O(N__14798),
            .I(\eeprom.n3086 ));
    InMux I__1987 (
            .O(N__14795),
            .I(N__14792));
    LocalMux I__1986 (
            .O(N__14792),
            .I(N__14789));
    Span4Mux_h I__1985 (
            .O(N__14789),
            .I(N__14786));
    Span4Mux_h I__1984 (
            .O(N__14786),
            .I(N__14783));
    Odrv4 I__1983 (
            .O(N__14783),
            .I(\eeprom.n3186 ));
    InMux I__1982 (
            .O(N__14780),
            .I(bfn_19_30_0_));
    InMux I__1981 (
            .O(N__14777),
            .I(\eeprom.n4123 ));
    CascadeMux I__1980 (
            .O(N__14774),
            .I(N__14770));
    CascadeMux I__1979 (
            .O(N__14773),
            .I(N__14767));
    InMux I__1978 (
            .O(N__14770),
            .I(N__14764));
    InMux I__1977 (
            .O(N__14767),
            .I(N__14760));
    LocalMux I__1976 (
            .O(N__14764),
            .I(N__14757));
    InMux I__1975 (
            .O(N__14763),
            .I(N__14754));
    LocalMux I__1974 (
            .O(N__14760),
            .I(N__14751));
    Odrv4 I__1973 (
            .O(N__14757),
            .I(\eeprom.n3117 ));
    LocalMux I__1972 (
            .O(N__14754),
            .I(\eeprom.n3117 ));
    Odrv4 I__1971 (
            .O(N__14751),
            .I(\eeprom.n3117 ));
    InMux I__1970 (
            .O(N__14744),
            .I(N__14741));
    LocalMux I__1969 (
            .O(N__14741),
            .I(N__14738));
    Odrv12 I__1968 (
            .O(N__14738),
            .I(\eeprom.n3184 ));
    InMux I__1967 (
            .O(N__14735),
            .I(\eeprom.n4124 ));
    InMux I__1966 (
            .O(N__14732),
            .I(\eeprom.n4125 ));
    InMux I__1965 (
            .O(N__14729),
            .I(\eeprom.n4126 ));
    InMux I__1964 (
            .O(N__14726),
            .I(\eeprom.n4127 ));
    CascadeMux I__1963 (
            .O(N__14723),
            .I(N__14720));
    InMux I__1962 (
            .O(N__14720),
            .I(N__14717));
    LocalMux I__1961 (
            .O(N__14717),
            .I(N__14713));
    InMux I__1960 (
            .O(N__14716),
            .I(N__14710));
    Odrv4 I__1959 (
            .O(N__14713),
            .I(\eeprom.n3007 ));
    LocalMux I__1958 (
            .O(N__14710),
            .I(\eeprom.n3007 ));
    InMux I__1957 (
            .O(N__14705),
            .I(N__14702));
    LocalMux I__1956 (
            .O(N__14702),
            .I(N__14699));
    Span4Mux_h I__1955 (
            .O(N__14699),
            .I(N__14696));
    Odrv4 I__1954 (
            .O(N__14696),
            .I(\eeprom.n3074 ));
    CascadeMux I__1953 (
            .O(N__14693),
            .I(\eeprom.n3007_cascade_ ));
    CascadeMux I__1952 (
            .O(N__14690),
            .I(N__14686));
    InMux I__1951 (
            .O(N__14689),
            .I(N__14683));
    InMux I__1950 (
            .O(N__14686),
            .I(N__14680));
    LocalMux I__1949 (
            .O(N__14683),
            .I(N__14677));
    LocalMux I__1948 (
            .O(N__14680),
            .I(\eeprom.n3006 ));
    Odrv4 I__1947 (
            .O(N__14677),
            .I(\eeprom.n3006 ));
    InMux I__1946 (
            .O(N__14672),
            .I(N__14669));
    LocalMux I__1945 (
            .O(N__14669),
            .I(\eeprom.n21_adj_336 ));
    CascadeMux I__1944 (
            .O(N__14666),
            .I(\eeprom.n3006_cascade_ ));
    InMux I__1943 (
            .O(N__14663),
            .I(N__14660));
    LocalMux I__1942 (
            .O(N__14660),
            .I(N__14657));
    Odrv4 I__1941 (
            .O(N__14657),
            .I(\eeprom.n18_adj_335 ));
    InMux I__1940 (
            .O(N__14654),
            .I(N__14651));
    LocalMux I__1939 (
            .O(N__14651),
            .I(\eeprom.n24_adj_340 ));
    CascadeMux I__1938 (
            .O(N__14648),
            .I(N__14645));
    InMux I__1937 (
            .O(N__14645),
            .I(N__14640));
    InMux I__1936 (
            .O(N__14644),
            .I(N__14637));
    InMux I__1935 (
            .O(N__14643),
            .I(N__14634));
    LocalMux I__1934 (
            .O(N__14640),
            .I(N__14631));
    LocalMux I__1933 (
            .O(N__14637),
            .I(N__14626));
    LocalMux I__1932 (
            .O(N__14634),
            .I(N__14626));
    Odrv4 I__1931 (
            .O(N__14631),
            .I(\eeprom.n3008 ));
    Odrv4 I__1930 (
            .O(N__14626),
            .I(\eeprom.n3008 ));
    InMux I__1929 (
            .O(N__14621),
            .I(N__14617));
    CascadeMux I__1928 (
            .O(N__14620),
            .I(N__14614));
    LocalMux I__1927 (
            .O(N__14617),
            .I(N__14611));
    InMux I__1926 (
            .O(N__14614),
            .I(N__14608));
    Odrv4 I__1925 (
            .O(N__14611),
            .I(\eeprom.n3005 ));
    LocalMux I__1924 (
            .O(N__14608),
            .I(\eeprom.n3005 ));
    CascadeMux I__1923 (
            .O(N__14603),
            .I(\eeprom.n3005_cascade_ ));
    InMux I__1922 (
            .O(N__14600),
            .I(N__14597));
    LocalMux I__1921 (
            .O(N__14597),
            .I(N__14594));
    Span4Mux_h I__1920 (
            .O(N__14594),
            .I(N__14591));
    Odrv4 I__1919 (
            .O(N__14591),
            .I(\eeprom.n3072 ));
    InMux I__1918 (
            .O(N__14588),
            .I(N__14585));
    LocalMux I__1917 (
            .O(N__14585),
            .I(\eeprom.n3082 ));
    CascadeMux I__1916 (
            .O(N__14582),
            .I(N__14577));
    InMux I__1915 (
            .O(N__14581),
            .I(N__14572));
    InMux I__1914 (
            .O(N__14580),
            .I(N__14572));
    InMux I__1913 (
            .O(N__14577),
            .I(N__14569));
    LocalMux I__1912 (
            .O(N__14572),
            .I(\eeprom.n3010 ));
    LocalMux I__1911 (
            .O(N__14569),
            .I(\eeprom.n3010 ));
    InMux I__1910 (
            .O(N__14564),
            .I(N__14561));
    LocalMux I__1909 (
            .O(N__14561),
            .I(N__14557));
    InMux I__1908 (
            .O(N__14560),
            .I(N__14554));
    Span12Mux_s6_v I__1907 (
            .O(N__14557),
            .I(N__14551));
    LocalMux I__1906 (
            .O(N__14554),
            .I(\eeprom.n3002 ));
    Odrv12 I__1905 (
            .O(N__14551),
            .I(\eeprom.n3002 ));
    CascadeMux I__1904 (
            .O(N__14546),
            .I(\eeprom.n3002_cascade_ ));
    CascadeMux I__1903 (
            .O(N__14543),
            .I(N__14540));
    InMux I__1902 (
            .O(N__14540),
            .I(N__14537));
    LocalMux I__1901 (
            .O(N__14537),
            .I(N__14534));
    Span4Mux_h I__1900 (
            .O(N__14534),
            .I(N__14531));
    Odrv4 I__1899 (
            .O(N__14531),
            .I(\eeprom.n20_adj_337 ));
    CascadeMux I__1898 (
            .O(N__14528),
            .I(N__14525));
    InMux I__1897 (
            .O(N__14525),
            .I(N__14522));
    LocalMux I__1896 (
            .O(N__14522),
            .I(N__14519));
    Span4Mux_h I__1895 (
            .O(N__14519),
            .I(N__14516));
    Odrv4 I__1894 (
            .O(N__14516),
            .I(\eeprom.n3078 ));
    InMux I__1893 (
            .O(N__14513),
            .I(N__14509));
    InMux I__1892 (
            .O(N__14512),
            .I(N__14505));
    LocalMux I__1891 (
            .O(N__14509),
            .I(N__14502));
    InMux I__1890 (
            .O(N__14508),
            .I(N__14499));
    LocalMux I__1889 (
            .O(N__14505),
            .I(\eeprom.n3016 ));
    Odrv4 I__1888 (
            .O(N__14502),
            .I(\eeprom.n3016 ));
    LocalMux I__1887 (
            .O(N__14499),
            .I(\eeprom.n3016 ));
    CascadeMux I__1886 (
            .O(N__14492),
            .I(N__14488));
    InMux I__1885 (
            .O(N__14491),
            .I(N__14484));
    InMux I__1884 (
            .O(N__14488),
            .I(N__14481));
    InMux I__1883 (
            .O(N__14487),
            .I(N__14478));
    LocalMux I__1882 (
            .O(N__14484),
            .I(N__14475));
    LocalMux I__1881 (
            .O(N__14481),
            .I(\eeprom.n3018 ));
    LocalMux I__1880 (
            .O(N__14478),
            .I(\eeprom.n3018 ));
    Odrv4 I__1879 (
            .O(N__14475),
            .I(\eeprom.n3018 ));
    CascadeMux I__1878 (
            .O(N__14468),
            .I(\eeprom.n2914_cascade_ ));
    InMux I__1877 (
            .O(N__14465),
            .I(N__14462));
    LocalMux I__1876 (
            .O(N__14462),
            .I(N__14459));
    Odrv4 I__1875 (
            .O(N__14459),
            .I(\eeprom.n3073 ));
    CascadeMux I__1874 (
            .O(N__14456),
            .I(N__14453));
    InMux I__1873 (
            .O(N__14453),
            .I(N__14449));
    CascadeMux I__1872 (
            .O(N__14452),
            .I(N__14446));
    LocalMux I__1871 (
            .O(N__14449),
            .I(N__14443));
    InMux I__1870 (
            .O(N__14446),
            .I(N__14439));
    Span4Mux_h I__1869 (
            .O(N__14443),
            .I(N__14436));
    InMux I__1868 (
            .O(N__14442),
            .I(N__14433));
    LocalMux I__1867 (
            .O(N__14439),
            .I(\eeprom.n3014 ));
    Odrv4 I__1866 (
            .O(N__14436),
            .I(\eeprom.n3014 ));
    LocalMux I__1865 (
            .O(N__14433),
            .I(\eeprom.n3014 ));
    InMux I__1864 (
            .O(N__14426),
            .I(N__14423));
    LocalMux I__1863 (
            .O(N__14423),
            .I(N__14419));
    InMux I__1862 (
            .O(N__14422),
            .I(N__14416));
    Span4Mux_h I__1861 (
            .O(N__14419),
            .I(N__14413));
    LocalMux I__1860 (
            .O(N__14416),
            .I(\eeprom.n3205 ));
    Odrv4 I__1859 (
            .O(N__14413),
            .I(\eeprom.n3205 ));
    InMux I__1858 (
            .O(N__14408),
            .I(N__14405));
    LocalMux I__1857 (
            .O(N__14405),
            .I(N__14402));
    Span4Mux_h I__1856 (
            .O(N__14402),
            .I(N__14399));
    Odrv4 I__1855 (
            .O(N__14399),
            .I(\eeprom.n3272 ));
    CascadeMux I__1854 (
            .O(N__14396),
            .I(\eeprom.n3205_cascade_ ));
    InMux I__1853 (
            .O(N__14393),
            .I(N__14389));
    InMux I__1852 (
            .O(N__14392),
            .I(N__14386));
    LocalMux I__1851 (
            .O(N__14389),
            .I(N__14383));
    LocalMux I__1850 (
            .O(N__14386),
            .I(\eeprom.n3204 ));
    Odrv4 I__1849 (
            .O(N__14383),
            .I(\eeprom.n3204 ));
    InMux I__1848 (
            .O(N__14378),
            .I(N__14375));
    LocalMux I__1847 (
            .O(N__14375),
            .I(N__14372));
    Span4Mux_h I__1846 (
            .O(N__14372),
            .I(N__14369));
    Odrv4 I__1845 (
            .O(N__14369),
            .I(\eeprom.n3271 ));
    CascadeMux I__1844 (
            .O(N__14366),
            .I(N__14363));
    InMux I__1843 (
            .O(N__14363),
            .I(N__14360));
    LocalMux I__1842 (
            .O(N__14360),
            .I(N__14355));
    InMux I__1841 (
            .O(N__14359),
            .I(N__14350));
    InMux I__1840 (
            .O(N__14358),
            .I(N__14350));
    Span4Mux_h I__1839 (
            .O(N__14355),
            .I(N__14347));
    LocalMux I__1838 (
            .O(N__14350),
            .I(\eeprom.n3207 ));
    Odrv4 I__1837 (
            .O(N__14347),
            .I(\eeprom.n3207 ));
    CascadeMux I__1836 (
            .O(N__14342),
            .I(N__14339));
    InMux I__1835 (
            .O(N__14339),
            .I(N__14336));
    LocalMux I__1834 (
            .O(N__14336),
            .I(N__14332));
    InMux I__1833 (
            .O(N__14335),
            .I(N__14329));
    Span4Mux_v I__1832 (
            .O(N__14332),
            .I(N__14326));
    LocalMux I__1831 (
            .O(N__14329),
            .I(\eeprom.n3017 ));
    Odrv4 I__1830 (
            .O(N__14326),
            .I(\eeprom.n3017 ));
    CascadeMux I__1829 (
            .O(N__14321),
            .I(\eeprom.n3017_cascade_ ));
    CascadeMux I__1828 (
            .O(N__14318),
            .I(\eeprom.n5147_cascade_ ));
    InMux I__1827 (
            .O(N__14315),
            .I(N__14311));
    CascadeMux I__1826 (
            .O(N__14314),
            .I(N__14308));
    LocalMux I__1825 (
            .O(N__14311),
            .I(N__14305));
    InMux I__1824 (
            .O(N__14308),
            .I(N__14301));
    Span4Mux_v I__1823 (
            .O(N__14305),
            .I(N__14298));
    InMux I__1822 (
            .O(N__14304),
            .I(N__14295));
    LocalMux I__1821 (
            .O(N__14301),
            .I(\eeprom.n3009 ));
    Odrv4 I__1820 (
            .O(N__14298),
            .I(\eeprom.n3009 ));
    LocalMux I__1819 (
            .O(N__14295),
            .I(\eeprom.n3009 ));
    InMux I__1818 (
            .O(N__14288),
            .I(N__14284));
    InMux I__1817 (
            .O(N__14287),
            .I(N__14281));
    LocalMux I__1816 (
            .O(N__14284),
            .I(N__14278));
    LocalMux I__1815 (
            .O(N__14281),
            .I(\eeprom.n3206 ));
    Odrv4 I__1814 (
            .O(N__14278),
            .I(\eeprom.n3206 ));
    CascadeMux I__1813 (
            .O(N__14273),
            .I(\eeprom.n20_adj_301_cascade_ ));
    InMux I__1812 (
            .O(N__14270),
            .I(N__14267));
    LocalMux I__1811 (
            .O(N__14267),
            .I(\eeprom.n16_adj_303 ));
    CascadeMux I__1810 (
            .O(N__14264),
            .I(N__14261));
    InMux I__1809 (
            .O(N__14261),
            .I(N__14256));
    InMux I__1808 (
            .O(N__14260),
            .I(N__14253));
    InMux I__1807 (
            .O(N__14259),
            .I(N__14250));
    LocalMux I__1806 (
            .O(N__14256),
            .I(N__14245));
    LocalMux I__1805 (
            .O(N__14253),
            .I(N__14245));
    LocalMux I__1804 (
            .O(N__14250),
            .I(\eeprom.n3212 ));
    Odrv4 I__1803 (
            .O(N__14245),
            .I(\eeprom.n3212 ));
    CascadeMux I__1802 (
            .O(N__14240),
            .I(\eeprom.n28_adj_305_cascade_ ));
    InMux I__1801 (
            .O(N__14237),
            .I(N__14234));
    LocalMux I__1800 (
            .O(N__14234),
            .I(\eeprom.n24_adj_304 ));
    CascadeMux I__1799 (
            .O(N__14231),
            .I(\eeprom.n3232_cascade_ ));
    InMux I__1798 (
            .O(N__14228),
            .I(N__14225));
    LocalMux I__1797 (
            .O(N__14225),
            .I(N__14222));
    Span4Mux_h I__1796 (
            .O(N__14222),
            .I(N__14219));
    Odrv4 I__1795 (
            .O(N__14219),
            .I(\eeprom.n3274 ));
    CascadeMux I__1794 (
            .O(N__14216),
            .I(N__14213));
    InMux I__1793 (
            .O(N__14213),
            .I(N__14210));
    LocalMux I__1792 (
            .O(N__14210),
            .I(N__14206));
    InMux I__1791 (
            .O(N__14209),
            .I(N__14203));
    Span4Mux_v I__1790 (
            .O(N__14206),
            .I(N__14200));
    LocalMux I__1789 (
            .O(N__14203),
            .I(\eeprom.n3306 ));
    Odrv4 I__1788 (
            .O(N__14200),
            .I(\eeprom.n3306 ));
    InMux I__1787 (
            .O(N__14195),
            .I(N__14191));
    CascadeMux I__1786 (
            .O(N__14194),
            .I(N__14188));
    LocalMux I__1785 (
            .O(N__14191),
            .I(N__14184));
    InMux I__1784 (
            .O(N__14188),
            .I(N__14181));
    InMux I__1783 (
            .O(N__14187),
            .I(N__14178));
    Odrv4 I__1782 (
            .O(N__14184),
            .I(\eeprom.n3305 ));
    LocalMux I__1781 (
            .O(N__14181),
            .I(\eeprom.n3305 ));
    LocalMux I__1780 (
            .O(N__14178),
            .I(\eeprom.n3305 ));
    CascadeMux I__1779 (
            .O(N__14171),
            .I(\eeprom.n3306_cascade_ ));
    CascadeMux I__1778 (
            .O(N__14168),
            .I(N__14165));
    InMux I__1777 (
            .O(N__14165),
            .I(N__14161));
    CascadeMux I__1776 (
            .O(N__14164),
            .I(N__14158));
    LocalMux I__1775 (
            .O(N__14161),
            .I(N__14154));
    InMux I__1774 (
            .O(N__14158),
            .I(N__14151));
    InMux I__1773 (
            .O(N__14157),
            .I(N__14148));
    Odrv4 I__1772 (
            .O(N__14154),
            .I(\eeprom.n3308 ));
    LocalMux I__1771 (
            .O(N__14151),
            .I(\eeprom.n3308 ));
    LocalMux I__1770 (
            .O(N__14148),
            .I(\eeprom.n3308 ));
    InMux I__1769 (
            .O(N__14141),
            .I(N__14138));
    LocalMux I__1768 (
            .O(N__14138),
            .I(\eeprom.n27 ));
    InMux I__1767 (
            .O(N__14135),
            .I(N__14132));
    LocalMux I__1766 (
            .O(N__14132),
            .I(N__14129));
    Odrv4 I__1765 (
            .O(N__14129),
            .I(\eeprom.n5309 ));
    CascadeMux I__1764 (
            .O(N__14126),
            .I(\eeprom.n18_adj_260_cascade_ ));
    InMux I__1763 (
            .O(N__14123),
            .I(N__14120));
    LocalMux I__1762 (
            .O(N__14120),
            .I(\eeprom.n24 ));
    InMux I__1761 (
            .O(N__14117),
            .I(N__14114));
    LocalMux I__1760 (
            .O(N__14114),
            .I(\eeprom.n22 ));
    CascadeMux I__1759 (
            .O(N__14111),
            .I(\eeprom.n26_adj_262_cascade_ ));
    CascadeMux I__1758 (
            .O(N__14108),
            .I(\eeprom.n3133_cascade_ ));
    CascadeMux I__1757 (
            .O(N__14105),
            .I(N__14102));
    InMux I__1756 (
            .O(N__14102),
            .I(N__14099));
    LocalMux I__1755 (
            .O(N__14099),
            .I(N__14096));
    Span4Mux_h I__1754 (
            .O(N__14096),
            .I(N__14093));
    Odrv4 I__1753 (
            .O(N__14093),
            .I(\eeprom.n3373 ));
    CascadeMux I__1752 (
            .O(N__14090),
            .I(N__14087));
    InMux I__1751 (
            .O(N__14087),
            .I(N__14084));
    LocalMux I__1750 (
            .O(N__14084),
            .I(N__14081));
    Span4Mux_h I__1749 (
            .O(N__14081),
            .I(N__14078));
    Odrv4 I__1748 (
            .O(N__14078),
            .I(\eeprom.n3369 ));
    InMux I__1747 (
            .O(N__14075),
            .I(N__14071));
    InMux I__1746 (
            .O(N__14074),
            .I(N__14068));
    LocalMux I__1745 (
            .O(N__14071),
            .I(N__14065));
    LocalMux I__1744 (
            .O(N__14068),
            .I(N__14062));
    Odrv4 I__1743 (
            .O(N__14065),
            .I(\eeprom.n3401 ));
    Odrv4 I__1742 (
            .O(N__14062),
            .I(\eeprom.n3401 ));
    CascadeMux I__1741 (
            .O(N__14057),
            .I(N__14053));
    InMux I__1740 (
            .O(N__14056),
            .I(N__14049));
    InMux I__1739 (
            .O(N__14053),
            .I(N__14046));
    InMux I__1738 (
            .O(N__14052),
            .I(N__14043));
    LocalMux I__1737 (
            .O(N__14049),
            .I(\eeprom.n3400 ));
    LocalMux I__1736 (
            .O(N__14046),
            .I(\eeprom.n3400 ));
    LocalMux I__1735 (
            .O(N__14043),
            .I(\eeprom.n3400 ));
    CascadeMux I__1734 (
            .O(N__14036),
            .I(N__14032));
    InMux I__1733 (
            .O(N__14035),
            .I(N__14028));
    InMux I__1732 (
            .O(N__14032),
            .I(N__14025));
    InMux I__1731 (
            .O(N__14031),
            .I(N__14022));
    LocalMux I__1730 (
            .O(N__14028),
            .I(\eeprom.n3399 ));
    LocalMux I__1729 (
            .O(N__14025),
            .I(\eeprom.n3399 ));
    LocalMux I__1728 (
            .O(N__14022),
            .I(\eeprom.n3399 ));
    CascadeMux I__1727 (
            .O(N__14015),
            .I(\eeprom.n3401_cascade_ ));
    InMux I__1726 (
            .O(N__14012),
            .I(N__14009));
    LocalMux I__1725 (
            .O(N__14009),
            .I(\eeprom.n27_adj_263 ));
    CascadeMux I__1724 (
            .O(N__14006),
            .I(N__14003));
    InMux I__1723 (
            .O(N__14003),
            .I(N__13998));
    InMux I__1722 (
            .O(N__14002),
            .I(N__13993));
    InMux I__1721 (
            .O(N__14001),
            .I(N__13993));
    LocalMux I__1720 (
            .O(N__13998),
            .I(\eeprom.n3402 ));
    LocalMux I__1719 (
            .O(N__13993),
            .I(\eeprom.n3402 ));
    CascadeMux I__1718 (
            .O(N__13988),
            .I(N__13985));
    InMux I__1717 (
            .O(N__13985),
            .I(N__13982));
    LocalMux I__1716 (
            .O(N__13982),
            .I(N__13979));
    Odrv4 I__1715 (
            .O(N__13979),
            .I(\eeprom.n3469 ));
    CascadeMux I__1714 (
            .O(N__13976),
            .I(N__13972));
    CascadeMux I__1713 (
            .O(N__13975),
            .I(N__13969));
    InMux I__1712 (
            .O(N__13972),
            .I(N__13965));
    InMux I__1711 (
            .O(N__13969),
            .I(N__13962));
    InMux I__1710 (
            .O(N__13968),
            .I(N__13959));
    LocalMux I__1709 (
            .O(N__13965),
            .I(\eeprom.n3307 ));
    LocalMux I__1708 (
            .O(N__13962),
            .I(\eeprom.n3307 ));
    LocalMux I__1707 (
            .O(N__13959),
            .I(\eeprom.n3307 ));
    InMux I__1706 (
            .O(N__13952),
            .I(N__13947));
    CascadeMux I__1705 (
            .O(N__13951),
            .I(N__13944));
    InMux I__1704 (
            .O(N__13950),
            .I(N__13941));
    LocalMux I__1703 (
            .O(N__13947),
            .I(N__13938));
    InMux I__1702 (
            .O(N__13944),
            .I(N__13935));
    LocalMux I__1701 (
            .O(N__13941),
            .I(N__13932));
    Odrv4 I__1700 (
            .O(N__13938),
            .I(\eeprom.n3311 ));
    LocalMux I__1699 (
            .O(N__13935),
            .I(\eeprom.n3311 ));
    Odrv4 I__1698 (
            .O(N__13932),
            .I(\eeprom.n3311 ));
    CascadeMux I__1697 (
            .O(N__13925),
            .I(N__13920));
    CascadeMux I__1696 (
            .O(N__13924),
            .I(N__13917));
    CascadeMux I__1695 (
            .O(N__13923),
            .I(N__13914));
    InMux I__1694 (
            .O(N__13920),
            .I(N__13911));
    InMux I__1693 (
            .O(N__13917),
            .I(N__13908));
    InMux I__1692 (
            .O(N__13914),
            .I(N__13905));
    LocalMux I__1691 (
            .O(N__13911),
            .I(\eeprom.n3312 ));
    LocalMux I__1690 (
            .O(N__13908),
            .I(\eeprom.n3312 ));
    LocalMux I__1689 (
            .O(N__13905),
            .I(\eeprom.n3312 ));
    InMux I__1688 (
            .O(N__13898),
            .I(N__13894));
    InMux I__1687 (
            .O(N__13897),
            .I(N__13891));
    LocalMux I__1686 (
            .O(N__13894),
            .I(N__13887));
    LocalMux I__1685 (
            .O(N__13891),
            .I(N__13884));
    InMux I__1684 (
            .O(N__13890),
            .I(N__13881));
    Span4Mux_v I__1683 (
            .O(N__13887),
            .I(N__13876));
    Span4Mux_h I__1682 (
            .O(N__13884),
            .I(N__13876));
    LocalMux I__1681 (
            .O(N__13881),
            .I(\eeprom.n3309 ));
    Odrv4 I__1680 (
            .O(N__13876),
            .I(\eeprom.n3309 ));
    CascadeMux I__1679 (
            .O(N__13871),
            .I(\eeprom.n28_cascade_ ));
    InMux I__1678 (
            .O(N__13868),
            .I(N__13865));
    LocalMux I__1677 (
            .O(N__13865),
            .I(\eeprom.n25 ));
    InMux I__1676 (
            .O(N__13862),
            .I(N__13859));
    LocalMux I__1675 (
            .O(N__13859),
            .I(N__13856));
    Span4Mux_v I__1674 (
            .O(N__13856),
            .I(N__13853));
    Odrv4 I__1673 (
            .O(N__13853),
            .I(\eeprom.n3385 ));
    CascadeMux I__1672 (
            .O(N__13850),
            .I(\eeprom.n3331_cascade_ ));
    CascadeMux I__1671 (
            .O(N__13847),
            .I(N__13844));
    InMux I__1670 (
            .O(N__13844),
            .I(N__13841));
    LocalMux I__1669 (
            .O(N__13841),
            .I(N__13838));
    Span4Mux_v I__1668 (
            .O(N__13838),
            .I(N__13835));
    Odrv4 I__1667 (
            .O(N__13835),
            .I(\eeprom.n3281 ));
    CascadeMux I__1666 (
            .O(N__13832),
            .I(N__13829));
    InMux I__1665 (
            .O(N__13829),
            .I(N__13826));
    LocalMux I__1664 (
            .O(N__13826),
            .I(N__13823));
    Odrv4 I__1663 (
            .O(N__13823),
            .I(\eeprom.n3485 ));
    CascadeMux I__1662 (
            .O(N__13820),
            .I(N__13815));
    InMux I__1661 (
            .O(N__13819),
            .I(N__13812));
    InMux I__1660 (
            .O(N__13818),
            .I(N__13809));
    InMux I__1659 (
            .O(N__13815),
            .I(N__13806));
    LocalMux I__1658 (
            .O(N__13812),
            .I(\eeprom.n3398 ));
    LocalMux I__1657 (
            .O(N__13809),
            .I(\eeprom.n3398 ));
    LocalMux I__1656 (
            .O(N__13806),
            .I(\eeprom.n3398 ));
    InMux I__1655 (
            .O(N__13799),
            .I(N__13795));
    InMux I__1654 (
            .O(N__13798),
            .I(N__13792));
    LocalMux I__1653 (
            .O(N__13795),
            .I(N__13789));
    LocalMux I__1652 (
            .O(N__13792),
            .I(N__13784));
    Span4Mux_h I__1651 (
            .O(N__13789),
            .I(N__13784));
    Odrv4 I__1650 (
            .O(N__13784),
            .I(\eeprom.n3397 ));
    CascadeMux I__1649 (
            .O(N__13781),
            .I(N__13776));
    InMux I__1648 (
            .O(N__13780),
            .I(N__13773));
    InMux I__1647 (
            .O(N__13779),
            .I(N__13770));
    InMux I__1646 (
            .O(N__13776),
            .I(N__13767));
    LocalMux I__1645 (
            .O(N__13773),
            .I(\eeprom.n3408 ));
    LocalMux I__1644 (
            .O(N__13770),
            .I(\eeprom.n3408 ));
    LocalMux I__1643 (
            .O(N__13767),
            .I(\eeprom.n3408 ));
    InMux I__1642 (
            .O(N__13760),
            .I(N__13756));
    CascadeMux I__1641 (
            .O(N__13759),
            .I(N__13752));
    LocalMux I__1640 (
            .O(N__13756),
            .I(N__13749));
    InMux I__1639 (
            .O(N__13755),
            .I(N__13746));
    InMux I__1638 (
            .O(N__13752),
            .I(N__13743));
    Odrv4 I__1637 (
            .O(N__13749),
            .I(\eeprom.n3411 ));
    LocalMux I__1636 (
            .O(N__13746),
            .I(\eeprom.n3411 ));
    LocalMux I__1635 (
            .O(N__13743),
            .I(\eeprom.n3411 ));
    CascadeMux I__1634 (
            .O(N__13736),
            .I(\eeprom.n18_cascade_ ));
    InMux I__1633 (
            .O(N__13733),
            .I(N__13730));
    LocalMux I__1632 (
            .O(N__13730),
            .I(\eeprom.n29 ));
    CascadeMux I__1631 (
            .O(N__13727),
            .I(\eeprom.n30_cascade_ ));
    CascadeMux I__1630 (
            .O(N__13724),
            .I(\eeprom.n3430_cascade_ ));
    InMux I__1629 (
            .O(N__13721),
            .I(N__13718));
    LocalMux I__1628 (
            .O(N__13718),
            .I(N__13715));
    Span4Mux_h I__1627 (
            .O(N__13715),
            .I(N__13712));
    Odrv4 I__1626 (
            .O(N__13712),
            .I(\eeprom.n3467 ));
    InMux I__1625 (
            .O(N__13709),
            .I(N__13706));
    LocalMux I__1624 (
            .O(N__13706),
            .I(N__13703));
    Span4Mux_h I__1623 (
            .O(N__13703),
            .I(N__13700));
    Odrv4 I__1622 (
            .O(N__13700),
            .I(\eeprom.n3466 ));
    CascadeMux I__1621 (
            .O(N__13697),
            .I(\eeprom.n3498_cascade_ ));
    CascadeMux I__1620 (
            .O(N__13694),
            .I(N__13691));
    InMux I__1619 (
            .O(N__13691),
            .I(N__13688));
    LocalMux I__1618 (
            .O(N__13688),
            .I(N__13685));
    Odrv4 I__1617 (
            .O(N__13685),
            .I(\eeprom.n28_adj_267 ));
    InMux I__1616 (
            .O(N__13682),
            .I(N__13679));
    LocalMux I__1615 (
            .O(N__13679),
            .I(N__13676));
    Odrv4 I__1614 (
            .O(N__13676),
            .I(\eeprom.n3476 ));
    InMux I__1613 (
            .O(N__13673),
            .I(N__13670));
    LocalMux I__1612 (
            .O(N__13670),
            .I(N__13667));
    Span4Mux_v I__1611 (
            .O(N__13667),
            .I(N__13664));
    Odrv4 I__1610 (
            .O(N__13664),
            .I(\eeprom.n3486 ));
    InMux I__1609 (
            .O(N__13661),
            .I(N__13658));
    LocalMux I__1608 (
            .O(N__13658),
            .I(N__13655));
    Span4Mux_h I__1607 (
            .O(N__13655),
            .I(N__13652));
    Odrv4 I__1606 (
            .O(N__13652),
            .I(\eeprom.n3468 ));
    CascadeMux I__1605 (
            .O(N__13649),
            .I(\eeprom.n3608_cascade_ ));
    InMux I__1604 (
            .O(N__13646),
            .I(N__13643));
    LocalMux I__1603 (
            .O(N__13643),
            .I(N__13640));
    Odrv4 I__1602 (
            .O(N__13640),
            .I(\eeprom.n3480 ));
    CascadeMux I__1601 (
            .O(N__13637),
            .I(\eeprom.n3512_cascade_ ));
    InMux I__1600 (
            .O(N__13634),
            .I(N__13631));
    LocalMux I__1599 (
            .O(N__13631),
            .I(\eeprom.n5175 ));
    CascadeMux I__1598 (
            .O(N__13628),
            .I(\eeprom.n5177_cascade_ ));
    InMux I__1597 (
            .O(N__13625),
            .I(N__13622));
    LocalMux I__1596 (
            .O(N__13622),
            .I(N__13619));
    Odrv4 I__1595 (
            .O(N__13619),
            .I(\eeprom.n31_adj_341 ));
    InMux I__1594 (
            .O(N__13616),
            .I(N__13613));
    LocalMux I__1593 (
            .O(N__13613),
            .I(N__13610));
    Odrv4 I__1592 (
            .O(N__13610),
            .I(\eeprom.n3598 ));
    InMux I__1591 (
            .O(N__13607),
            .I(N__13604));
    LocalMux I__1590 (
            .O(N__13604),
            .I(N__13601));
    Odrv12 I__1589 (
            .O(N__13601),
            .I(\eeprom.n3483 ));
    CascadeMux I__1588 (
            .O(N__13598),
            .I(\eeprom.n5031_cascade_ ));
    InMux I__1587 (
            .O(N__13595),
            .I(N__13592));
    LocalMux I__1586 (
            .O(N__13592),
            .I(\eeprom.n5161 ));
    InMux I__1585 (
            .O(N__13589),
            .I(N__13586));
    LocalMux I__1584 (
            .O(N__13586),
            .I(\eeprom.n29_adj_274 ));
    InMux I__1583 (
            .O(N__13583),
            .I(N__13580));
    LocalMux I__1582 (
            .O(N__13580),
            .I(N__13576));
    InMux I__1581 (
            .O(N__13579),
            .I(N__13573));
    Odrv4 I__1580 (
            .O(N__13576),
            .I(\eeprom.n3612 ));
    LocalMux I__1579 (
            .O(N__13573),
            .I(\eeprom.n3612 ));
    CascadeMux I__1578 (
            .O(N__13568),
            .I(N__13564));
    InMux I__1577 (
            .O(N__13567),
            .I(N__13561));
    InMux I__1576 (
            .O(N__13564),
            .I(N__13558));
    LocalMux I__1575 (
            .O(N__13561),
            .I(N__13552));
    LocalMux I__1574 (
            .O(N__13558),
            .I(N__13552));
    InMux I__1573 (
            .O(N__13557),
            .I(N__13549));
    Odrv4 I__1572 (
            .O(N__13552),
            .I(\eeprom.n3617 ));
    LocalMux I__1571 (
            .O(N__13549),
            .I(\eeprom.n3617 ));
    InMux I__1570 (
            .O(N__13544),
            .I(N__13541));
    LocalMux I__1569 (
            .O(N__13541),
            .I(N__13538));
    Odrv4 I__1568 (
            .O(N__13538),
            .I(\eeprom.n3596 ));
    CascadeMux I__1567 (
            .O(N__13535),
            .I(\eeprom.n3609_cascade_ ));
    CascadeMux I__1566 (
            .O(N__13532),
            .I(\eeprom.n5021_cascade_ ));
    InMux I__1565 (
            .O(N__13529),
            .I(N__13526));
    LocalMux I__1564 (
            .O(N__13526),
            .I(\eeprom.n5023 ));
    InMux I__1563 (
            .O(N__13523),
            .I(N__13520));
    LocalMux I__1562 (
            .O(N__13520),
            .I(N__13517));
    Span4Mux_h I__1561 (
            .O(N__13517),
            .I(N__13514));
    Odrv4 I__1560 (
            .O(N__13514),
            .I(\eeprom.n3474 ));
    InMux I__1559 (
            .O(N__13511),
            .I(N__13506));
    CascadeMux I__1558 (
            .O(N__13510),
            .I(N__13503));
    CascadeMux I__1557 (
            .O(N__13509),
            .I(N__13500));
    LocalMux I__1556 (
            .O(N__13506),
            .I(N__13497));
    InMux I__1555 (
            .O(N__13503),
            .I(N__13494));
    InMux I__1554 (
            .O(N__13500),
            .I(N__13491));
    Odrv4 I__1553 (
            .O(N__13497),
            .I(\eeprom.n3407 ));
    LocalMux I__1552 (
            .O(N__13494),
            .I(\eeprom.n3407 ));
    LocalMux I__1551 (
            .O(N__13491),
            .I(\eeprom.n3407 ));
    CascadeMux I__1550 (
            .O(N__13484),
            .I(\eeprom.n5019_cascade_ ));
    CascadeMux I__1549 (
            .O(N__13481),
            .I(\eeprom.n28_adj_342_cascade_ ));
    InMux I__1548 (
            .O(N__13478),
            .I(N__13474));
    InMux I__1547 (
            .O(N__13477),
            .I(N__13471));
    LocalMux I__1546 (
            .O(N__13474),
            .I(N__13468));
    LocalMux I__1545 (
            .O(N__13471),
            .I(\eeprom.n3615 ));
    Odrv4 I__1544 (
            .O(N__13468),
            .I(\eeprom.n3615 ));
    CascadeMux I__1543 (
            .O(N__13463),
            .I(\eeprom.n3628_cascade_ ));
    InMux I__1542 (
            .O(N__13460),
            .I(N__13457));
    LocalMux I__1541 (
            .O(N__13457),
            .I(\eeprom.n1204 ));
    CascadeMux I__1540 (
            .O(N__13454),
            .I(\eeprom.n3714_cascade_ ));
    CascadeMux I__1539 (
            .O(N__13451),
            .I(N__13447));
    InMux I__1538 (
            .O(N__13450),
            .I(N__13444));
    InMux I__1537 (
            .O(N__13447),
            .I(N__13441));
    LocalMux I__1536 (
            .O(N__13444),
            .I(\eeprom.n1201 ));
    LocalMux I__1535 (
            .O(N__13441),
            .I(\eeprom.n1201 ));
    CascadeMux I__1534 (
            .O(N__13436),
            .I(N__13431));
    InMux I__1533 (
            .O(N__13435),
            .I(N__13421));
    InMux I__1532 (
            .O(N__13434),
            .I(N__13421));
    InMux I__1531 (
            .O(N__13431),
            .I(N__13416));
    InMux I__1530 (
            .O(N__13430),
            .I(N__13416));
    InMux I__1529 (
            .O(N__13429),
            .I(N__13407));
    InMux I__1528 (
            .O(N__13428),
            .I(N__13407));
    InMux I__1527 (
            .O(N__13427),
            .I(N__13407));
    InMux I__1526 (
            .O(N__13426),
            .I(N__13407));
    LocalMux I__1525 (
            .O(N__13421),
            .I(\eeprom.n3628 ));
    LocalMux I__1524 (
            .O(N__13416),
            .I(\eeprom.n3628 ));
    LocalMux I__1523 (
            .O(N__13407),
            .I(\eeprom.n3628 ));
    CascadeMux I__1522 (
            .O(N__13400),
            .I(\eeprom.n5025_cascade_ ));
    CascadeMux I__1521 (
            .O(N__13397),
            .I(\eeprom.n5027_cascade_ ));
    CascadeMux I__1520 (
            .O(N__13394),
            .I(\eeprom.n5029_cascade_ ));
    CascadeMux I__1519 (
            .O(N__13391),
            .I(\eeprom.n3712_cascade_ ));
    InMux I__1518 (
            .O(N__13388),
            .I(N__13385));
    LocalMux I__1517 (
            .O(N__13385),
            .I(\eeprom.n1207 ));
    CascadeMux I__1516 (
            .O(N__13382),
            .I(N__13379));
    InMux I__1515 (
            .O(N__13379),
            .I(N__13375));
    InMux I__1514 (
            .O(N__13378),
            .I(N__13372));
    LocalMux I__1513 (
            .O(N__13375),
            .I(\eeprom.n3618 ));
    LocalMux I__1512 (
            .O(N__13372),
            .I(\eeprom.n3618 ));
    CascadeMux I__1511 (
            .O(N__13367),
            .I(\eeprom.n3717_cascade_ ));
    InMux I__1510 (
            .O(N__13364),
            .I(N__13361));
    LocalMux I__1509 (
            .O(N__13361),
            .I(\eeprom.n1208 ));
    CascadeMux I__1508 (
            .O(N__13358),
            .I(\eeprom.n5362_cascade_ ));
    CascadeMux I__1507 (
            .O(N__13355),
            .I(N__13352));
    InMux I__1506 (
            .O(N__13352),
            .I(N__13349));
    LocalMux I__1505 (
            .O(N__13349),
            .I(\eeprom.n1206 ));
    InMux I__1504 (
            .O(N__13346),
            .I(N__13343));
    LocalMux I__1503 (
            .O(N__13343),
            .I(\eeprom.n1205 ));
    CascadeMux I__1502 (
            .O(N__13340),
            .I(N__13336));
    CascadeMux I__1501 (
            .O(N__13339),
            .I(N__13333));
    InMux I__1500 (
            .O(N__13336),
            .I(N__13330));
    InMux I__1499 (
            .O(N__13333),
            .I(N__13326));
    LocalMux I__1498 (
            .O(N__13330),
            .I(N__13323));
    InMux I__1497 (
            .O(N__13329),
            .I(N__13320));
    LocalMux I__1496 (
            .O(N__13326),
            .I(\eeprom.n3616 ));
    Odrv4 I__1495 (
            .O(N__13323),
            .I(\eeprom.n3616 ));
    LocalMux I__1494 (
            .O(N__13320),
            .I(\eeprom.n3616 ));
    CascadeMux I__1493 (
            .O(N__13313),
            .I(\eeprom.n3715_cascade_ ));
    InMux I__1492 (
            .O(N__13310),
            .I(N__13307));
    LocalMux I__1491 (
            .O(N__13307),
            .I(\eeprom.n5017 ));
    InMux I__1490 (
            .O(N__13304),
            .I(\eeprom.n4116 ));
    InMux I__1489 (
            .O(N__13301),
            .I(\eeprom.n4117 ));
    InMux I__1488 (
            .O(N__13298),
            .I(\eeprom.n4118 ));
    InMux I__1487 (
            .O(N__13295),
            .I(\eeprom.n4119 ));
    InMux I__1486 (
            .O(N__13292),
            .I(N__13289));
    LocalMux I__1485 (
            .O(N__13289),
            .I(N__13286));
    Span4Mux_h I__1484 (
            .O(N__13286),
            .I(N__13283));
    Odrv4 I__1483 (
            .O(N__13283),
            .I(\eeprom.n3070 ));
    InMux I__1482 (
            .O(N__13280),
            .I(bfn_18_31_0_));
    CascadeMux I__1481 (
            .O(N__13277),
            .I(N__13274));
    InMux I__1480 (
            .O(N__13274),
            .I(N__13271));
    LocalMux I__1479 (
            .O(N__13271),
            .I(N__13268));
    Span4Mux_h I__1478 (
            .O(N__13268),
            .I(N__13265));
    Odrv4 I__1477 (
            .O(N__13265),
            .I(\eeprom.n3069 ));
    InMux I__1476 (
            .O(N__13262),
            .I(\eeprom.n4121 ));
    InMux I__1475 (
            .O(N__13259),
            .I(\eeprom.n4122 ));
    InMux I__1474 (
            .O(N__13256),
            .I(N__13253));
    LocalMux I__1473 (
            .O(N__13253),
            .I(\eeprom.n3071 ));
    CascadeMux I__1472 (
            .O(N__13250),
            .I(N__13247));
    InMux I__1471 (
            .O(N__13247),
            .I(N__13242));
    InMux I__1470 (
            .O(N__13246),
            .I(N__13239));
    InMux I__1469 (
            .O(N__13245),
            .I(N__13236));
    LocalMux I__1468 (
            .O(N__13242),
            .I(N__13231));
    LocalMux I__1467 (
            .O(N__13239),
            .I(N__13231));
    LocalMux I__1466 (
            .O(N__13236),
            .I(\eeprom.n3004 ));
    Odrv4 I__1465 (
            .O(N__13231),
            .I(\eeprom.n3004 ));
    InMux I__1464 (
            .O(N__13226),
            .I(N__13222));
    InMux I__1463 (
            .O(N__13225),
            .I(N__13219));
    LocalMux I__1462 (
            .O(N__13222),
            .I(N__13215));
    LocalMux I__1461 (
            .O(N__13219),
            .I(N__13212));
    InMux I__1460 (
            .O(N__13218),
            .I(N__13209));
    Odrv4 I__1459 (
            .O(N__13215),
            .I(\eeprom.n3613 ));
    Odrv4 I__1458 (
            .O(N__13212),
            .I(\eeprom.n3613 ));
    LocalMux I__1457 (
            .O(N__13209),
            .I(\eeprom.n3613 ));
    CascadeMux I__1456 (
            .O(N__13202),
            .I(N__13199));
    InMux I__1455 (
            .O(N__13199),
            .I(N__13196));
    LocalMux I__1454 (
            .O(N__13196),
            .I(\eeprom.n1202 ));
    InMux I__1453 (
            .O(N__13193),
            .I(N__13190));
    LocalMux I__1452 (
            .O(N__13190),
            .I(\eeprom.n3083 ));
    InMux I__1451 (
            .O(N__13187),
            .I(\eeprom.n4107 ));
    InMux I__1450 (
            .O(N__13184),
            .I(\eeprom.n4108 ));
    InMux I__1449 (
            .O(N__13181),
            .I(N__13178));
    LocalMux I__1448 (
            .O(N__13178),
            .I(N__13175));
    Odrv4 I__1447 (
            .O(N__13175),
            .I(\eeprom.n3081 ));
    InMux I__1446 (
            .O(N__13172),
            .I(\eeprom.n4109 ));
    InMux I__1445 (
            .O(N__13169),
            .I(\eeprom.n4110 ));
    InMux I__1444 (
            .O(N__13166),
            .I(N__13163));
    LocalMux I__1443 (
            .O(N__13163),
            .I(\eeprom.n3079 ));
    InMux I__1442 (
            .O(N__13160),
            .I(\eeprom.n4111 ));
    InMux I__1441 (
            .O(N__13157),
            .I(bfn_18_30_0_));
    CascadeMux I__1440 (
            .O(N__13154),
            .I(N__13151));
    InMux I__1439 (
            .O(N__13151),
            .I(N__13148));
    LocalMux I__1438 (
            .O(N__13148),
            .I(N__13145));
    Odrv4 I__1437 (
            .O(N__13145),
            .I(\eeprom.n3077 ));
    InMux I__1436 (
            .O(N__13142),
            .I(\eeprom.n4113 ));
    InMux I__1435 (
            .O(N__13139),
            .I(N__13136));
    LocalMux I__1434 (
            .O(N__13136),
            .I(N__13133));
    Odrv12 I__1433 (
            .O(N__13133),
            .I(\eeprom.n3076 ));
    InMux I__1432 (
            .O(N__13130),
            .I(\eeprom.n4114 ));
    InMux I__1431 (
            .O(N__13127),
            .I(N__13124));
    LocalMux I__1430 (
            .O(N__13124),
            .I(N__13121));
    Odrv4 I__1429 (
            .O(N__13121),
            .I(\eeprom.n3075 ));
    InMux I__1428 (
            .O(N__13118),
            .I(\eeprom.n4115 ));
    CascadeMux I__1427 (
            .O(N__13115),
            .I(\eeprom.n3034_cascade_ ));
    InMux I__1426 (
            .O(N__13112),
            .I(bfn_18_29_0_));
    InMux I__1425 (
            .O(N__13109),
            .I(N__13106));
    LocalMux I__1424 (
            .O(N__13106),
            .I(\eeprom.n3085 ));
    InMux I__1423 (
            .O(N__13103),
            .I(\eeprom.n4105 ));
    CascadeMux I__1422 (
            .O(N__13100),
            .I(N__13097));
    InMux I__1421 (
            .O(N__13097),
            .I(N__13094));
    LocalMux I__1420 (
            .O(N__13094),
            .I(N__13091));
    Odrv4 I__1419 (
            .O(N__13091),
            .I(\eeprom.n3084 ));
    InMux I__1418 (
            .O(N__13088),
            .I(\eeprom.n4106 ));
    InMux I__1417 (
            .O(N__13085),
            .I(N__13082));
    LocalMux I__1416 (
            .O(N__13082),
            .I(N__13079));
    Odrv4 I__1415 (
            .O(N__13079),
            .I(\eeprom.n3270 ));
    CascadeMux I__1414 (
            .O(N__13076),
            .I(\eeprom.n3203_cascade_ ));
    CascadeMux I__1413 (
            .O(N__13073),
            .I(\eeprom.n3113_cascade_ ));
    CascadeMux I__1412 (
            .O(N__13070),
            .I(\eeprom.n5305_cascade_ ));
    InMux I__1411 (
            .O(N__13067),
            .I(N__13064));
    LocalMux I__1410 (
            .O(N__13064),
            .I(N__13061));
    Odrv4 I__1409 (
            .O(N__13061),
            .I(\eeprom.n3273 ));
    CascadeMux I__1408 (
            .O(N__13058),
            .I(\eeprom.n3206_cascade_ ));
    CascadeMux I__1407 (
            .O(N__13055),
            .I(\eeprom.n3108_cascade_ ));
    CascadeMux I__1406 (
            .O(N__13052),
            .I(N__13049));
    InMux I__1405 (
            .O(N__13049),
            .I(N__13045));
    InMux I__1404 (
            .O(N__13048),
            .I(N__13042));
    LocalMux I__1403 (
            .O(N__13045),
            .I(N__13039));
    LocalMux I__1402 (
            .O(N__13042),
            .I(N__13036));
    Span4Mux_v I__1401 (
            .O(N__13039),
            .I(N__13030));
    Span4Mux_h I__1400 (
            .O(N__13036),
            .I(N__13030));
    InMux I__1399 (
            .O(N__13035),
            .I(N__13027));
    Odrv4 I__1398 (
            .O(N__13030),
            .I(\eeprom.n3202 ));
    LocalMux I__1397 (
            .O(N__13027),
            .I(\eeprom.n3202 ));
    CascadeMux I__1396 (
            .O(N__13022),
            .I(N__13018));
    InMux I__1395 (
            .O(N__13021),
            .I(N__13015));
    InMux I__1394 (
            .O(N__13018),
            .I(N__13012));
    LocalMux I__1393 (
            .O(N__13015),
            .I(N__13008));
    LocalMux I__1392 (
            .O(N__13012),
            .I(N__13005));
    InMux I__1391 (
            .O(N__13011),
            .I(N__13002));
    Odrv4 I__1390 (
            .O(N__13008),
            .I(\eeprom.n3201 ));
    Odrv4 I__1389 (
            .O(N__13005),
            .I(\eeprom.n3201 ));
    LocalMux I__1388 (
            .O(N__13002),
            .I(\eeprom.n3201 ));
    CascadeMux I__1387 (
            .O(N__12995),
            .I(N__12992));
    InMux I__1386 (
            .O(N__12992),
            .I(N__12989));
    LocalMux I__1385 (
            .O(N__12989),
            .I(N__12985));
    InMux I__1384 (
            .O(N__12988),
            .I(N__12982));
    Odrv4 I__1383 (
            .O(N__12985),
            .I(\eeprom.n3203 ));
    LocalMux I__1382 (
            .O(N__12982),
            .I(\eeprom.n3203 ));
    CascadeMux I__1381 (
            .O(N__12977),
            .I(N__12974));
    InMux I__1380 (
            .O(N__12974),
            .I(N__12970));
    CascadeMux I__1379 (
            .O(N__12973),
            .I(N__12967));
    LocalMux I__1378 (
            .O(N__12970),
            .I(N__12964));
    InMux I__1377 (
            .O(N__12967),
            .I(N__12961));
    Span4Mux_v I__1376 (
            .O(N__12964),
            .I(N__12958));
    LocalMux I__1375 (
            .O(N__12961),
            .I(\eeprom.n3200 ));
    Odrv4 I__1374 (
            .O(N__12958),
            .I(\eeprom.n3200 ));
    CascadeMux I__1373 (
            .O(N__12953),
            .I(\eeprom.n3200_cascade_ ));
    InMux I__1372 (
            .O(N__12950),
            .I(N__12947));
    LocalMux I__1371 (
            .O(N__12947),
            .I(N__12944));
    Span4Mux_h I__1370 (
            .O(N__12944),
            .I(N__12941));
    Odrv4 I__1369 (
            .O(N__12941),
            .I(\eeprom.n3286 ));
    InMux I__1368 (
            .O(N__12938),
            .I(N__12935));
    LocalMux I__1367 (
            .O(N__12935),
            .I(N__12932));
    Span4Mux_h I__1366 (
            .O(N__12932),
            .I(N__12929));
    Odrv4 I__1365 (
            .O(N__12929),
            .I(\eeprom.n3280 ));
    InMux I__1364 (
            .O(N__12926),
            .I(N__12923));
    LocalMux I__1363 (
            .O(N__12923),
            .I(N__12920));
    Span4Mux_h I__1362 (
            .O(N__12920),
            .I(N__12917));
    Odrv4 I__1361 (
            .O(N__12917),
            .I(\eeprom.n3275 ));
    InMux I__1360 (
            .O(N__12914),
            .I(N__12911));
    LocalMux I__1359 (
            .O(N__12911),
            .I(N__12908));
    Span4Mux_h I__1358 (
            .O(N__12908),
            .I(N__12905));
    Odrv4 I__1357 (
            .O(N__12905),
            .I(\eeprom.n3276 ));
    InMux I__1356 (
            .O(N__12902),
            .I(N__12899));
    LocalMux I__1355 (
            .O(N__12899),
            .I(N__12896));
    Span4Mux_h I__1354 (
            .O(N__12896),
            .I(N__12893));
    Odrv4 I__1353 (
            .O(N__12893),
            .I(\eeprom.n3279 ));
    CascadeMux I__1352 (
            .O(N__12890),
            .I(\eeprom.n3204_cascade_ ));
    InMux I__1351 (
            .O(N__12887),
            .I(N__12884));
    LocalMux I__1350 (
            .O(N__12884),
            .I(N__12881));
    Span4Mux_v I__1349 (
            .O(N__12881),
            .I(N__12878));
    Odrv4 I__1348 (
            .O(N__12878),
            .I(\eeprom.n3267 ));
    CascadeMux I__1347 (
            .O(N__12875),
            .I(\eeprom.n3299_cascade_ ));
    CascadeMux I__1346 (
            .O(N__12872),
            .I(N__12868));
    InMux I__1345 (
            .O(N__12871),
            .I(N__12865));
    InMux I__1344 (
            .O(N__12868),
            .I(N__12862));
    LocalMux I__1343 (
            .O(N__12865),
            .I(N__12859));
    LocalMux I__1342 (
            .O(N__12862),
            .I(N__12854));
    Span4Mux_v I__1341 (
            .O(N__12859),
            .I(N__12854));
    Odrv4 I__1340 (
            .O(N__12854),
            .I(\eeprom.n3298 ));
    InMux I__1339 (
            .O(N__12851),
            .I(N__12848));
    LocalMux I__1338 (
            .O(N__12848),
            .I(\eeprom.n3379 ));
    InMux I__1337 (
            .O(N__12845),
            .I(N__12841));
    CascadeMux I__1336 (
            .O(N__12844),
            .I(N__12838));
    LocalMux I__1335 (
            .O(N__12841),
            .I(N__12835));
    InMux I__1334 (
            .O(N__12838),
            .I(N__12832));
    Span4Mux_v I__1333 (
            .O(N__12835),
            .I(N__12829));
    LocalMux I__1332 (
            .O(N__12832),
            .I(\eeprom.n3299 ));
    Odrv4 I__1331 (
            .O(N__12829),
            .I(\eeprom.n3299 ));
    InMux I__1330 (
            .O(N__12824),
            .I(N__12821));
    LocalMux I__1329 (
            .O(N__12821),
            .I(N__12818));
    Odrv4 I__1328 (
            .O(N__12818),
            .I(\eeprom.n3366 ));
    InMux I__1327 (
            .O(N__12815),
            .I(N__12812));
    LocalMux I__1326 (
            .O(N__12812),
            .I(N__12809));
    Span4Mux_v I__1325 (
            .O(N__12809),
            .I(N__12806));
    Odrv4 I__1324 (
            .O(N__12806),
            .I(\eeprom.n3269 ));
    CascadeMux I__1323 (
            .O(N__12803),
            .I(N__12800));
    InMux I__1322 (
            .O(N__12800),
            .I(N__12797));
    LocalMux I__1321 (
            .O(N__12797),
            .I(N__12793));
    InMux I__1320 (
            .O(N__12796),
            .I(N__12790));
    Odrv4 I__1319 (
            .O(N__12793),
            .I(\eeprom.n3301 ));
    LocalMux I__1318 (
            .O(N__12790),
            .I(\eeprom.n3301 ));
    CascadeMux I__1317 (
            .O(N__12785),
            .I(\eeprom.n3301_cascade_ ));
    InMux I__1316 (
            .O(N__12782),
            .I(N__12779));
    LocalMux I__1315 (
            .O(N__12779),
            .I(N__12776));
    Odrv4 I__1314 (
            .O(N__12776),
            .I(\eeprom.n3368 ));
    InMux I__1313 (
            .O(N__12773),
            .I(N__12770));
    LocalMux I__1312 (
            .O(N__12770),
            .I(N__12767));
    Odrv4 I__1311 (
            .O(N__12767),
            .I(\eeprom.n3374 ));
    CascadeMux I__1310 (
            .O(N__12764),
            .I(N__12761));
    InMux I__1309 (
            .O(N__12761),
            .I(N__12758));
    LocalMux I__1308 (
            .O(N__12758),
            .I(N__12754));
    CascadeMux I__1307 (
            .O(N__12757),
            .I(N__12751));
    Span4Mux_v I__1306 (
            .O(N__12754),
            .I(N__12747));
    InMux I__1305 (
            .O(N__12751),
            .I(N__12744));
    InMux I__1304 (
            .O(N__12750),
            .I(N__12741));
    Odrv4 I__1303 (
            .O(N__12747),
            .I(\eeprom.n3406 ));
    LocalMux I__1302 (
            .O(N__12744),
            .I(\eeprom.n3406 ));
    LocalMux I__1301 (
            .O(N__12741),
            .I(\eeprom.n3406 ));
    CascadeMux I__1300 (
            .O(N__12734),
            .I(N__12731));
    InMux I__1299 (
            .O(N__12731),
            .I(N__12728));
    LocalMux I__1298 (
            .O(N__12728),
            .I(N__12725));
    Odrv4 I__1297 (
            .O(N__12725),
            .I(\eeprom.n3370 ));
    InMux I__1296 (
            .O(N__12722),
            .I(N__12719));
    LocalMux I__1295 (
            .O(N__12719),
            .I(N__12716));
    Span4Mux_v I__1294 (
            .O(N__12716),
            .I(N__12713));
    Odrv4 I__1293 (
            .O(N__12713),
            .I(\eeprom.n3268 ));
    InMux I__1292 (
            .O(N__12710),
            .I(N__12707));
    LocalMux I__1291 (
            .O(N__12707),
            .I(N__12702));
    InMux I__1290 (
            .O(N__12706),
            .I(N__12697));
    InMux I__1289 (
            .O(N__12705),
            .I(N__12697));
    Odrv4 I__1288 (
            .O(N__12702),
            .I(\eeprom.n3300 ));
    LocalMux I__1287 (
            .O(N__12697),
            .I(\eeprom.n3300 ));
    InMux I__1286 (
            .O(N__12692),
            .I(N__12689));
    LocalMux I__1285 (
            .O(N__12689),
            .I(N__12686));
    Span4Mux_h I__1284 (
            .O(N__12686),
            .I(N__12683));
    Odrv4 I__1283 (
            .O(N__12683),
            .I(\eeprom.n3376 ));
    CascadeMux I__1282 (
            .O(N__12680),
            .I(N__12677));
    InMux I__1281 (
            .O(N__12677),
            .I(N__12674));
    LocalMux I__1280 (
            .O(N__12674),
            .I(N__12671));
    Span4Mux_v I__1279 (
            .O(N__12671),
            .I(N__12668));
    Odrv4 I__1278 (
            .O(N__12668),
            .I(\eeprom.n3380 ));
    CascadeMux I__1277 (
            .O(N__12665),
            .I(N__12661));
    InMux I__1276 (
            .O(N__12664),
            .I(N__12658));
    InMux I__1275 (
            .O(N__12661),
            .I(N__12655));
    LocalMux I__1274 (
            .O(N__12658),
            .I(\eeprom.n3412 ));
    LocalMux I__1273 (
            .O(N__12655),
            .I(\eeprom.n3412 ));
    CascadeMux I__1272 (
            .O(N__12650),
            .I(\eeprom.n3412_cascade_ ));
    InMux I__1271 (
            .O(N__12647),
            .I(N__12644));
    LocalMux I__1270 (
            .O(N__12644),
            .I(\eeprom.n3479 ));
    InMux I__1269 (
            .O(N__12641),
            .I(N__12638));
    LocalMux I__1268 (
            .O(N__12638),
            .I(N__12635));
    Odrv4 I__1267 (
            .O(N__12635),
            .I(\eeprom.n3375 ));
    InMux I__1266 (
            .O(N__12632),
            .I(N__12629));
    LocalMux I__1265 (
            .O(N__12629),
            .I(N__12626));
    Odrv4 I__1264 (
            .O(N__12626),
            .I(\eeprom.n3378 ));
    CascadeMux I__1263 (
            .O(N__12623),
            .I(N__12619));
    InMux I__1262 (
            .O(N__12622),
            .I(N__12616));
    InMux I__1261 (
            .O(N__12619),
            .I(N__12613));
    LocalMux I__1260 (
            .O(N__12616),
            .I(\eeprom.n3410 ));
    LocalMux I__1259 (
            .O(N__12613),
            .I(\eeprom.n3410 ));
    InMux I__1258 (
            .O(N__12608),
            .I(N__12605));
    LocalMux I__1257 (
            .O(N__12605),
            .I(\eeprom.n3477 ));
    CascadeMux I__1256 (
            .O(N__12602),
            .I(\eeprom.n3410_cascade_ ));
    InMux I__1255 (
            .O(N__12599),
            .I(N__12596));
    LocalMux I__1254 (
            .O(N__12596),
            .I(\eeprom.n3465 ));
    InMux I__1253 (
            .O(N__12593),
            .I(N__12590));
    LocalMux I__1252 (
            .O(N__12590),
            .I(N__12587));
    Span4Mux_h I__1251 (
            .O(N__12587),
            .I(N__12584));
    Odrv4 I__1250 (
            .O(N__12584),
            .I(\eeprom.n3367 ));
    CascadeMux I__1249 (
            .O(N__12581),
            .I(\eeprom.n3505_cascade_ ));
    InMux I__1248 (
            .O(N__12578),
            .I(N__12575));
    LocalMux I__1247 (
            .O(N__12575),
            .I(\eeprom.n30_adj_273 ));
    InMux I__1246 (
            .O(N__12572),
            .I(N__12569));
    LocalMux I__1245 (
            .O(N__12569),
            .I(\eeprom.n3478 ));
    InMux I__1244 (
            .O(N__12566),
            .I(N__12563));
    LocalMux I__1243 (
            .O(N__12563),
            .I(\eeprom.n3472 ));
    InMux I__1242 (
            .O(N__12560),
            .I(N__12557));
    LocalMux I__1241 (
            .O(N__12557),
            .I(\eeprom.n3484 ));
    CascadeMux I__1240 (
            .O(N__12554),
            .I(N__12551));
    InMux I__1239 (
            .O(N__12551),
            .I(N__12548));
    LocalMux I__1238 (
            .O(N__12548),
            .I(\eeprom.n3475 ));
    CascadeMux I__1237 (
            .O(N__12545),
            .I(\eeprom.n3507_cascade_ ));
    InMux I__1236 (
            .O(N__12542),
            .I(N__12539));
    LocalMux I__1235 (
            .O(N__12539),
            .I(\eeprom.n31 ));
    CascadeMux I__1234 (
            .O(N__12536),
            .I(N__12533));
    InMux I__1233 (
            .O(N__12533),
            .I(N__12530));
    LocalMux I__1232 (
            .O(N__12530),
            .I(\eeprom.n3482 ));
    CascadeMux I__1231 (
            .O(N__12527),
            .I(\eeprom.n3514_cascade_ ));
    CascadeMux I__1230 (
            .O(N__12524),
            .I(\eeprom.n5323_cascade_ ));
    InMux I__1229 (
            .O(N__12521),
            .I(N__12518));
    LocalMux I__1228 (
            .O(N__12518),
            .I(\eeprom.n5321 ));
    InMux I__1227 (
            .O(N__12515),
            .I(N__12512));
    LocalMux I__1226 (
            .O(N__12512),
            .I(\eeprom.n4753 ));
    InMux I__1225 (
            .O(N__12509),
            .I(N__12506));
    LocalMux I__1224 (
            .O(N__12506),
            .I(\eeprom.n3605 ));
    CascadeMux I__1223 (
            .O(N__12503),
            .I(N__12500));
    InMux I__1222 (
            .O(N__12500),
            .I(N__12497));
    LocalMux I__1221 (
            .O(N__12497),
            .I(N__12494));
    Span4Mux_v I__1220 (
            .O(N__12494),
            .I(N__12491));
    Odrv4 I__1219 (
            .O(N__12491),
            .I(\eeprom.n3471 ));
    CascadeMux I__1218 (
            .O(N__12488),
            .I(\eeprom.n32_cascade_ ));
    CascadeMux I__1217 (
            .O(N__12485),
            .I(\eeprom.n3529_cascade_ ));
    InMux I__1216 (
            .O(N__12482),
            .I(N__12479));
    LocalMux I__1215 (
            .O(N__12479),
            .I(\eeprom.n3481 ));
    CascadeMux I__1214 (
            .O(N__12476),
            .I(\eeprom.n3513_cascade_ ));
    InMux I__1213 (
            .O(N__12473),
            .I(N__12470));
    LocalMux I__1212 (
            .O(N__12470),
            .I(N__12467));
    Odrv4 I__1211 (
            .O(N__12467),
            .I(\eeprom.n3473 ));
    InMux I__1210 (
            .O(N__12464),
            .I(N__12458));
    InMux I__1209 (
            .O(N__12463),
            .I(N__12458));
    LocalMux I__1208 (
            .O(N__12458),
            .I(N__12454));
    InMux I__1207 (
            .O(N__12457),
            .I(N__12451));
    Odrv4 I__1206 (
            .O(N__12454),
            .I(blink_counter_24));
    LocalMux I__1205 (
            .O(N__12451),
            .I(blink_counter_24));
    InMux I__1204 (
            .O(N__12446),
            .I(N__12439));
    InMux I__1203 (
            .O(N__12445),
            .I(N__12439));
    InMux I__1202 (
            .O(N__12444),
            .I(N__12436));
    LocalMux I__1201 (
            .O(N__12439),
            .I(blink_counter_22));
    LocalMux I__1200 (
            .O(N__12436),
            .I(blink_counter_22));
    CascadeMux I__1199 (
            .O(N__12431),
            .I(N__12427));
    CascadeMux I__1198 (
            .O(N__12430),
            .I(N__12424));
    InMux I__1197 (
            .O(N__12427),
            .I(N__12418));
    InMux I__1196 (
            .O(N__12424),
            .I(N__12418));
    InMux I__1195 (
            .O(N__12423),
            .I(N__12415));
    LocalMux I__1194 (
            .O(N__12418),
            .I(blink_counter_23));
    LocalMux I__1193 (
            .O(N__12415),
            .I(blink_counter_23));
    InMux I__1192 (
            .O(N__12410),
            .I(N__12403));
    InMux I__1191 (
            .O(N__12409),
            .I(N__12403));
    InMux I__1190 (
            .O(N__12408),
            .I(N__12400));
    LocalMux I__1189 (
            .O(N__12403),
            .I(blink_counter_21));
    LocalMux I__1188 (
            .O(N__12400),
            .I(blink_counter_21));
    InMux I__1187 (
            .O(N__12395),
            .I(N__12392));
    LocalMux I__1186 (
            .O(N__12392),
            .I(N__12389));
    Span4Mux_v I__1185 (
            .O(N__12389),
            .I(N__12386));
    Odrv4 I__1184 (
            .O(N__12386),
            .I(n5420));
    CascadeMux I__1183 (
            .O(N__12383),
            .I(N__12380));
    InMux I__1182 (
            .O(N__12380),
            .I(N__12377));
    LocalMux I__1181 (
            .O(N__12377),
            .I(\eeprom.n1203 ));
    CascadeMux I__1180 (
            .O(N__12374),
            .I(\eeprom.n3713_cascade_ ));
    CascadeMux I__1179 (
            .O(N__12371),
            .I(\eeprom.n3618_cascade_ ));
    CascadeMux I__1178 (
            .O(N__12368),
            .I(\eeprom.n3615_cascade_ ));
    CascadeMux I__1177 (
            .O(N__12365),
            .I(\eeprom.n5221_cascade_ ));
    InMux I__1176 (
            .O(N__12362),
            .I(N__12359));
    LocalMux I__1175 (
            .O(N__12359),
            .I(\eeprom.n5225 ));
    CascadeMux I__1174 (
            .O(N__12356),
            .I(N__12353));
    InMux I__1173 (
            .O(N__12353),
            .I(N__12349));
    InMux I__1172 (
            .O(N__12352),
            .I(N__12345));
    LocalMux I__1171 (
            .O(N__12349),
            .I(N__12342));
    InMux I__1170 (
            .O(N__12348),
            .I(N__12339));
    LocalMux I__1169 (
            .O(N__12345),
            .I(\eeprom.n3614 ));
    Odrv4 I__1168 (
            .O(N__12342),
            .I(\eeprom.n3614 ));
    LocalMux I__1167 (
            .O(N__12339),
            .I(\eeprom.n3614 ));
    InMux I__1166 (
            .O(N__12332),
            .I(\eeprom.n3966 ));
    InMux I__1165 (
            .O(N__12329),
            .I(\eeprom.n3967 ));
    InMux I__1164 (
            .O(N__12326),
            .I(\eeprom.n3968 ));
    InMux I__1163 (
            .O(N__12323),
            .I(\eeprom.n3969 ));
    InMux I__1162 (
            .O(N__12320),
            .I(\eeprom.n3970 ));
    InMux I__1161 (
            .O(N__12317),
            .I(\eeprom.n3971 ));
    InMux I__1160 (
            .O(N__12314),
            .I(\eeprom.n3972 ));
    InMux I__1159 (
            .O(N__12311),
            .I(N__12308));
    LocalMux I__1158 (
            .O(N__12308),
            .I(N__12305));
    Span4Mux_v I__1157 (
            .O(N__12305),
            .I(N__12302));
    Odrv4 I__1156 (
            .O(N__12302),
            .I(n5421));
    InMux I__1155 (
            .O(N__12299),
            .I(\eeprom.n4155 ));
    InMux I__1154 (
            .O(N__12296),
            .I(\eeprom.n4156 ));
    InMux I__1153 (
            .O(N__12293),
            .I(bfn_17_29_0_));
    InMux I__1152 (
            .O(N__12290),
            .I(\eeprom.n4158 ));
    InMux I__1151 (
            .O(N__12287),
            .I(\eeprom.n4159 ));
    InMux I__1150 (
            .O(N__12284),
            .I(\eeprom.n4160 ));
    InMux I__1149 (
            .O(N__12281),
            .I(\eeprom.n4161 ));
    InMux I__1148 (
            .O(N__12278),
            .I(bfn_18_17_0_));
    InMux I__1147 (
            .O(N__12275),
            .I(\eeprom.n4146 ));
    InMux I__1146 (
            .O(N__12272),
            .I(\eeprom.n4147 ));
    InMux I__1145 (
            .O(N__12269),
            .I(\eeprom.n4148 ));
    InMux I__1144 (
            .O(N__12266),
            .I(bfn_17_28_0_));
    CascadeMux I__1143 (
            .O(N__12263),
            .I(N__12260));
    InMux I__1142 (
            .O(N__12260),
            .I(N__12257));
    LocalMux I__1141 (
            .O(N__12257),
            .I(N__12254));
    Odrv4 I__1140 (
            .O(N__12254),
            .I(\eeprom.n3277 ));
    InMux I__1139 (
            .O(N__12251),
            .I(\eeprom.n4150 ));
    InMux I__1138 (
            .O(N__12248),
            .I(\eeprom.n4151 ));
    InMux I__1137 (
            .O(N__12245),
            .I(\eeprom.n4152 ));
    InMux I__1136 (
            .O(N__12242),
            .I(\eeprom.n4153 ));
    InMux I__1135 (
            .O(N__12239),
            .I(\eeprom.n4154 ));
    InMux I__1134 (
            .O(N__12236),
            .I(\eeprom.n4179 ));
    InMux I__1133 (
            .O(N__12233),
            .I(\eeprom.n4180 ));
    InMux I__1132 (
            .O(N__12230),
            .I(\eeprom.n4181 ));
    InMux I__1131 (
            .O(N__12227),
            .I(\eeprom.n4182 ));
    InMux I__1130 (
            .O(N__12224),
            .I(bfn_17_27_0_));
    InMux I__1129 (
            .O(N__12221),
            .I(\eeprom.n4142 ));
    InMux I__1128 (
            .O(N__12218),
            .I(\eeprom.n4143 ));
    InMux I__1127 (
            .O(N__12215),
            .I(\eeprom.n4144 ));
    InMux I__1126 (
            .O(N__12212),
            .I(\eeprom.n4145 ));
    InMux I__1125 (
            .O(N__12209),
            .I(\eeprom.n4170 ));
    InMux I__1124 (
            .O(N__12206),
            .I(\eeprom.n4171 ));
    InMux I__1123 (
            .O(N__12203),
            .I(\eeprom.n4172 ));
    InMux I__1122 (
            .O(N__12200),
            .I(\eeprom.n4173 ));
    InMux I__1121 (
            .O(N__12197),
            .I(\eeprom.n4174 ));
    CascadeMux I__1120 (
            .O(N__12194),
            .I(N__12191));
    InMux I__1119 (
            .O(N__12191),
            .I(N__12188));
    LocalMux I__1118 (
            .O(N__12188),
            .I(N__12185));
    Odrv4 I__1117 (
            .O(N__12185),
            .I(\eeprom.n3372 ));
    InMux I__1116 (
            .O(N__12182),
            .I(\eeprom.n4175 ));
    InMux I__1115 (
            .O(N__12179),
            .I(\eeprom.n4176 ));
    InMux I__1114 (
            .O(N__12176),
            .I(bfn_17_26_0_));
    InMux I__1113 (
            .O(N__12173),
            .I(\eeprom.n4178 ));
    InMux I__1112 (
            .O(N__12170),
            .I(bfn_17_24_0_));
    InMux I__1111 (
            .O(N__12167),
            .I(\eeprom.n4162 ));
    InMux I__1110 (
            .O(N__12164),
            .I(\eeprom.n4163 ));
    InMux I__1109 (
            .O(N__12161),
            .I(\eeprom.n4164 ));
    InMux I__1108 (
            .O(N__12158),
            .I(\eeprom.n4165 ));
    InMux I__1107 (
            .O(N__12155),
            .I(\eeprom.n4166 ));
    InMux I__1106 (
            .O(N__12152),
            .I(\eeprom.n4167 ));
    InMux I__1105 (
            .O(N__12149),
            .I(\eeprom.n4168 ));
    InMux I__1104 (
            .O(N__12146),
            .I(bfn_17_25_0_));
    InMux I__1103 (
            .O(N__12143),
            .I(\eeprom.n4197 ));
    InMux I__1102 (
            .O(N__12140),
            .I(bfn_17_23_0_));
    InMux I__1101 (
            .O(N__12137),
            .I(\eeprom.n4199 ));
    InMux I__1100 (
            .O(N__12134),
            .I(\eeprom.n4200 ));
    InMux I__1099 (
            .O(N__12131),
            .I(\eeprom.n4201 ));
    InMux I__1098 (
            .O(N__12128),
            .I(\eeprom.n4202 ));
    InMux I__1097 (
            .O(N__12125),
            .I(\eeprom.n4203 ));
    InMux I__1096 (
            .O(N__12122),
            .I(\eeprom.n4204 ));
    InMux I__1095 (
            .O(N__12119),
            .I(\eeprom.n4188 ));
    InMux I__1094 (
            .O(N__12116),
            .I(\eeprom.n4189 ));
    InMux I__1093 (
            .O(N__12113),
            .I(bfn_17_22_0_));
    InMux I__1092 (
            .O(N__12110),
            .I(\eeprom.n4191 ));
    InMux I__1091 (
            .O(N__12107),
            .I(\eeprom.n4192 ));
    InMux I__1090 (
            .O(N__12104),
            .I(\eeprom.n4193 ));
    InMux I__1089 (
            .O(N__12101),
            .I(\eeprom.n4194 ));
    InMux I__1088 (
            .O(N__12098),
            .I(\eeprom.n4195 ));
    InMux I__1087 (
            .O(N__12095),
            .I(\eeprom.n4196 ));
    InMux I__1086 (
            .O(N__12092),
            .I(n3928));
    InMux I__1085 (
            .O(N__12089),
            .I(bfn_17_20_0_));
    InMux I__1084 (
            .O(N__12086),
            .I(n3930));
    InMux I__1083 (
            .O(N__12083),
            .I(N__12080));
    LocalMux I__1082 (
            .O(N__12080),
            .I(N__12077));
    Span4Mux_v I__1081 (
            .O(N__12077),
            .I(N__12073));
    InMux I__1080 (
            .O(N__12076),
            .I(N__12070));
    Odrv4 I__1079 (
            .O(N__12073),
            .I(blink_counter_25));
    LocalMux I__1078 (
            .O(N__12070),
            .I(blink_counter_25));
    InMux I__1077 (
            .O(N__12065),
            .I(bfn_17_21_0_));
    InMux I__1076 (
            .O(N__12062),
            .I(\eeprom.n4183 ));
    InMux I__1075 (
            .O(N__12059),
            .I(\eeprom.n4184 ));
    InMux I__1074 (
            .O(N__12056),
            .I(\eeprom.n4185 ));
    InMux I__1073 (
            .O(N__12053),
            .I(\eeprom.n4186 ));
    InMux I__1072 (
            .O(N__12050),
            .I(\eeprom.n4187 ));
    InMux I__1071 (
            .O(N__12047),
            .I(N__12044));
    LocalMux I__1070 (
            .O(N__12044),
            .I(n12));
    InMux I__1069 (
            .O(N__12041),
            .I(n3919));
    InMux I__1068 (
            .O(N__12038),
            .I(N__12035));
    LocalMux I__1067 (
            .O(N__12035),
            .I(n11_adj_364));
    InMux I__1066 (
            .O(N__12032),
            .I(n3920));
    InMux I__1065 (
            .O(N__12029),
            .I(N__12026));
    LocalMux I__1064 (
            .O(N__12026),
            .I(n10_adj_363));
    InMux I__1063 (
            .O(N__12023),
            .I(bfn_17_19_0_));
    InMux I__1062 (
            .O(N__12020),
            .I(N__12017));
    LocalMux I__1061 (
            .O(N__12017),
            .I(n9));
    InMux I__1060 (
            .O(N__12014),
            .I(n3922));
    InMux I__1059 (
            .O(N__12011),
            .I(N__12008));
    LocalMux I__1058 (
            .O(N__12008),
            .I(n8_adj_362));
    InMux I__1057 (
            .O(N__12005),
            .I(n3923));
    InMux I__1056 (
            .O(N__12002),
            .I(N__11999));
    LocalMux I__1055 (
            .O(N__11999),
            .I(n7));
    InMux I__1054 (
            .O(N__11996),
            .I(n3924));
    InMux I__1053 (
            .O(N__11993),
            .I(N__11990));
    LocalMux I__1052 (
            .O(N__11990),
            .I(n6));
    InMux I__1051 (
            .O(N__11987),
            .I(n3925));
    InMux I__1050 (
            .O(N__11984),
            .I(n3926));
    InMux I__1049 (
            .O(N__11981),
            .I(n3927));
    InMux I__1048 (
            .O(N__11978),
            .I(N__11975));
    LocalMux I__1047 (
            .O(N__11975),
            .I(n20));
    InMux I__1046 (
            .O(N__11972),
            .I(n3911));
    InMux I__1045 (
            .O(N__11969),
            .I(N__11966));
    LocalMux I__1044 (
            .O(N__11966),
            .I(n19));
    InMux I__1043 (
            .O(N__11963),
            .I(n3912));
    InMux I__1042 (
            .O(N__11960),
            .I(N__11957));
    LocalMux I__1041 (
            .O(N__11957),
            .I(n18));
    InMux I__1040 (
            .O(N__11954),
            .I(bfn_17_18_0_));
    InMux I__1039 (
            .O(N__11951),
            .I(N__11948));
    LocalMux I__1038 (
            .O(N__11948),
            .I(n17));
    InMux I__1037 (
            .O(N__11945),
            .I(n3914));
    InMux I__1036 (
            .O(N__11942),
            .I(N__11939));
    LocalMux I__1035 (
            .O(N__11939),
            .I(n16));
    InMux I__1034 (
            .O(N__11936),
            .I(n3915));
    InMux I__1033 (
            .O(N__11933),
            .I(N__11930));
    LocalMux I__1032 (
            .O(N__11930),
            .I(n15));
    InMux I__1031 (
            .O(N__11927),
            .I(n3916));
    InMux I__1030 (
            .O(N__11924),
            .I(N__11921));
    LocalMux I__1029 (
            .O(N__11921),
            .I(n14));
    InMux I__1028 (
            .O(N__11918),
            .I(n3917));
    InMux I__1027 (
            .O(N__11915),
            .I(N__11912));
    LocalMux I__1026 (
            .O(N__11912),
            .I(n13));
    InMux I__1025 (
            .O(N__11909),
            .I(n3918));
    IoInMux I__1024 (
            .O(N__11906),
            .I(N__11903));
    LocalMux I__1023 (
            .O(N__11903),
            .I(N__11900));
    Span4Mux_s2_v I__1022 (
            .O(N__11900),
            .I(N__11897));
    Sp12to4 I__1021 (
            .O(N__11897),
            .I(N__11894));
    Span12Mux_h I__1020 (
            .O(N__11894),
            .I(N__11891));
    Odrv12 I__1019 (
            .O(N__11891),
            .I(LED_c));
    InMux I__1018 (
            .O(N__11888),
            .I(N__11885));
    LocalMux I__1017 (
            .O(N__11885),
            .I(n26));
    InMux I__1016 (
            .O(N__11882),
            .I(bfn_17_17_0_));
    InMux I__1015 (
            .O(N__11879),
            .I(N__11876));
    LocalMux I__1014 (
            .O(N__11876),
            .I(n25));
    InMux I__1013 (
            .O(N__11873),
            .I(n3906));
    InMux I__1012 (
            .O(N__11870),
            .I(N__11867));
    LocalMux I__1011 (
            .O(N__11867),
            .I(n24));
    InMux I__1010 (
            .O(N__11864),
            .I(n3907));
    InMux I__1009 (
            .O(N__11861),
            .I(N__11858));
    LocalMux I__1008 (
            .O(N__11858),
            .I(n23));
    InMux I__1007 (
            .O(N__11855),
            .I(n3908));
    InMux I__1006 (
            .O(N__11852),
            .I(N__11849));
    LocalMux I__1005 (
            .O(N__11849),
            .I(n22));
    InMux I__1004 (
            .O(N__11846),
            .I(n3909));
    InMux I__1003 (
            .O(N__11843),
            .I(N__11840));
    LocalMux I__1002 (
            .O(N__11840),
            .I(n21));
    InMux I__1001 (
            .O(N__11837),
            .I(n3910));
    IoInMux I__1000 (
            .O(N__11834),
            .I(N__11831));
    LocalMux I__999 (
            .O(N__11831),
            .I(N__11828));
    IoSpan4Mux I__998 (
            .O(N__11828),
            .I(N__11825));
    IoSpan4Mux I__997 (
            .O(N__11825),
            .I(N__11822));
    IoSpan4Mux I__996 (
            .O(N__11822),
            .I(N__11819));
    Odrv4 I__995 (
            .O(N__11819),
            .I(CLK_pad_gb_input));
    INV \INVeeprom.i2c.write_enable_132C  (
            .O(\INVeeprom.i2c.write_enable_132C_net ),
            .I(N__29683));
    INV \INVeeprom.i2c.sda_out_133C  (
            .O(\INVeeprom.i2c.sda_out_133C_net ),
            .I(N__29656));
    INV \INVeeprom.i2c.i2c_scl_enable_124C  (
            .O(\INVeeprom.i2c.i2c_scl_enable_124C_net ),
            .I(N__29696));
    defparam IN_MUX_bfv_27_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_27_23_0_));
    defparam IN_MUX_bfv_27_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_24_0_ (
            .carryinitin(\eeprom.n4249 ),
            .carryinitout(bfn_27_24_0_));
    defparam IN_MUX_bfv_27_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_25_0_ (
            .carryinitin(\eeprom.n4257 ),
            .carryinitout(bfn_27_25_0_));
    defparam IN_MUX_bfv_27_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_26_0_ (
            .carryinitin(\eeprom.n4265 ),
            .carryinitout(bfn_27_26_0_));
    defparam IN_MUX_bfv_20_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_17_0_));
    defparam IN_MUX_bfv_20_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_18_0_ (
            .carryinitin(\eeprom.n4235 ),
            .carryinitout(bfn_20_18_0_));
    defparam IN_MUX_bfv_20_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_19_0_));
    defparam IN_MUX_bfv_20_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_20_0_ (
            .carryinitin(\eeprom.n4212 ),
            .carryinitout(bfn_20_20_0_));
    defparam IN_MUX_bfv_20_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_21_0_ (
            .carryinitin(\eeprom.n4220 ),
            .carryinitout(bfn_20_21_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(\eeprom.n4190 ),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(\eeprom.n4198 ),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(\eeprom.n4169 ),
            .carryinitout(bfn_17_25_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(\eeprom.n4177 ),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_17_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_27_0_));
    defparam IN_MUX_bfv_17_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_28_0_ (
            .carryinitin(\eeprom.n4149 ),
            .carryinitout(bfn_17_28_0_));
    defparam IN_MUX_bfv_17_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_29_0_ (
            .carryinitin(\eeprom.n4157 ),
            .carryinitout(bfn_17_29_0_));
    defparam IN_MUX_bfv_19_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_30_0_));
    defparam IN_MUX_bfv_19_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_31_0_ (
            .carryinitin(\eeprom.n4130 ),
            .carryinitout(bfn_19_31_0_));
    defparam IN_MUX_bfv_19_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_32_0_ (
            .carryinitin(\eeprom.n4138 ),
            .carryinitout(bfn_19_32_0_));
    defparam IN_MUX_bfv_18_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_29_0_));
    defparam IN_MUX_bfv_18_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_30_0_ (
            .carryinitin(\eeprom.n4112 ),
            .carryinitout(bfn_18_30_0_));
    defparam IN_MUX_bfv_18_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_31_0_ (
            .carryinitin(\eeprom.n4120 ),
            .carryinitout(bfn_18_31_0_));
    defparam IN_MUX_bfv_20_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_29_0_));
    defparam IN_MUX_bfv_20_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_30_0_ (
            .carryinitin(\eeprom.n4095 ),
            .carryinitout(bfn_20_30_0_));
    defparam IN_MUX_bfv_20_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_31_0_ (
            .carryinitin(\eeprom.n4103 ),
            .carryinitout(bfn_20_31_0_));
    defparam IN_MUX_bfv_21_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_27_0_));
    defparam IN_MUX_bfv_21_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_28_0_ (
            .carryinitin(\eeprom.n4079 ),
            .carryinitout(bfn_21_28_0_));
    defparam IN_MUX_bfv_21_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_29_0_ (
            .carryinitin(\eeprom.n4087 ),
            .carryinitout(bfn_21_29_0_));
    defparam IN_MUX_bfv_22_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_25_0_));
    defparam IN_MUX_bfv_22_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_26_0_ (
            .carryinitin(\eeprom.n4064 ),
            .carryinitout(bfn_22_26_0_));
    defparam IN_MUX_bfv_21_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_23_0_));
    defparam IN_MUX_bfv_21_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_24_0_ (
            .carryinitin(\eeprom.n4050 ),
            .carryinitout(bfn_21_24_0_));
    defparam IN_MUX_bfv_24_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_23_0_));
    defparam IN_MUX_bfv_24_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_24_0_ (
            .carryinitin(\eeprom.n4037 ),
            .carryinitout(bfn_24_24_0_));
    defparam IN_MUX_bfv_22_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_22_0_));
    defparam IN_MUX_bfv_22_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_23_0_ (
            .carryinitin(\eeprom.n4025 ),
            .carryinitout(bfn_22_23_0_));
    defparam IN_MUX_bfv_21_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_20_0_));
    defparam IN_MUX_bfv_21_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_21_0_ (
            .carryinitin(\eeprom.n4014 ),
            .carryinitout(bfn_21_21_0_));
    defparam IN_MUX_bfv_22_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_17_0_));
    defparam IN_MUX_bfv_22_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_18_0_ (
            .carryinitin(\eeprom.n4004 ),
            .carryinitout(bfn_22_18_0_));
    defparam IN_MUX_bfv_24_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_17_0_));
    defparam IN_MUX_bfv_24_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_18_0_ (
            .carryinitin(\eeprom.n3995 ),
            .carryinitout(bfn_24_18_0_));
    defparam IN_MUX_bfv_23_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_18_0_));
    defparam IN_MUX_bfv_23_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_19_0_ (
            .carryinitin(\eeprom.n3987 ),
            .carryinitout(bfn_23_19_0_));
    defparam IN_MUX_bfv_24_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_20_0_));
    defparam IN_MUX_bfv_27_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_27_17_0_));
    defparam IN_MUX_bfv_30_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_30_20_0_));
    defparam IN_MUX_bfv_26_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_21_0_));
    defparam IN_MUX_bfv_26_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_22_0_ (
            .carryinitin(\eeprom.n3938 ),
            .carryinitout(bfn_26_22_0_));
    defparam IN_MUX_bfv_26_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_23_0_ (
            .carryinitin(\eeprom.n3946 ),
            .carryinitout(bfn_26_23_0_));
    defparam IN_MUX_bfv_26_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_24_0_ (
            .carryinitin(\eeprom.n3954 ),
            .carryinitout(bfn_26_24_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_28_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_28_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_28_21_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(n3913),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(n3921),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(n3929),
            .carryinitout(bfn_17_20_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__11834),
            .GLOBALBUFFEROUTPUT(CLK_N));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam i4592_3_lut_LC_15_19_3.C_ON=1'b0;
    defparam i4592_3_lut_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam i4592_3_lut_LC_15_19_3.LUT_INIT=16'b0001000110111011;
    LogicCell40 i4592_3_lut_LC_15_19_3 (
            .in0(N__12083),
            .in1(N__12395),
            .in2(_gnd_net_),
            .in3(N__12311),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i0_LC_17_17_0.C_ON=1'b1;
    defparam blink_counter_227__i0_LC_17_17_0.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i0_LC_17_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i0_LC_17_17_0 (
            .in0(_gnd_net_),
            .in1(N__11888),
            .in2(_gnd_net_),
            .in3(N__11882),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(n3906),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i1_LC_17_17_1.C_ON=1'b1;
    defparam blink_counter_227__i1_LC_17_17_1.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i1_LC_17_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i1_LC_17_17_1 (
            .in0(_gnd_net_),
            .in1(N__11879),
            .in2(_gnd_net_),
            .in3(N__11873),
            .lcout(n25),
            .ltout(),
            .carryin(n3906),
            .carryout(n3907),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i2_LC_17_17_2.C_ON=1'b1;
    defparam blink_counter_227__i2_LC_17_17_2.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i2_LC_17_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i2_LC_17_17_2 (
            .in0(_gnd_net_),
            .in1(N__11870),
            .in2(_gnd_net_),
            .in3(N__11864),
            .lcout(n24),
            .ltout(),
            .carryin(n3907),
            .carryout(n3908),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i3_LC_17_17_3.C_ON=1'b1;
    defparam blink_counter_227__i3_LC_17_17_3.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i3_LC_17_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i3_LC_17_17_3 (
            .in0(_gnd_net_),
            .in1(N__11861),
            .in2(_gnd_net_),
            .in3(N__11855),
            .lcout(n23),
            .ltout(),
            .carryin(n3908),
            .carryout(n3909),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i4_LC_17_17_4.C_ON=1'b1;
    defparam blink_counter_227__i4_LC_17_17_4.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i4_LC_17_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i4_LC_17_17_4 (
            .in0(_gnd_net_),
            .in1(N__11852),
            .in2(_gnd_net_),
            .in3(N__11846),
            .lcout(n22),
            .ltout(),
            .carryin(n3909),
            .carryout(n3910),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i5_LC_17_17_5.C_ON=1'b1;
    defparam blink_counter_227__i5_LC_17_17_5.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i5_LC_17_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i5_LC_17_17_5 (
            .in0(_gnd_net_),
            .in1(N__11843),
            .in2(_gnd_net_),
            .in3(N__11837),
            .lcout(n21),
            .ltout(),
            .carryin(n3910),
            .carryout(n3911),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i6_LC_17_17_6.C_ON=1'b1;
    defparam blink_counter_227__i6_LC_17_17_6.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i6_LC_17_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i6_LC_17_17_6 (
            .in0(_gnd_net_),
            .in1(N__11978),
            .in2(_gnd_net_),
            .in3(N__11972),
            .lcout(n20),
            .ltout(),
            .carryin(n3911),
            .carryout(n3912),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i7_LC_17_17_7.C_ON=1'b1;
    defparam blink_counter_227__i7_LC_17_17_7.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i7_LC_17_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i7_LC_17_17_7 (
            .in0(_gnd_net_),
            .in1(N__11969),
            .in2(_gnd_net_),
            .in3(N__11963),
            .lcout(n19),
            .ltout(),
            .carryin(n3912),
            .carryout(n3913),
            .clk(N__29856),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i8_LC_17_18_0.C_ON=1'b1;
    defparam blink_counter_227__i8_LC_17_18_0.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i8_LC_17_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i8_LC_17_18_0 (
            .in0(_gnd_net_),
            .in1(N__11960),
            .in2(_gnd_net_),
            .in3(N__11954),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(n3914),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i9_LC_17_18_1.C_ON=1'b1;
    defparam blink_counter_227__i9_LC_17_18_1.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i9_LC_17_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i9_LC_17_18_1 (
            .in0(_gnd_net_),
            .in1(N__11951),
            .in2(_gnd_net_),
            .in3(N__11945),
            .lcout(n17),
            .ltout(),
            .carryin(n3914),
            .carryout(n3915),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i10_LC_17_18_2.C_ON=1'b1;
    defparam blink_counter_227__i10_LC_17_18_2.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i10_LC_17_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i10_LC_17_18_2 (
            .in0(_gnd_net_),
            .in1(N__11942),
            .in2(_gnd_net_),
            .in3(N__11936),
            .lcout(n16),
            .ltout(),
            .carryin(n3915),
            .carryout(n3916),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i11_LC_17_18_3.C_ON=1'b1;
    defparam blink_counter_227__i11_LC_17_18_3.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i11_LC_17_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i11_LC_17_18_3 (
            .in0(_gnd_net_),
            .in1(N__11933),
            .in2(_gnd_net_),
            .in3(N__11927),
            .lcout(n15),
            .ltout(),
            .carryin(n3916),
            .carryout(n3917),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i12_LC_17_18_4.C_ON=1'b1;
    defparam blink_counter_227__i12_LC_17_18_4.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i12_LC_17_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i12_LC_17_18_4 (
            .in0(_gnd_net_),
            .in1(N__11924),
            .in2(_gnd_net_),
            .in3(N__11918),
            .lcout(n14),
            .ltout(),
            .carryin(n3917),
            .carryout(n3918),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i13_LC_17_18_5.C_ON=1'b1;
    defparam blink_counter_227__i13_LC_17_18_5.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i13_LC_17_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i13_LC_17_18_5 (
            .in0(_gnd_net_),
            .in1(N__11915),
            .in2(_gnd_net_),
            .in3(N__11909),
            .lcout(n13),
            .ltout(),
            .carryin(n3918),
            .carryout(n3919),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i14_LC_17_18_6.C_ON=1'b1;
    defparam blink_counter_227__i14_LC_17_18_6.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i14_LC_17_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i14_LC_17_18_6 (
            .in0(_gnd_net_),
            .in1(N__12047),
            .in2(_gnd_net_),
            .in3(N__12041),
            .lcout(n12),
            .ltout(),
            .carryin(n3919),
            .carryout(n3920),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i15_LC_17_18_7.C_ON=1'b1;
    defparam blink_counter_227__i15_LC_17_18_7.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i15_LC_17_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i15_LC_17_18_7 (
            .in0(_gnd_net_),
            .in1(N__12038),
            .in2(_gnd_net_),
            .in3(N__12032),
            .lcout(n11_adj_364),
            .ltout(),
            .carryin(n3920),
            .carryout(n3921),
            .clk(N__29857),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i16_LC_17_19_0.C_ON=1'b1;
    defparam blink_counter_227__i16_LC_17_19_0.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i16_LC_17_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i16_LC_17_19_0 (
            .in0(_gnd_net_),
            .in1(N__12029),
            .in2(_gnd_net_),
            .in3(N__12023),
            .lcout(n10_adj_363),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(n3922),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i17_LC_17_19_1.C_ON=1'b1;
    defparam blink_counter_227__i17_LC_17_19_1.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i17_LC_17_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i17_LC_17_19_1 (
            .in0(_gnd_net_),
            .in1(N__12020),
            .in2(_gnd_net_),
            .in3(N__12014),
            .lcout(n9),
            .ltout(),
            .carryin(n3922),
            .carryout(n3923),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i18_LC_17_19_2.C_ON=1'b1;
    defparam blink_counter_227__i18_LC_17_19_2.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i18_LC_17_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i18_LC_17_19_2 (
            .in0(_gnd_net_),
            .in1(N__12011),
            .in2(_gnd_net_),
            .in3(N__12005),
            .lcout(n8_adj_362),
            .ltout(),
            .carryin(n3923),
            .carryout(n3924),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i19_LC_17_19_3.C_ON=1'b1;
    defparam blink_counter_227__i19_LC_17_19_3.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i19_LC_17_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i19_LC_17_19_3 (
            .in0(_gnd_net_),
            .in1(N__12002),
            .in2(_gnd_net_),
            .in3(N__11996),
            .lcout(n7),
            .ltout(),
            .carryin(n3924),
            .carryout(n3925),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i20_LC_17_19_4.C_ON=1'b1;
    defparam blink_counter_227__i20_LC_17_19_4.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i20_LC_17_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i20_LC_17_19_4 (
            .in0(_gnd_net_),
            .in1(N__11993),
            .in2(_gnd_net_),
            .in3(N__11987),
            .lcout(n6),
            .ltout(),
            .carryin(n3925),
            .carryout(n3926),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i21_LC_17_19_5.C_ON=1'b1;
    defparam blink_counter_227__i21_LC_17_19_5.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i21_LC_17_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i21_LC_17_19_5 (
            .in0(_gnd_net_),
            .in1(N__12408),
            .in2(_gnd_net_),
            .in3(N__11984),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n3926),
            .carryout(n3927),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i22_LC_17_19_6.C_ON=1'b1;
    defparam blink_counter_227__i22_LC_17_19_6.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i22_LC_17_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i22_LC_17_19_6 (
            .in0(_gnd_net_),
            .in1(N__12444),
            .in2(_gnd_net_),
            .in3(N__11981),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n3927),
            .carryout(n3928),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i23_LC_17_19_7.C_ON=1'b1;
    defparam blink_counter_227__i23_LC_17_19_7.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i23_LC_17_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i23_LC_17_19_7 (
            .in0(_gnd_net_),
            .in1(N__12423),
            .in2(_gnd_net_),
            .in3(N__12092),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n3928),
            .carryout(n3929),
            .clk(N__29858),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i24_LC_17_20_0.C_ON=1'b1;
    defparam blink_counter_227__i24_LC_17_20_0.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i24_LC_17_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i24_LC_17_20_0 (
            .in0(_gnd_net_),
            .in1(N__12457),
            .in2(_gnd_net_),
            .in3(N__12089),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(n3930),
            .clk(N__29859),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_227__i25_LC_17_20_1.C_ON=1'b0;
    defparam blink_counter_227__i25_LC_17_20_1.SEQ_MODE=4'b1000;
    defparam blink_counter_227__i25_LC_17_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_227__i25_LC_17_20_1 (
            .in0(_gnd_net_),
            .in1(N__12076),
            .in2(_gnd_net_),
            .in3(N__12086),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29859),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_2_lut_LC_17_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_2_lut_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_2_lut_LC_17_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_2_lut_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(N__23421),
            .in2(_gnd_net_),
            .in3(N__12065),
            .lcout(\eeprom.n3486 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\eeprom.n4183 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_3_lut_LC_17_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_3_lut_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_3_lut_LC_17_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_3_lut_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__28538),
            .in2(N__16664),
            .in3(N__12062),
            .lcout(\eeprom.n3485 ),
            .ltout(),
            .carryin(\eeprom.n4183 ),
            .carryout(\eeprom.n4184 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_4_lut_LC_17_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_4_lut_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_4_lut_LC_17_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_4_lut_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16166),
            .in3(N__12059),
            .lcout(\eeprom.n3484 ),
            .ltout(),
            .carryin(\eeprom.n4184 ),
            .carryout(\eeprom.n4185 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_5_lut_LC_17_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_5_lut_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_5_lut_LC_17_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_5_lut_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16625),
            .in3(N__12056),
            .lcout(\eeprom.n3483 ),
            .ltout(),
            .carryin(\eeprom.n4185 ),
            .carryout(\eeprom.n4186 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_6_lut_LC_17_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_6_lut_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_6_lut_LC_17_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_6_lut_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17228),
            .in3(N__12053),
            .lcout(\eeprom.n3482 ),
            .ltout(),
            .carryin(\eeprom.n4186 ),
            .carryout(\eeprom.n4187 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_7_lut_LC_17_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_7_lut_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_7_lut_LC_17_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_7_lut_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(N__16183),
            .in2(_gnd_net_),
            .in3(N__12050),
            .lcout(\eeprom.n3481 ),
            .ltout(),
            .carryin(\eeprom.n4187 ),
            .carryout(\eeprom.n4188 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_8_lut_LC_17_21_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_8_lut_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_8_lut_LC_17_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_8_lut_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16511),
            .in3(N__12119),
            .lcout(\eeprom.n3480 ),
            .ltout(),
            .carryin(\eeprom.n4188 ),
            .carryout(\eeprom.n4189 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_9_lut_LC_17_21_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_9_lut_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_9_lut_LC_17_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_9_lut_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(N__28539),
            .in2(N__12665),
            .in3(N__12116),
            .lcout(\eeprom.n3479 ),
            .ltout(),
            .carryin(\eeprom.n4189 ),
            .carryout(\eeprom.n4190 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_10_lut_LC_17_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_10_lut_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_10_lut_LC_17_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_10_lut_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__28764),
            .in2(N__13759),
            .in3(N__12113),
            .lcout(\eeprom.n3478 ),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\eeprom.n4191 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_11_lut_LC_17_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_11_lut_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_11_lut_LC_17_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_11_lut_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__28768),
            .in2(N__12623),
            .in3(N__12110),
            .lcout(\eeprom.n3477 ),
            .ltout(),
            .carryin(\eeprom.n4191 ),
            .carryout(\eeprom.n4192 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_12_lut_LC_17_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_12_lut_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_12_lut_LC_17_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_12_lut_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(N__28765),
            .in2(N__17033),
            .in3(N__12107),
            .lcout(\eeprom.n3476 ),
            .ltout(),
            .carryin(\eeprom.n4192 ),
            .carryout(\eeprom.n4193 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_13_lut_LC_17_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_13_lut_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_13_lut_LC_17_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_13_lut_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(N__28769),
            .in2(N__13781),
            .in3(N__12104),
            .lcout(\eeprom.n3475 ),
            .ltout(),
            .carryin(\eeprom.n4193 ),
            .carryout(\eeprom.n4194 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_14_lut_LC_17_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_14_lut_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_14_lut_LC_17_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_14_lut_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(N__28766),
            .in2(N__13510),
            .in3(N__12101),
            .lcout(\eeprom.n3474 ),
            .ltout(),
            .carryin(\eeprom.n4194 ),
            .carryout(\eeprom.n4195 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_15_lut_LC_17_22_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_15_lut_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_15_lut_LC_17_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_15_lut_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(N__28770),
            .in2(N__12757),
            .in3(N__12098),
            .lcout(\eeprom.n3473 ),
            .ltout(),
            .carryin(\eeprom.n4195 ),
            .carryout(\eeprom.n4196 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_16_lut_LC_17_22_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_16_lut_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_16_lut_LC_17_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_16_lut_LC_17_22_6  (
            .in0(_gnd_net_),
            .in1(N__28767),
            .in2(N__16751),
            .in3(N__12095),
            .lcout(\eeprom.n3472 ),
            .ltout(),
            .carryin(\eeprom.n4196 ),
            .carryout(\eeprom.n4197 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_17_lut_LC_17_22_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_17_lut_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_17_lut_LC_17_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_17_lut_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(N__28771),
            .in2(N__16710),
            .in3(N__12143),
            .lcout(\eeprom.n3471 ),
            .ltout(),
            .carryin(\eeprom.n4197 ),
            .carryout(\eeprom.n4198 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_18_lut_LC_17_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_18_lut_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_18_lut_LC_17_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_18_lut_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__28772),
            .in2(N__19262),
            .in3(N__12140),
            .lcout(\eeprom.n3470 ),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\eeprom.n4199 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_19_lut_LC_17_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_19_lut_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_19_lut_LC_17_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_19_lut_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__28777),
            .in2(N__14006),
            .in3(N__12137),
            .lcout(\eeprom.n3469 ),
            .ltout(),
            .carryin(\eeprom.n4199 ),
            .carryout(\eeprom.n4200 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_20_lut_LC_17_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_20_lut_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_20_lut_LC_17_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_20_lut_LC_17_23_2  (
            .in0(_gnd_net_),
            .in1(N__14074),
            .in2(N__28874),
            .in3(N__12134),
            .lcout(\eeprom.n3468 ),
            .ltout(),
            .carryin(\eeprom.n4200 ),
            .carryout(\eeprom.n4201 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_21_lut_LC_17_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_21_lut_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_21_lut_LC_17_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_21_lut_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(N__28781),
            .in2(N__14057),
            .in3(N__12131),
            .lcout(\eeprom.n3467 ),
            .ltout(),
            .carryin(\eeprom.n4201 ),
            .carryout(\eeprom.n4202 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_22_lut_LC_17_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_22_lut_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_22_lut_LC_17_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_22_lut_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(N__28773),
            .in2(N__14036),
            .in3(N__12128),
            .lcout(\eeprom.n3466 ),
            .ltout(),
            .carryin(\eeprom.n4202 ),
            .carryout(\eeprom.n4203 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_23_lut_LC_17_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2290_23_lut_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_23_lut_LC_17_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2290_23_lut_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__13818),
            .in2(N__28873),
            .in3(N__12125),
            .lcout(\eeprom.n3465 ),
            .ltout(),
            .carryin(\eeprom.n4203 ),
            .carryout(\eeprom.n4204 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2290_24_lut_LC_17_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2290_24_lut_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2290_24_lut_LC_17_23_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2290_24_lut_LC_17_23_6  (
            .in0(N__28782),
            .in1(N__13798),
            .in2(N__19223),
            .in3(N__12122),
            .lcout(\eeprom.n3496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2232_3_lut_LC_17_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2232_3_lut_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2232_3_lut_LC_17_23_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2232_3_lut_LC_17_23_7  (
            .in0(_gnd_net_),
            .in1(N__14195),
            .in2(N__12194),
            .in3(N__17155),
            .lcout(\eeprom.n3404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_2_lut_LC_17_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_2_lut_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_2_lut_LC_17_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_2_lut_LC_17_24_0  (
            .in0(_gnd_net_),
            .in1(N__22659),
            .in2(_gnd_net_),
            .in3(N__12170),
            .lcout(\eeprom.n3386 ),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(\eeprom.n4162 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_3_lut_LC_17_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_3_lut_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_3_lut_LC_17_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_3_lut_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__28783),
            .in2(N__16880),
            .in3(N__12167),
            .lcout(\eeprom.n3385 ),
            .ltout(),
            .carryin(\eeprom.n4162 ),
            .carryout(\eeprom.n4163 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_4_lut_LC_17_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_4_lut_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_4_lut_LC_17_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_4_lut_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(N__16951),
            .in2(_gnd_net_),
            .in3(N__12164),
            .lcout(\eeprom.n3384 ),
            .ltout(),
            .carryin(\eeprom.n4163 ),
            .carryout(\eeprom.n4164 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_5_lut_LC_17_24_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_5_lut_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_5_lut_LC_17_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_5_lut_LC_17_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16910),
            .in3(N__12161),
            .lcout(\eeprom.n3383 ),
            .ltout(),
            .carryin(\eeprom.n4164 ),
            .carryout(\eeprom.n4165 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_6_lut_LC_17_24_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_6_lut_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_6_lut_LC_17_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_6_lut_LC_17_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17660),
            .in3(N__12158),
            .lcout(\eeprom.n3382 ),
            .ltout(),
            .carryin(\eeprom.n4165 ),
            .carryout(\eeprom.n4166 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_7_lut_LC_17_24_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_7_lut_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_7_lut_LC_17_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_7_lut_LC_17_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16934),
            .in3(N__12155),
            .lcout(\eeprom.n3381 ),
            .ltout(),
            .carryin(\eeprom.n4166 ),
            .carryout(\eeprom.n4167 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_8_lut_LC_17_24_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_8_lut_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_8_lut_LC_17_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_8_lut_LC_17_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16583),
            .in3(N__12152),
            .lcout(\eeprom.n3380 ),
            .ltout(),
            .carryin(\eeprom.n4167 ),
            .carryout(\eeprom.n4168 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_9_lut_LC_17_24_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_9_lut_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_9_lut_LC_17_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_9_lut_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(N__28784),
            .in2(N__13923),
            .in3(N__12149),
            .lcout(\eeprom.n3379 ),
            .ltout(),
            .carryin(\eeprom.n4168 ),
            .carryout(\eeprom.n4169 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_10_lut_LC_17_25_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_10_lut_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_10_lut_LC_17_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_10_lut_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(N__28875),
            .in2(N__13951),
            .in3(N__12146),
            .lcout(\eeprom.n3378 ),
            .ltout(),
            .carryin(bfn_17_25_0_),
            .carryout(\eeprom.n4170 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_11_lut_LC_17_25_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_11_lut_LC_17_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_11_lut_LC_17_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_11_lut_LC_17_25_1  (
            .in0(_gnd_net_),
            .in1(N__28878),
            .in2(N__17180),
            .in3(N__12209),
            .lcout(\eeprom.n3377 ),
            .ltout(),
            .carryin(\eeprom.n4170 ),
            .carryout(\eeprom.n4171 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_12_lut_LC_17_25_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_12_lut_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_12_lut_LC_17_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_12_lut_LC_17_25_2  (
            .in0(_gnd_net_),
            .in1(N__13890),
            .in2(N__28928),
            .in3(N__12206),
            .lcout(\eeprom.n3376 ),
            .ltout(),
            .carryin(\eeprom.n4171 ),
            .carryout(\eeprom.n4172 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_13_lut_LC_17_25_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_13_lut_LC_17_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_13_lut_LC_17_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_13_lut_LC_17_25_3  (
            .in0(_gnd_net_),
            .in1(N__28882),
            .in2(N__14164),
            .in3(N__12203),
            .lcout(\eeprom.n3375 ),
            .ltout(),
            .carryin(\eeprom.n4172 ),
            .carryout(\eeprom.n4173 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_14_lut_LC_17_25_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_14_lut_LC_17_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_14_lut_LC_17_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_14_lut_LC_17_25_4  (
            .in0(_gnd_net_),
            .in1(N__28876),
            .in2(N__13975),
            .in3(N__12200),
            .lcout(\eeprom.n3374 ),
            .ltout(),
            .carryin(\eeprom.n4173 ),
            .carryout(\eeprom.n4174 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_15_lut_LC_17_25_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_15_lut_LC_17_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_15_lut_LC_17_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_15_lut_LC_17_25_5  (
            .in0(_gnd_net_),
            .in1(N__28883),
            .in2(N__14216),
            .in3(N__12197),
            .lcout(\eeprom.n3373 ),
            .ltout(),
            .carryin(\eeprom.n4174 ),
            .carryout(\eeprom.n4175 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_16_lut_LC_17_25_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_16_lut_LC_17_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_16_lut_LC_17_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_16_lut_LC_17_25_6  (
            .in0(_gnd_net_),
            .in1(N__28877),
            .in2(N__14194),
            .in3(N__12182),
            .lcout(\eeprom.n3372 ),
            .ltout(),
            .carryin(\eeprom.n4175 ),
            .carryout(\eeprom.n4176 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_17_lut_LC_17_25_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_17_lut_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_17_lut_LC_17_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_17_lut_LC_17_25_7  (
            .in0(_gnd_net_),
            .in1(N__28884),
            .in2(N__16820),
            .in3(N__12179),
            .lcout(\eeprom.n3371 ),
            .ltout(),
            .carryin(\eeprom.n4176 ),
            .carryout(\eeprom.n4177 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_18_lut_LC_17_26_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_18_lut_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_18_lut_LC_17_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_18_lut_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__28365),
            .in2(N__16847),
            .in3(N__12176),
            .lcout(\eeprom.n3370 ),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(\eeprom.n4178 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_19_lut_LC_17_26_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_19_lut_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_19_lut_LC_17_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_19_lut_LC_17_26_1  (
            .in0(_gnd_net_),
            .in1(N__28885),
            .in2(N__16785),
            .in3(N__12173),
            .lcout(\eeprom.n3369 ),
            .ltout(),
            .carryin(\eeprom.n4178 ),
            .carryout(\eeprom.n4179 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_20_lut_LC_17_26_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_20_lut_LC_17_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_20_lut_LC_17_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_20_lut_LC_17_26_2  (
            .in0(_gnd_net_),
            .in1(N__28366),
            .in2(N__12803),
            .in3(N__12236),
            .lcout(\eeprom.n3368 ),
            .ltout(),
            .carryin(\eeprom.n4179 ),
            .carryout(\eeprom.n4180 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_21_lut_LC_17_26_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_21_lut_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_21_lut_LC_17_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_21_lut_LC_17_26_3  (
            .in0(_gnd_net_),
            .in1(N__12710),
            .in2(N__28543),
            .in3(N__12233),
            .lcout(\eeprom.n3367 ),
            .ltout(),
            .carryin(\eeprom.n4180 ),
            .carryout(\eeprom.n4181 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_22_lut_LC_17_26_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2223_22_lut_LC_17_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_22_lut_LC_17_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2223_22_lut_LC_17_26_4  (
            .in0(_gnd_net_),
            .in1(N__12845),
            .in2(N__28929),
            .in3(N__12230),
            .lcout(\eeprom.n3366 ),
            .ltout(),
            .carryin(\eeprom.n4181 ),
            .carryout(\eeprom.n4182 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2223_23_lut_LC_17_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2223_23_lut_LC_17_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2223_23_lut_LC_17_26_5 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \eeprom.rem_4_add_2223_23_lut_LC_17_26_5  (
            .in0(N__28370),
            .in1(N__17159),
            .in2(N__12872),
            .in3(N__12227),
            .lcout(\eeprom.n3397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2169_3_lut_LC_17_26_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2169_3_lut_LC_17_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2169_3_lut_LC_17_26_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2169_3_lut_LC_17_26_7  (
            .in0(_gnd_net_),
            .in1(N__18186),
            .in2(N__12263),
            .in3(N__17782),
            .lcout(\eeprom.n3309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_2_lut_LC_17_27_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_2_lut_LC_17_27_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_2_lut_LC_17_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_2_lut_LC_17_27_0  (
            .in0(_gnd_net_),
            .in1(N__24231),
            .in2(_gnd_net_),
            .in3(N__12224),
            .lcout(\eeprom.n3286 ),
            .ltout(),
            .carryin(bfn_17_27_0_),
            .carryout(\eeprom.n4142 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_3_lut_LC_17_27_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_3_lut_LC_17_27_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_3_lut_LC_17_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_3_lut_LC_17_27_1  (
            .in0(_gnd_net_),
            .in1(N__28371),
            .in2(N__16989),
            .in3(N__12221),
            .lcout(\eeprom.n3285 ),
            .ltout(),
            .carryin(\eeprom.n4142 ),
            .carryout(\eeprom.n4143 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_4_lut_LC_17_27_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_4_lut_LC_17_27_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_4_lut_LC_17_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_4_lut_LC_17_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17327),
            .in3(N__12218),
            .lcout(\eeprom.n3284 ),
            .ltout(),
            .carryin(\eeprom.n4143 ),
            .carryout(\eeprom.n4144 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_5_lut_LC_17_27_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_5_lut_LC_17_27_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_5_lut_LC_17_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_5_lut_LC_17_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17495),
            .in3(N__12215),
            .lcout(\eeprom.n3283 ),
            .ltout(),
            .carryin(\eeprom.n4144 ),
            .carryout(\eeprom.n4145 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_6_lut_LC_17_27_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_6_lut_LC_17_27_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_6_lut_LC_17_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_6_lut_LC_17_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17402),
            .in3(N__12212),
            .lcout(\eeprom.n3282 ),
            .ltout(),
            .carryin(\eeprom.n4145 ),
            .carryout(\eeprom.n4146 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_7_lut_LC_17_27_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_7_lut_LC_17_27_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_7_lut_LC_17_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_7_lut_LC_17_27_5  (
            .in0(_gnd_net_),
            .in1(N__17513),
            .in2(_gnd_net_),
            .in3(N__12275),
            .lcout(\eeprom.n3281 ),
            .ltout(),
            .carryin(\eeprom.n4146 ),
            .carryout(\eeprom.n4147 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_8_lut_LC_17_27_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_8_lut_LC_17_27_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_8_lut_LC_17_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_8_lut_LC_17_27_6  (
            .in0(_gnd_net_),
            .in1(N__17584),
            .in2(_gnd_net_),
            .in3(N__12272),
            .lcout(\eeprom.n3280 ),
            .ltout(),
            .carryin(\eeprom.n4147 ),
            .carryout(\eeprom.n4148 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_9_lut_LC_17_27_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_9_lut_LC_17_27_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_9_lut_LC_17_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_9_lut_LC_17_27_7  (
            .in0(_gnd_net_),
            .in1(N__14259),
            .in2(N__28544),
            .in3(N__12269),
            .lcout(\eeprom.n3279 ),
            .ltout(),
            .carryin(\eeprom.n4148 ),
            .carryout(\eeprom.n4149 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_10_lut_LC_17_28_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_10_lut_LC_17_28_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_10_lut_LC_17_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_10_lut_LC_17_28_0  (
            .in0(_gnd_net_),
            .in1(N__18224),
            .in2(N__28930),
            .in3(N__12266),
            .lcout(\eeprom.n3278 ),
            .ltout(),
            .carryin(bfn_17_28_0_),
            .carryout(\eeprom.n4150 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_11_lut_LC_17_28_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_11_lut_LC_17_28_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_11_lut_LC_17_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_11_lut_LC_17_28_1  (
            .in0(_gnd_net_),
            .in1(N__28892),
            .in2(N__18194),
            .in3(N__12251),
            .lcout(\eeprom.n3277 ),
            .ltout(),
            .carryin(\eeprom.n4150 ),
            .carryout(\eeprom.n4151 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_12_lut_LC_17_28_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_12_lut_LC_17_28_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_12_lut_LC_17_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_12_lut_LC_17_28_2  (
            .in0(_gnd_net_),
            .in1(N__28375),
            .in2(N__17836),
            .in3(N__12248),
            .lcout(\eeprom.n3276 ),
            .ltout(),
            .carryin(\eeprom.n4151 ),
            .carryout(\eeprom.n4152 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_13_lut_LC_17_28_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_13_lut_LC_17_28_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_13_lut_LC_17_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_13_lut_LC_17_28_3  (
            .in0(_gnd_net_),
            .in1(N__17251),
            .in2(N__28545),
            .in3(N__12245),
            .lcout(\eeprom.n3275 ),
            .ltout(),
            .carryin(\eeprom.n4152 ),
            .carryout(\eeprom.n4153 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_14_lut_LC_17_28_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_14_lut_LC_17_28_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_14_lut_LC_17_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_14_lut_LC_17_28_4  (
            .in0(_gnd_net_),
            .in1(N__28379),
            .in2(N__14366),
            .in3(N__12242),
            .lcout(\eeprom.n3274 ),
            .ltout(),
            .carryin(\eeprom.n4153 ),
            .carryout(\eeprom.n4154 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_15_lut_LC_17_28_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_15_lut_LC_17_28_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_15_lut_LC_17_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_15_lut_LC_17_28_5  (
            .in0(_gnd_net_),
            .in1(N__14288),
            .in2(N__28546),
            .in3(N__12239),
            .lcout(\eeprom.n3273 ),
            .ltout(),
            .carryin(\eeprom.n4154 ),
            .carryout(\eeprom.n4155 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_16_lut_LC_17_28_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_16_lut_LC_17_28_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_16_lut_LC_17_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_16_lut_LC_17_28_6  (
            .in0(_gnd_net_),
            .in1(N__14426),
            .in2(N__28931),
            .in3(N__12299),
            .lcout(\eeprom.n3272 ),
            .ltout(),
            .carryin(\eeprom.n4155 ),
            .carryout(\eeprom.n4156 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_17_lut_LC_17_28_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_17_lut_LC_17_28_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_17_lut_LC_17_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_17_lut_LC_17_28_7  (
            .in0(_gnd_net_),
            .in1(N__14393),
            .in2(N__28547),
            .in3(N__12296),
            .lcout(\eeprom.n3271 ),
            .ltout(),
            .carryin(\eeprom.n4156 ),
            .carryout(\eeprom.n4157 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_18_lut_LC_17_29_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_18_lut_LC_17_29_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_18_lut_LC_17_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_18_lut_LC_17_29_0  (
            .in0(_gnd_net_),
            .in1(N__28386),
            .in2(N__12995),
            .in3(N__12293),
            .lcout(\eeprom.n3270 ),
            .ltout(),
            .carryin(bfn_17_29_0_),
            .carryout(\eeprom.n4158 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_19_lut_LC_17_29_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_19_lut_LC_17_29_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_19_lut_LC_17_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_19_lut_LC_17_29_1  (
            .in0(_gnd_net_),
            .in1(N__13048),
            .in2(N__28548),
            .in3(N__12290),
            .lcout(\eeprom.n3269 ),
            .ltout(),
            .carryin(\eeprom.n4158 ),
            .carryout(\eeprom.n4159 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_20_lut_LC_17_29_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_20_lut_LC_17_29_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_20_lut_LC_17_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_20_lut_LC_17_29_2  (
            .in0(_gnd_net_),
            .in1(N__28390),
            .in2(N__13022),
            .in3(N__12287),
            .lcout(\eeprom.n3268 ),
            .ltout(),
            .carryin(\eeprom.n4159 ),
            .carryout(\eeprom.n4160 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_21_lut_LC_17_29_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2156_21_lut_LC_17_29_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_21_lut_LC_17_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2156_21_lut_LC_17_29_3  (
            .in0(_gnd_net_),
            .in1(N__28391),
            .in2(N__12977),
            .in3(N__12284),
            .lcout(\eeprom.n3267 ),
            .ltout(),
            .carryin(\eeprom.n4160 ),
            .carryout(\eeprom.n4161 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2156_22_lut_LC_17_29_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2156_22_lut_LC_17_29_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2156_22_lut_LC_17_29_4 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2156_22_lut_LC_17_29_4  (
            .in0(N__28392),
            .in1(N__15082),
            .in2(N__17786),
            .in3(N__12281),
            .lcout(\eeprom.n3298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1960_3_lut_LC_17_30_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1960_3_lut_LC_17_30_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1960_3_lut_LC_17_30_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1960_3_lut_LC_17_30_0  (
            .in0(_gnd_net_),
            .in1(N__19748),
            .in2(N__18824),
            .in3(N__18779),
            .lcout(\eeprom.n3004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_2_lut_LC_18_17_0 .C_ON=1'b1;
    defparam \eeprom.add_823_2_lut_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_2_lut_LC_18_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_823_2_lut_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__21577),
            .in2(_gnd_net_),
            .in3(N__12278),
            .lcout(\eeprom.n1208 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\eeprom.n3966 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_3_lut_LC_18_17_1 .C_ON=1'b1;
    defparam \eeprom.add_823_3_lut_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_3_lut_LC_18_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_823_3_lut_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__13378),
            .in2(N__28537),
            .in3(N__12332),
            .lcout(\eeprom.n1207 ),
            .ltout(),
            .carryin(\eeprom.n3966 ),
            .carryout(\eeprom.n3967 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_4_lut_LC_18_17_2 .C_ON=1'b1;
    defparam \eeprom.add_823_4_lut_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_4_lut_LC_18_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_823_4_lut_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13568),
            .in3(N__12329),
            .lcout(\eeprom.n1206 ),
            .ltout(),
            .carryin(\eeprom.n3967 ),
            .carryout(\eeprom.n3968 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_5_lut_LC_18_17_3 .C_ON=1'b1;
    defparam \eeprom.add_823_5_lut_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_5_lut_LC_18_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_823_5_lut_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13340),
            .in3(N__12326),
            .lcout(\eeprom.n1205 ),
            .ltout(),
            .carryin(\eeprom.n3968 ),
            .carryout(\eeprom.n3969 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_6_lut_LC_18_17_4 .C_ON=1'b1;
    defparam \eeprom.add_823_6_lut_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_6_lut_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_823_6_lut_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__13478),
            .in2(_gnd_net_),
            .in3(N__12323),
            .lcout(\eeprom.n1204 ),
            .ltout(),
            .carryin(\eeprom.n3969 ),
            .carryout(\eeprom.n3970 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_7_lut_LC_18_17_5 .C_ON=1'b1;
    defparam \eeprom.add_823_7_lut_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_7_lut_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_823_7_lut_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12356),
            .in3(N__12320),
            .lcout(\eeprom.n1203 ),
            .ltout(),
            .carryin(\eeprom.n3970 ),
            .carryout(\eeprom.n3971 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_8_lut_LC_18_17_6 .C_ON=1'b1;
    defparam \eeprom.add_823_8_lut_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_8_lut_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_823_8_lut_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__13225),
            .in2(_gnd_net_),
            .in3(N__12317),
            .lcout(\eeprom.n1202 ),
            .ltout(),
            .carryin(\eeprom.n3971 ),
            .carryout(\eeprom.n3972 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_823_9_lut_LC_18_17_7 .C_ON=1'b0;
    defparam \eeprom.add_823_9_lut_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_823_9_lut_LC_18_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \eeprom.add_823_9_lut_LC_18_17_7  (
            .in0(N__28356),
            .in1(N__13583),
            .in2(_gnd_net_),
            .in3(N__12314),
            .lcout(\eeprom.n1201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4591_4_lut_LC_18_18_1.C_ON=1'b0;
    defparam i4591_4_lut_LC_18_18_1.SEQ_MODE=4'b0000;
    defparam i4591_4_lut_LC_18_18_1.LUT_INIT=16'b1111111010110000;
    LogicCell40 i4591_4_lut_LC_18_18_1 (
            .in0(N__12464),
            .in1(N__12446),
            .in2(N__12431),
            .in3(N__12410),
            .lcout(n5421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4738_1_lut_2_lut_LC_18_18_2 .C_ON=1'b0;
    defparam \eeprom.i4738_1_lut_2_lut_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4738_1_lut_2_lut_LC_18_18_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i4738_1_lut_2_lut_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13451),
            .in3(N__13435),
            .lcout(\eeprom.n5568 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4590_4_lut_LC_18_18_3.C_ON=1'b0;
    defparam i4590_4_lut_LC_18_18_3.SEQ_MODE=4'b0000;
    defparam i4590_4_lut_LC_18_18_3.LUT_INIT=16'b1101110101000000;
    LogicCell40 i4590_4_lut_LC_18_18_3 (
            .in0(N__12463),
            .in1(N__12445),
            .in2(N__12430),
            .in3(N__12409),
            .lcout(n5420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2445_3_lut_LC_18_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2445_3_lut_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2445_3_lut_LC_18_18_4 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \eeprom.rem_4_i2445_3_lut_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__12352),
            .in2(N__12383),
            .in3(N__13434),
            .lcout(\eeprom.n3713 ),
            .ltout(\eeprom.n3713_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4732_1_lut_LC_18_18_5 .C_ON=1'b0;
    defparam \eeprom.i4732_1_lut_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4732_1_lut_LC_18_18_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4732_1_lut_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12374),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2382_3_lut_LC_18_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2382_3_lut_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2382_3_lut_LC_18_18_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i2382_3_lut_LC_18_18_6  (
            .in0(N__15485),
            .in1(N__29459),
            .in2(_gnd_net_),
            .in3(N__16328),
            .lcout(\eeprom.n3618 ),
            .ltout(\eeprom.n3618_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_100_LC_18_18_7 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_100_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_100_LC_18_18_7 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \eeprom.i1_4_lut_adj_100_LC_18_18_7  (
            .in0(N__21576),
            .in1(N__12509),
            .in2(N__12371),
            .in3(N__12362),
            .lcout(\eeprom.n5017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2379_3_lut_LC_18_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2379_3_lut_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2379_3_lut_LC_18_19_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2379_3_lut_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__15854),
            .in2(N__16323),
            .in3(N__15880),
            .lcout(\eeprom.n3615 ),
            .ltout(\eeprom.n3615_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_89_LC_18_19_1 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_89_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_89_LC_18_19_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_89_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12368),
            .in3(N__13218),
            .lcout(),
            .ltout(\eeprom.n5221_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_99_LC_18_19_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_99_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_99_LC_18_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_99_LC_18_19_2  (
            .in0(N__12348),
            .in1(N__13557),
            .in2(N__12365),
            .in3(N__13329),
            .lcout(\eeprom.n5225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2378_3_lut_LC_18_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2378_3_lut_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2378_3_lut_LC_18_19_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2378_3_lut_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__15841),
            .in2(N__15815),
            .in3(N__16300),
            .lcout(\eeprom.n3614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2369_3_lut_LC_18_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2369_3_lut_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2369_3_lut_LC_18_19_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2369_3_lut_LC_18_19_4  (
            .in0(N__16064),
            .in1(_gnd_net_),
            .in2(N__16324),
            .in3(N__16046),
            .lcout(\eeprom.n3605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2380_3_lut_LC_18_19_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2380_3_lut_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2380_3_lut_LC_18_19_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2380_3_lut_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__15436),
            .in2(N__15410),
            .in3(N__16301),
            .lcout(\eeprom.n3616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2299_3_lut_LC_18_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2299_3_lut_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2299_3_lut_LC_18_19_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2299_3_lut_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__16715),
            .in2(N__12503),
            .in3(N__19221),
            .lcout(\eeprom.n3503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i14_3_lut_LC_18_20_0 .C_ON=1'b0;
    defparam \eeprom.i14_3_lut_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i14_3_lut_LC_18_20_0 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \eeprom.i14_3_lut_LC_18_20_0  (
            .in0(N__16129),
            .in1(_gnd_net_),
            .in2(N__13694),
            .in3(N__16062),
            .lcout(),
            .ltout(\eeprom.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i17_4_lut_LC_18_20_1 .C_ON=1'b0;
    defparam \eeprom.i17_4_lut_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i17_4_lut_LC_18_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i17_4_lut_LC_18_20_1  (
            .in0(N__12542),
            .in1(N__12578),
            .in2(N__12488),
            .in3(N__13589),
            .lcout(\eeprom.n3529 ),
            .ltout(\eeprom.n3529_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2377_3_lut_LC_18_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2377_3_lut_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2377_3_lut_LC_18_20_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2377_3_lut_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__15793),
            .in2(N__12485),
            .in3(N__15779),
            .lcout(\eeprom.n3613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2309_3_lut_LC_18_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2309_3_lut_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2309_3_lut_LC_18_20_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2309_3_lut_LC_18_20_4  (
            .in0(N__12482),
            .in1(_gnd_net_),
            .in2(N__16187),
            .in3(N__19194),
            .lcout(\eeprom.n3513 ),
            .ltout(\eeprom.n3513_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_19_LC_18_20_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_19_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_19_LC_18_20_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_19_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12476),
            .in3(N__15831),
            .lcout(\eeprom.n5321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2301_3_lut_LC_18_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2301_3_lut_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2301_3_lut_LC_18_20_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2301_3_lut_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__12473),
            .in2(N__12764),
            .in3(N__19195),
            .lcout(\eeprom.n3505 ),
            .ltout(\eeprom.n3505_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_22_LC_18_20_7 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_22_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_22_LC_18_20_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_22_LC_18_20_7  (
            .in0(N__15727),
            .in1(N__15993),
            .in2(N__12581),
            .in3(N__12515),
            .lcout(\eeprom.n30_adj_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4682_3_lut_LC_18_21_0 .C_ON=1'b0;
    defparam \eeprom.i4682_3_lut_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4682_3_lut_LC_18_21_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.i4682_3_lut_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__12572),
            .in2(N__19206),
            .in3(N__13760),
            .lcout(\eeprom.n3510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2300_3_lut_LC_18_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2300_3_lut_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2300_3_lut_LC_18_21_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2300_3_lut_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__12566),
            .in2(N__16750),
            .in3(N__19172),
            .lcout(\eeprom.n3504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2312_3_lut_LC_18_21_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2312_3_lut_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2312_3_lut_LC_18_21_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2312_3_lut_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__16165),
            .in2(N__19205),
            .in3(N__12560),
            .lcout(\eeprom.n3516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2303_3_lut_LC_18_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2303_3_lut_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2303_3_lut_LC_18_21_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2303_3_lut_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(N__13780),
            .in2(N__12554),
            .in3(N__19173),
            .lcout(\eeprom.n3507 ),
            .ltout(\eeprom.n3507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_adj_23_LC_18_21_4 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_adj_23_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_adj_23_LC_18_21_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_adj_23_LC_18_21_4  (
            .in0(N__15690),
            .in1(N__15609),
            .in2(N__12545),
            .in3(N__15654),
            .lcout(\eeprom.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2310_3_lut_LC_18_21_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2310_3_lut_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2310_3_lut_LC_18_21_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2310_3_lut_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(N__17227),
            .in2(N__12536),
            .in3(N__19168),
            .lcout(\eeprom.n3514 ),
            .ltout(\eeprom.n3514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_20_LC_18_21_6 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_20_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_20_LC_18_21_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_20_LC_18_21_6  (
            .in0(N__15870),
            .in1(_gnd_net_),
            .in2(N__12527),
            .in3(N__15426),
            .lcout(),
            .ltout(\eeprom.n5323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_21_LC_18_21_7 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_21_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_21_LC_18_21_7 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_21_LC_18_21_7  (
            .in0(N__29457),
            .in1(N__15465),
            .in2(N__12524),
            .in3(N__12521),
            .lcout(\eeprom.n4753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_LC_18_22_0 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_LC_18_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_LC_18_22_0  (
            .in0(N__12664),
            .in1(N__12750),
            .in2(N__13509),
            .in3(N__12622),
            .lcout(\eeprom.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2236_3_lut_LC_18_22_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2236_3_lut_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2236_3_lut_LC_18_22_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2236_3_lut_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__13898),
            .in2(N__17157),
            .in3(N__12692),
            .lcout(\eeprom.n3408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2240_3_lut_LC_18_22_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2240_3_lut_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2240_3_lut_LC_18_22_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2240_3_lut_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__16582),
            .in2(N__12680),
            .in3(N__17132),
            .lcout(\eeprom.n3412 ),
            .ltout(\eeprom.n3412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2307_3_lut_LC_18_22_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2307_3_lut_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2307_3_lut_LC_18_22_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2307_3_lut_LC_18_22_3  (
            .in0(N__19188),
            .in1(_gnd_net_),
            .in2(N__12650),
            .in3(N__12647),
            .lcout(\eeprom.n3511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2235_3_lut_LC_18_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2235_3_lut_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2235_3_lut_LC_18_22_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2235_3_lut_LC_18_22_4  (
            .in0(N__12641),
            .in1(_gnd_net_),
            .in2(N__14168),
            .in3(N__17136),
            .lcout(\eeprom.n3407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2238_3_lut_LC_18_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2238_3_lut_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2238_3_lut_LC_18_22_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2238_3_lut_LC_18_22_5  (
            .in0(N__12632),
            .in1(_gnd_net_),
            .in2(N__17156),
            .in3(N__13952),
            .lcout(\eeprom.n3410 ),
            .ltout(\eeprom.n3410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2305_3_lut_LC_18_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2305_3_lut_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2305_3_lut_LC_18_22_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2305_3_lut_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(N__12608),
            .in2(N__12602),
            .in3(N__19189),
            .lcout(\eeprom.n3509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2293_3_lut_LC_18_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2293_3_lut_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2293_3_lut_LC_18_22_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2293_3_lut_LC_18_22_7  (
            .in0(N__13819),
            .in1(_gnd_net_),
            .in2(N__19215),
            .in3(N__12599),
            .lcout(\eeprom.n3497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2227_3_lut_LC_18_23_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2227_3_lut_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2227_3_lut_LC_18_23_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2227_3_lut_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(N__12706),
            .in2(N__17158),
            .in3(N__12593),
            .lcout(\eeprom.n3399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2159_3_lut_LC_18_23_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2159_3_lut_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2159_3_lut_LC_18_23_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2159_3_lut_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(N__12887),
            .in2(N__12973),
            .in3(N__17764),
            .lcout(\eeprom.n3299 ),
            .ltout(\eeprom.n3299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_LC_18_23_2 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_LC_18_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_LC_18_23_2  (
            .in0(N__12796),
            .in1(N__12705),
            .in2(N__12875),
            .in3(N__12871),
            .lcout(\eeprom.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4681_3_lut_LC_18_23_3 .C_ON=1'b0;
    defparam \eeprom.i4681_3_lut_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4681_3_lut_LC_18_23_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.i4681_3_lut_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__12851),
            .in2(N__13925),
            .in3(N__17140),
            .lcout(\eeprom.n3411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2226_3_lut_LC_18_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2226_3_lut_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2226_3_lut_LC_18_23_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2226_3_lut_LC_18_23_4  (
            .in0(N__17146),
            .in1(_gnd_net_),
            .in2(N__12844),
            .in3(N__12824),
            .lcout(\eeprom.n3398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2161_3_lut_LC_18_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2161_3_lut_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2161_3_lut_LC_18_23_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2161_3_lut_LC_18_23_5  (
            .in0(N__12815),
            .in1(_gnd_net_),
            .in2(N__13052),
            .in3(N__17763),
            .lcout(\eeprom.n3301 ),
            .ltout(\eeprom.n3301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2228_3_lut_LC_18_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2228_3_lut_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2228_3_lut_LC_18_23_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2228_3_lut_LC_18_23_6  (
            .in0(N__17145),
            .in1(_gnd_net_),
            .in2(N__12785),
            .in3(N__12782),
            .lcout(\eeprom.n3400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2234_3_lut_LC_18_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2234_3_lut_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2234_3_lut_LC_18_23_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2234_3_lut_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__12773),
            .in2(N__13976),
            .in3(N__17141),
            .lcout(\eeprom.n3406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2230_3_lut_LC_18_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2230_3_lut_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2230_3_lut_LC_18_24_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2230_3_lut_LC_18_24_0  (
            .in0(_gnd_net_),
            .in1(N__16840),
            .in2(N__12734),
            .in3(N__17149),
            .lcout(\eeprom.n3402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2160_3_lut_LC_18_24_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2160_3_lut_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2160_3_lut_LC_18_24_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2160_3_lut_LC_18_24_1  (
            .in0(_gnd_net_),
            .in1(N__12722),
            .in2(N__17775),
            .in3(N__13021),
            .lcout(\eeprom.n3300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2092_3_lut_LC_18_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2092_3_lut_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2092_3_lut_LC_18_24_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2092_3_lut_LC_18_24_2  (
            .in0(_gnd_net_),
            .in1(N__15151),
            .in2(N__15125),
            .in3(N__17947),
            .lcout(\eeprom.n3200 ),
            .ltout(\eeprom.n3200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_38_LC_18_24_3 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_38_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_38_LC_18_24_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_adj_38_LC_18_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12953),
            .in3(N__15083),
            .lcout(\eeprom.n16_adj_303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2178_3_lut_LC_18_24_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2178_3_lut_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2178_3_lut_LC_18_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i2178_3_lut_LC_18_24_4  (
            .in0(N__12950),
            .in1(N__24235),
            .in2(_gnd_net_),
            .in3(N__17744),
            .lcout(\eeprom.n3318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2172_rep_14_3_lut_LC_18_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2172_rep_14_3_lut_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2172_rep_14_3_lut_LC_18_24_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2172_rep_14_3_lut_LC_18_24_5  (
            .in0(_gnd_net_),
            .in1(N__12938),
            .in2(N__17774),
            .in3(N__17585),
            .lcout(\eeprom.n3312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2167_3_lut_LC_18_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2167_3_lut_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2167_3_lut_LC_18_24_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2167_3_lut_LC_18_24_7  (
            .in0(N__17252),
            .in1(_gnd_net_),
            .in2(N__17776),
            .in3(N__12926),
            .lcout(\eeprom.n3307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2168_3_lut_LC_18_25_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2168_3_lut_LC_18_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2168_3_lut_LC_18_25_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2168_3_lut_LC_18_25_0  (
            .in0(_gnd_net_),
            .in1(N__17837),
            .in2(N__17777),
            .in3(N__12914),
            .lcout(\eeprom.n3308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2171_3_lut_LC_18_25_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2171_3_lut_LC_18_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2171_3_lut_LC_18_25_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2171_3_lut_LC_18_25_1  (
            .in0(_gnd_net_),
            .in1(N__12902),
            .in2(N__14264),
            .in3(N__17758),
            .lcout(\eeprom.n3311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2096_3_lut_LC_18_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2096_3_lut_LC_18_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2096_3_lut_LC_18_25_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2096_3_lut_LC_18_25_2  (
            .in0(_gnd_net_),
            .in1(N__15290),
            .in2(N__15323),
            .in3(N__17946),
            .lcout(\eeprom.n3204 ),
            .ltout(\eeprom.n3204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_adj_39_LC_18_25_3 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_adj_39_LC_18_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_adj_39_LC_18_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_adj_39_LC_18_25_3  (
            .in0(N__12988),
            .in1(N__13035),
            .in2(N__12890),
            .in3(N__13011),
            .lcout(\eeprom.n24_adj_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2098_3_lut_LC_18_25_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2098_3_lut_LC_18_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2098_3_lut_LC_18_25_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \eeprom.rem_4_i2098_3_lut_LC_18_25_4  (
            .in0(_gnd_net_),
            .in1(N__17945),
            .in2(N__14915),
            .in3(N__14891),
            .lcout(\eeprom.n3206 ),
            .ltout(\eeprom.n3206_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2165_3_lut_LC_18_25_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2165_3_lut_LC_18_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2165_3_lut_LC_18_25_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2165_3_lut_LC_18_25_5  (
            .in0(_gnd_net_),
            .in1(N__13067),
            .in2(N__13058),
            .in3(N__17754),
            .lcout(\eeprom.n3305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2032_3_lut_LC_18_25_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2032_3_lut_LC_18_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2032_3_lut_LC_18_25_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2032_3_lut_LC_18_25_6  (
            .in0(_gnd_net_),
            .in1(N__13139),
            .in2(N__14314),
            .in3(N__18146),
            .lcout(\eeprom.n3108 ),
            .ltout(\eeprom.n3108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_LC_18_25_7 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_LC_18_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_LC_18_25_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_LC_18_25_7  (
            .in0(N__17292),
            .in1(N__14997),
            .in2(N__13055),
            .in3(N__14910),
            .lcout(\eeprom.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i8_4_lut_LC_18_26_0 .C_ON=1'b0;
    defparam \eeprom.i8_4_lut_LC_18_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i8_4_lut_LC_18_26_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i8_4_lut_LC_18_26_0  (
            .in0(N__15183),
            .in1(N__15141),
            .in2(N__15104),
            .in3(N__15226),
            .lcout(\eeprom.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2094_3_lut_LC_18_26_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2094_3_lut_LC_18_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2094_3_lut_LC_18_26_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \eeprom.rem_4_i2094_3_lut_LC_18_26_2  (
            .in0(_gnd_net_),
            .in1(N__17933),
            .in2(N__15230),
            .in3(N__15206),
            .lcout(\eeprom.n3202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2093_3_lut_LC_18_26_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2093_3_lut_LC_18_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2093_3_lut_LC_18_26_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \eeprom.rem_4_i2093_3_lut_LC_18_26_3  (
            .in0(N__17934),
            .in1(_gnd_net_),
            .in2(N__15170),
            .in3(N__15184),
            .lcout(\eeprom.n3201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2110_3_lut_LC_18_26_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2110_3_lut_LC_18_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2110_3_lut_LC_18_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i2110_3_lut_LC_18_26_4  (
            .in0(N__14795),
            .in1(N__22407),
            .in2(_gnd_net_),
            .in3(N__17926),
            .lcout(\eeprom.n3218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2095_3_lut_LC_18_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2095_3_lut_LC_18_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2095_3_lut_LC_18_26_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2095_3_lut_LC_18_26_5  (
            .in0(_gnd_net_),
            .in1(N__15245),
            .in2(N__17953),
            .in3(N__15275),
            .lcout(\eeprom.n3203 ),
            .ltout(\eeprom.n3203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2162_3_lut_LC_18_26_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2162_3_lut_LC_18_26_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2162_3_lut_LC_18_26_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2162_3_lut_LC_18_26_6  (
            .in0(_gnd_net_),
            .in1(N__13085),
            .in2(N__13076),
            .in3(N__17772),
            .lcout(\eeprom.n3302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2102_3_lut_LC_18_26_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2102_3_lut_LC_18_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2102_3_lut_LC_18_26_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2102_3_lut_LC_18_26_7  (
            .in0(_gnd_net_),
            .in1(N__14998),
            .in2(N__17952),
            .in3(N__14975),
            .lcout(\eeprom.n3210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2025_3_lut_LC_18_27_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2025_3_lut_LC_18_27_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2025_3_lut_LC_18_27_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2025_3_lut_LC_18_27_0  (
            .in0(_gnd_net_),
            .in1(N__14560),
            .in2(N__13277),
            .in3(N__18124),
            .lcout(\eeprom.n3101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2104_3_lut_LC_18_27_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2104_3_lut_LC_18_27_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2104_3_lut_LC_18_27_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2104_3_lut_LC_18_27_1  (
            .in0(_gnd_net_),
            .in1(N__15049),
            .in2(N__15035),
            .in3(N__17954),
            .lcout(\eeprom.n3212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2040_3_lut_LC_18_27_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2040_3_lut_LC_18_27_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2040_3_lut_LC_18_27_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2040_3_lut_LC_18_27_2  (
            .in0(_gnd_net_),
            .in1(N__14335),
            .in2(N__13100),
            .in3(N__18119),
            .lcout(\eeprom.n3116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2037_3_lut_LC_18_27_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2037_3_lut_LC_18_27_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2037_3_lut_LC_18_27_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2037_3_lut_LC_18_27_4  (
            .in0(_gnd_net_),
            .in1(N__13181),
            .in2(N__14452),
            .in3(N__18120),
            .lcout(\eeprom.n3113 ),
            .ltout(\eeprom.n3113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_13_LC_18_27_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_13_LC_18_27_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_13_LC_18_27_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_13_LC_18_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13073),
            .in3(N__17529),
            .lcout(),
            .ltout(\eeprom.n5305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_14_LC_18_27_6 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_14_LC_18_27_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_14_LC_18_27_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_14_LC_18_27_6  (
            .in0(N__14763),
            .in1(N__17616),
            .in2(N__13070),
            .in3(N__17433),
            .lcout(\eeprom.n5309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2026_3_lut_LC_18_27_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2026_3_lut_LC_18_27_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2026_3_lut_LC_18_27_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2026_3_lut_LC_18_27_7  (
            .in0(_gnd_net_),
            .in1(N__13292),
            .in2(N__18142),
            .in3(N__14827),
            .lcout(\eeprom.n3102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2033_3_lut_LC_18_28_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2033_3_lut_LC_18_28_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2033_3_lut_LC_18_28_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2033_3_lut_LC_18_28_0  (
            .in0(_gnd_net_),
            .in1(N__14581),
            .in2(N__13154),
            .in3(N__18101),
            .lcout(\eeprom.n3109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2035_3_lut_LC_18_28_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2035_3_lut_LC_18_28_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2035_3_lut_LC_18_28_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2035_3_lut_LC_18_28_1  (
            .in0(_gnd_net_),
            .in1(N__14843),
            .in2(N__18133),
            .in3(N__13166),
            .lcout(\eeprom.n3111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2041_3_lut_LC_18_28_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2041_3_lut_LC_18_28_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2041_3_lut_LC_18_28_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2041_3_lut_LC_18_28_2  (
            .in0(_gnd_net_),
            .in1(N__13109),
            .in2(N__14492),
            .in3(N__18100),
            .lcout(\eeprom.n3117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2031_3_lut_LC_18_28_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2031_3_lut_LC_18_28_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2031_3_lut_LC_18_28_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2031_3_lut_LC_18_28_3  (
            .in0(_gnd_net_),
            .in1(N__13127),
            .in2(N__18134),
            .in3(N__14644),
            .lcout(\eeprom.n3107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i8_4_lut_adj_79_LC_18_28_4 .C_ON=1'b0;
    defparam \eeprom.i8_4_lut_adj_79_LC_18_28_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i8_4_lut_adj_79_LC_18_28_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i8_4_lut_adj_79_LC_18_28_4  (
            .in0(N__14716),
            .in1(N__14817),
            .in2(N__14620),
            .in3(N__13246),
            .lcout(\eeprom.n21_adj_336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_88_LC_18_28_6 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_88_LC_18_28_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_88_LC_18_28_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_88_LC_18_28_6  (
            .in0(N__14842),
            .in1(N__14580),
            .in2(N__14543),
            .in3(N__14654),
            .lcout(\eeprom.n3034 ),
            .ltout(\eeprom.n3034_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2039_3_lut_LC_18_28_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2039_3_lut_LC_18_28_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2039_3_lut_LC_18_28_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2039_3_lut_LC_18_28_7  (
            .in0(_gnd_net_),
            .in1(N__13193),
            .in2(N__13115),
            .in3(N__14512),
            .lcout(\eeprom.n3115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_2_lut_LC_18_29_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_2_lut_LC_18_29_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_2_lut_LC_18_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_2_lut_LC_18_29_0  (
            .in0(_gnd_net_),
            .in1(N__24196),
            .in2(_gnd_net_),
            .in3(N__13112),
            .lcout(\eeprom.n3086 ),
            .ltout(),
            .carryin(bfn_18_29_0_),
            .carryout(\eeprom.n4105 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_3_lut_LC_18_29_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_3_lut_LC_18_29_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_3_lut_LC_18_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_3_lut_LC_18_29_1  (
            .in0(_gnd_net_),
            .in1(N__14491),
            .in2(N__28560),
            .in3(N__13103),
            .lcout(\eeprom.n3085 ),
            .ltout(),
            .carryin(\eeprom.n4105 ),
            .carryout(\eeprom.n4106 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_4_lut_LC_18_29_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_4_lut_LC_18_29_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_4_lut_LC_18_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_4_lut_LC_18_29_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14342),
            .in3(N__13088),
            .lcout(\eeprom.n3084 ),
            .ltout(),
            .carryin(\eeprom.n4106 ),
            .carryout(\eeprom.n4107 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_5_lut_LC_18_29_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_5_lut_LC_18_29_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_5_lut_LC_18_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_5_lut_LC_18_29_3  (
            .in0(_gnd_net_),
            .in1(N__14513),
            .in2(_gnd_net_),
            .in3(N__13187),
            .lcout(\eeprom.n3083 ),
            .ltout(),
            .carryin(\eeprom.n4107 ),
            .carryout(\eeprom.n4108 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_6_lut_LC_18_29_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_6_lut_LC_18_29_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_6_lut_LC_18_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_6_lut_LC_18_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18281),
            .in3(N__13184),
            .lcout(\eeprom.n3082 ),
            .ltout(),
            .carryin(\eeprom.n4108 ),
            .carryout(\eeprom.n4109 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_7_lut_LC_18_29_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_7_lut_LC_18_29_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_7_lut_LC_18_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_7_lut_LC_18_29_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14456),
            .in3(N__13172),
            .lcout(\eeprom.n3081 ),
            .ltout(),
            .carryin(\eeprom.n4109 ),
            .carryout(\eeprom.n4110 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_8_lut_LC_18_29_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_8_lut_LC_18_29_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_8_lut_LC_18_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_8_lut_LC_18_29_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18260),
            .in3(N__13169),
            .lcout(\eeprom.n3080 ),
            .ltout(),
            .carryin(\eeprom.n4110 ),
            .carryout(\eeprom.n4111 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_9_lut_LC_18_29_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_9_lut_LC_18_29_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_9_lut_LC_18_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_9_lut_LC_18_29_7  (
            .in0(_gnd_net_),
            .in1(N__14841),
            .in2(N__28561),
            .in3(N__13160),
            .lcout(\eeprom.n3079 ),
            .ltout(),
            .carryin(\eeprom.n4111 ),
            .carryout(\eeprom.n4112 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_10_lut_LC_18_30_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_10_lut_LC_18_30_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_10_lut_LC_18_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_10_lut_LC_18_30_0  (
            .in0(_gnd_net_),
            .in1(N__28896),
            .in2(N__18017),
            .in3(N__13157),
            .lcout(\eeprom.n3078 ),
            .ltout(),
            .carryin(bfn_18_30_0_),
            .carryout(\eeprom.n4113 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_11_lut_LC_18_30_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_11_lut_LC_18_30_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_11_lut_LC_18_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_11_lut_LC_18_30_1  (
            .in0(_gnd_net_),
            .in1(N__28904),
            .in2(N__14582),
            .in3(N__13142),
            .lcout(\eeprom.n3077 ),
            .ltout(),
            .carryin(\eeprom.n4113 ),
            .carryout(\eeprom.n4114 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_12_lut_LC_18_30_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_12_lut_LC_18_30_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_12_lut_LC_18_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_12_lut_LC_18_30_2  (
            .in0(_gnd_net_),
            .in1(N__14315),
            .in2(N__28934),
            .in3(N__13130),
            .lcout(\eeprom.n3076 ),
            .ltout(),
            .carryin(\eeprom.n4114 ),
            .carryout(\eeprom.n4115 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_13_lut_LC_18_30_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_13_lut_LC_18_30_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_13_lut_LC_18_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_13_lut_LC_18_30_3  (
            .in0(_gnd_net_),
            .in1(N__28908),
            .in2(N__14648),
            .in3(N__13118),
            .lcout(\eeprom.n3075 ),
            .ltout(),
            .carryin(\eeprom.n4115 ),
            .carryout(\eeprom.n4116 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_14_lut_LC_18_30_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_14_lut_LC_18_30_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_14_lut_LC_18_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_14_lut_LC_18_30_4  (
            .in0(_gnd_net_),
            .in1(N__28897),
            .in2(N__14723),
            .in3(N__13304),
            .lcout(\eeprom.n3074 ),
            .ltout(),
            .carryin(\eeprom.n4116 ),
            .carryout(\eeprom.n4117 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_15_lut_LC_18_30_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_15_lut_LC_18_30_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_15_lut_LC_18_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_15_lut_LC_18_30_5  (
            .in0(_gnd_net_),
            .in1(N__14689),
            .in2(N__28932),
            .in3(N__13301),
            .lcout(\eeprom.n3073 ),
            .ltout(),
            .carryin(\eeprom.n4117 ),
            .carryout(\eeprom.n4118 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_16_lut_LC_18_30_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_16_lut_LC_18_30_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_16_lut_LC_18_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_16_lut_LC_18_30_6  (
            .in0(_gnd_net_),
            .in1(N__14621),
            .in2(N__28935),
            .in3(N__13298),
            .lcout(\eeprom.n3072 ),
            .ltout(),
            .carryin(\eeprom.n4118 ),
            .carryout(\eeprom.n4119 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_17_lut_LC_18_30_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_17_lut_LC_18_30_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_17_lut_LC_18_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_17_lut_LC_18_30_7  (
            .in0(_gnd_net_),
            .in1(N__13245),
            .in2(N__28933),
            .in3(N__13295),
            .lcout(\eeprom.n3071 ),
            .ltout(),
            .carryin(\eeprom.n4119 ),
            .carryout(\eeprom.n4120 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_18_lut_LC_18_31_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_18_lut_LC_18_31_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_18_lut_LC_18_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_18_lut_LC_18_31_0  (
            .in0(_gnd_net_),
            .in1(N__14828),
            .in2(N__28936),
            .in3(N__13280),
            .lcout(\eeprom.n3070 ),
            .ltout(),
            .carryin(bfn_18_31_0_),
            .carryout(\eeprom.n4121 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_19_lut_LC_18_31_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2022_19_lut_LC_18_31_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_19_lut_LC_18_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2022_19_lut_LC_18_31_1  (
            .in0(_gnd_net_),
            .in1(N__14564),
            .in2(N__28937),
            .in3(N__13262),
            .lcout(\eeprom.n3069 ),
            .ltout(),
            .carryin(\eeprom.n4121 ),
            .carryout(\eeprom.n4122 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2022_20_lut_LC_18_31_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2022_20_lut_LC_18_31_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2022_20_lut_LC_18_31_2 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2022_20_lut_LC_18_31_2  (
            .in0(N__28915),
            .in1(N__18673),
            .in2(N__18145),
            .in3(N__13259),
            .lcout(\eeprom.n3100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2027_3_lut_LC_18_31_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2027_3_lut_LC_18_31_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2027_3_lut_LC_18_31_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2027_3_lut_LC_18_31_5  (
            .in0(_gnd_net_),
            .in1(N__13256),
            .in2(N__13250),
            .in3(N__18138),
            .lcout(\eeprom.n3103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2444_3_lut_LC_19_17_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2444_3_lut_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2444_3_lut_LC_19_17_1 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \eeprom.rem_4_i2444_3_lut_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(N__13226),
            .in2(N__13202),
            .in3(N__13429),
            .lcout(\eeprom.n3712 ),
            .ltout(\eeprom.n3712_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4735_1_lut_LC_19_17_2 .C_ON=1'b0;
    defparam \eeprom.i4735_1_lut_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4735_1_lut_LC_19_17_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4735_1_lut_LC_19_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13391),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2449_3_lut_LC_19_17_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2449_3_lut_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2449_3_lut_LC_19_17_3 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \eeprom.rem_4_i2449_3_lut_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__13388),
            .in2(N__13382),
            .in3(N__13428),
            .lcout(\eeprom.n3717 ),
            .ltout(\eeprom.n3717_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4720_1_lut_LC_19_17_4 .C_ON=1'b0;
    defparam \eeprom.i4720_1_lut_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4720_1_lut_LC_19_17_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4720_1_lut_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13367),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2450_rep_4_3_lut_LC_19_17_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2450_rep_4_3_lut_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2450_rep_4_3_lut_LC_19_17_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \eeprom.rem_4_i2450_rep_4_3_lut_LC_19_17_5  (
            .in0(N__13364),
            .in1(N__21578),
            .in2(_gnd_net_),
            .in3(N__13426),
            .lcout(\eeprom.n5362 ),
            .ltout(\eeprom.n5362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4717_1_lut_LC_19_17_6 .C_ON=1'b0;
    defparam \eeprom.i4717_1_lut_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4717_1_lut_LC_19_17_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4717_1_lut_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13358),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2448_3_lut_LC_19_17_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2448_3_lut_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2448_3_lut_LC_19_17_7 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \eeprom.rem_4_i2448_3_lut_LC_19_17_7  (
            .in0(_gnd_net_),
            .in1(N__13567),
            .in2(N__13355),
            .in3(N__13427),
            .lcout(\eeprom.n3716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2447_3_lut_LC_19_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2447_3_lut_LC_19_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2447_3_lut_LC_19_18_0 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \eeprom.rem_4_i2447_3_lut_LC_19_18_0  (
            .in0(_gnd_net_),
            .in1(N__13346),
            .in2(N__13339),
            .in3(N__13430),
            .lcout(\eeprom.n3715 ),
            .ltout(\eeprom.n3715_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4726_1_lut_LC_19_18_1 .C_ON=1'b0;
    defparam \eeprom.i4726_1_lut_LC_19_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4726_1_lut_LC_19_18_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4726_1_lut_LC_19_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13313),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_101_LC_19_18_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_101_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_101_LC_19_18_2 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \eeprom.i1_4_lut_adj_101_LC_19_18_2  (
            .in0(N__16329),
            .in1(N__15935),
            .in2(N__19088),
            .in3(N__13310),
            .lcout(),
            .ltout(\eeprom.n5019_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_103_LC_19_18_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_103_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_103_LC_19_18_3 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \eeprom.i1_4_lut_adj_103_LC_19_18_3  (
            .in0(N__16424),
            .in1(N__16403),
            .in2(N__13484),
            .in3(N__16330),
            .lcout(),
            .ltout(\eeprom.n28_adj_342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_104_LC_19_18_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_104_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_104_LC_19_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_104_LC_19_18_4  (
            .in0(N__13544),
            .in1(N__16211),
            .in2(N__13481),
            .in3(N__13595),
            .lcout(\eeprom.n3628 ),
            .ltout(\eeprom.n3628_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2446_3_lut_LC_19_18_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2446_3_lut_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2446_3_lut_LC_19_18_5 .LUT_INIT=16'b0000010111110101;
    LogicCell40 \eeprom.rem_4_i2446_3_lut_LC_19_18_5  (
            .in0(N__13477),
            .in1(_gnd_net_),
            .in2(N__13463),
            .in3(N__13460),
            .lcout(\eeprom.n3714 ),
            .ltout(\eeprom.n3714_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4729_1_lut_LC_19_18_6 .C_ON=1'b0;
    defparam \eeprom.i4729_1_lut_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4729_1_lut_LC_19_18_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4729_1_lut_LC_19_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13454),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4741_2_lut_LC_19_18_7 .C_ON=1'b0;
    defparam \eeprom.i4741_2_lut_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4741_2_lut_LC_19_18_7 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \eeprom.i4741_2_lut_LC_19_18_7  (
            .in0(N__13450),
            .in1(_gnd_net_),
            .in2(N__13436),
            .in3(_gnd_net_),
            .lcout(\eeprom.n3711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_93_LC_19_19_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_93_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_93_LC_19_19_0 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \eeprom.i1_4_lut_adj_93_LC_19_19_0  (
            .in0(N__15977),
            .in1(N__16003),
            .in2(N__16321),
            .in3(N__13529),
            .lcout(),
            .ltout(\eeprom.n5025_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_94_LC_19_19_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_94_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_94_LC_19_19_1 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \eeprom.i1_4_lut_adj_94_LC_19_19_1  (
            .in0(N__15961),
            .in1(N__15947),
            .in2(N__13400),
            .in3(N__16297),
            .lcout(),
            .ltout(\eeprom.n5027_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_95_LC_19_19_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_95_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_95_LC_19_19_2 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \eeprom.i1_4_lut_adj_95_LC_19_19_2  (
            .in0(N__16298),
            .in1(N__15893),
            .in2(N__13397),
            .in3(N__15920),
            .lcout(),
            .ltout(\eeprom.n5029_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_98_LC_19_19_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_98_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_98_LC_19_19_3 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \eeprom.i1_4_lut_adj_98_LC_19_19_3  (
            .in0(N__16466),
            .in1(N__16486),
            .in2(N__13394),
            .in3(N__16299),
            .lcout(),
            .ltout(\eeprom.n5031_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_102_LC_19_19_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_102_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_102_LC_19_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_102_LC_19_19_4  (
            .in0(N__13579),
            .in1(N__13616),
            .in2(N__13598),
            .in3(N__13625),
            .lcout(\eeprom.n5161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_24_LC_19_19_5 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_24_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_24_LC_19_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_24_LC_19_19_5  (
            .in0(N__15960),
            .in1(N__15915),
            .in2(N__16487),
            .in3(N__19084),
            .lcout(\eeprom.n29_adj_274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2376_3_lut_LC_19_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2376_3_lut_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2376_3_lut_LC_19_19_6 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \eeprom.rem_4_i2376_3_lut_LC_19_19_6  (
            .in0(N__15757),
            .in1(N__15743),
            .in2(N__16322),
            .in3(_gnd_net_),
            .lcout(\eeprom.n3612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2381_3_lut_LC_19_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2381_3_lut_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2381_3_lut_LC_19_19_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2381_3_lut_LC_19_19_7  (
            .in0(_gnd_net_),
            .in1(N__15469),
            .in2(N__15449),
            .in3(N__16290),
            .lcout(\eeprom.n3617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2360_3_lut_LC_19_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2360_3_lut_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2360_3_lut_LC_19_20_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2360_3_lut_LC_19_20_0  (
            .in0(N__16364),
            .in1(_gnd_net_),
            .in2(N__16319),
            .in3(N__16390),
            .lcout(\eeprom.n3596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2373_3_lut_LC_19_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2373_3_lut_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2373_3_lut_LC_19_20_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2373_3_lut_LC_19_20_1  (
            .in0(_gnd_net_),
            .in1(N__15655),
            .in2(N__15635),
            .in3(N__16277),
            .lcout(),
            .ltout(\eeprom.n3609_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_91_LC_19_20_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_91_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_91_LC_19_20_2 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \eeprom.i1_4_lut_adj_91_LC_19_20_2  (
            .in0(N__16278),
            .in1(N__16130),
            .in2(N__13535),
            .in3(N__16100),
            .lcout(),
            .ltout(\eeprom.n5021_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_92_LC_19_20_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_92_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_92_LC_19_20_3 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \eeprom.i1_4_lut_adj_92_LC_19_20_3  (
            .in0(N__16091),
            .in1(N__16073),
            .in2(N__13532),
            .in3(N__16279),
            .lcout(\eeprom.n5023 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2302_3_lut_LC_19_20_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2302_3_lut_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2302_3_lut_LC_19_20_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2302_3_lut_LC_19_20_5  (
            .in0(_gnd_net_),
            .in1(N__13523),
            .in2(N__19220),
            .in3(N__13511),
            .lcout(\eeprom.n3506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2314_rep_5_3_lut_LC_19_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2314_rep_5_3_lut_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2314_rep_5_3_lut_LC_19_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i2314_rep_5_3_lut_LC_19_20_6  (
            .in0(N__13673),
            .in1(N__23426),
            .in2(_gnd_net_),
            .in3(N__19196),
            .lcout(\eeprom.n3518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2296_3_lut_LC_19_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2296_3_lut_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2296_3_lut_LC_19_20_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2296_3_lut_LC_19_20_7  (
            .in0(N__14075),
            .in1(_gnd_net_),
            .in2(N__19219),
            .in3(N__13661),
            .lcout(\eeprom.n3500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2372_3_lut_LC_19_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2372_3_lut_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2372_3_lut_LC_19_21_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2372_3_lut_LC_19_21_0  (
            .in0(N__15593),
            .in1(_gnd_net_),
            .in2(N__15619),
            .in3(N__16283),
            .lcout(),
            .ltout(\eeprom.n3608_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_90_LC_19_21_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_90_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_90_LC_19_21_1 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \eeprom.i1_4_lut_adj_90_LC_19_21_1  (
            .in0(N__16284),
            .in1(N__15671),
            .in2(N__13649),
            .in3(N__15691),
            .lcout(\eeprom.n5175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2308_3_lut_LC_19_21_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2308_3_lut_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2308_3_lut_LC_19_21_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2308_3_lut_LC_19_21_2  (
            .in0(_gnd_net_),
            .in1(N__13646),
            .in2(N__19204),
            .in3(N__16510),
            .lcout(\eeprom.n3512 ),
            .ltout(\eeprom.n3512_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_96_LC_19_21_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_96_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_96_LC_19_21_3 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \eeprom.i1_4_lut_adj_96_LC_19_21_3  (
            .in0(N__16285),
            .in1(N__15713),
            .in2(N__13637),
            .in3(N__13634),
            .lcout(),
            .ltout(\eeprom.n5177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_97_LC_19_21_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_97_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_97_LC_19_21_4 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \eeprom.i1_4_lut_adj_97_LC_19_21_4  (
            .in0(N__16031),
            .in1(N__16013),
            .in2(N__13628),
            .in3(N__16289),
            .lcout(\eeprom.n31_adj_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2362_3_lut_LC_19_21_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2362_3_lut_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2362_3_lut_LC_19_21_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2362_3_lut_LC_19_21_5  (
            .in0(_gnd_net_),
            .in1(N__16433),
            .in2(N__16320),
            .in3(N__16453),
            .lcout(\eeprom.n3598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2311_3_lut_LC_19_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2311_3_lut_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2311_3_lut_LC_19_21_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2311_3_lut_LC_19_21_6  (
            .in0(_gnd_net_),
            .in1(N__13607),
            .in2(N__19203),
            .in3(N__16618),
            .lcout(\eeprom.n3515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2313_3_lut_LC_19_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2313_3_lut_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2313_3_lut_LC_19_21_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2313_3_lut_LC_19_21_7  (
            .in0(_gnd_net_),
            .in1(N__16657),
            .in2(N__13832),
            .in3(N__19161),
            .lcout(\eeprom.n3517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_LC_19_22_1 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_LC_19_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_LC_19_22_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_LC_19_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13820),
            .in3(N__13799),
            .lcout(),
            .ltout(\eeprom.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_LC_19_22_2 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_LC_19_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_LC_19_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_LC_19_22_2  (
            .in0(N__13779),
            .in1(N__13755),
            .in2(N__13736),
            .in3(N__17022),
            .lcout(),
            .ltout(\eeprom.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i16_4_lut_LC_19_22_3 .C_ON=1'b0;
    defparam \eeprom.i16_4_lut_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i16_4_lut_LC_19_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i16_4_lut_LC_19_22_3  (
            .in0(N__13733),
            .in1(N__14012),
            .in2(N__13727),
            .in3(N__16682),
            .lcout(\eeprom.n3430 ),
            .ltout(\eeprom.n3430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2295_3_lut_LC_19_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2295_3_lut_LC_19_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2295_3_lut_LC_19_22_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2295_3_lut_LC_19_22_4  (
            .in0(_gnd_net_),
            .in1(N__14056),
            .in2(N__13724),
            .in3(N__13721),
            .lcout(\eeprom.n3499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2294_3_lut_LC_19_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2294_3_lut_LC_19_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2294_3_lut_LC_19_22_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2294_3_lut_LC_19_22_5  (
            .in0(_gnd_net_),
            .in1(N__14035),
            .in2(N__19222),
            .in3(N__13709),
            .lcout(\eeprom.n3498 ),
            .ltout(\eeprom.n3498_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_18_LC_19_22_6 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_18_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_18_LC_19_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_18_LC_19_22_6  (
            .in0(N__16351),
            .in1(N__16380),
            .in2(N__13697),
            .in3(N__16449),
            .lcout(\eeprom.n28_adj_267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2304_3_lut_LC_19_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2304_3_lut_LC_19_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2304_3_lut_LC_19_22_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2304_3_lut_LC_19_22_7  (
            .in0(N__19214),
            .in1(_gnd_net_),
            .in2(N__17029),
            .in3(N__13682),
            .lcout(\eeprom.n3508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2233_3_lut_LC_19_23_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2233_3_lut_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2233_3_lut_LC_19_23_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2233_3_lut_LC_19_23_1  (
            .in0(_gnd_net_),
            .in1(N__14209),
            .in2(N__14105),
            .in3(N__17147),
            .lcout(\eeprom.n3405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2229_3_lut_LC_19_23_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2229_3_lut_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2229_3_lut_LC_19_23_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \eeprom.rem_4_i2229_3_lut_LC_19_23_2  (
            .in0(N__17148),
            .in1(_gnd_net_),
            .in2(N__14090),
            .in3(N__16790),
            .lcout(\eeprom.n3401 ),
            .ltout(\eeprom.n3401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_17_LC_19_23_3 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_17_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_17_LC_19_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_17_LC_19_23_3  (
            .in0(N__14052),
            .in1(N__14031),
            .in2(N__14015),
            .in3(N__14001),
            .lcout(\eeprom.n27_adj_263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2297_3_lut_LC_19_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2297_3_lut_LC_19_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2297_3_lut_LC_19_23_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i2297_3_lut_LC_19_23_4  (
            .in0(N__14002),
            .in1(_gnd_net_),
            .in2(N__13988),
            .in3(N__19190),
            .lcout(\eeprom.n3501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_111_LC_19_23_5 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_111_LC_19_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_111_LC_19_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_111_LC_19_23_5  (
            .in0(N__13968),
            .in1(N__13950),
            .in2(N__13924),
            .in3(N__13897),
            .lcout(),
            .ltout(\eeprom.n28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i15_4_lut_LC_19_23_6 .C_ON=1'b0;
    defparam \eeprom.i15_4_lut_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i15_4_lut_LC_19_23_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i15_4_lut_LC_19_23_6  (
            .in0(N__14141),
            .in1(N__16757),
            .in2(N__13871),
            .in3(N__13868),
            .lcout(\eeprom.n3331 ),
            .ltout(\eeprom.n3331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2245_3_lut_LC_19_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2245_3_lut_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2245_3_lut_LC_19_23_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2245_3_lut_LC_19_23_7  (
            .in0(_gnd_net_),
            .in1(N__13862),
            .in2(N__13850),
            .in3(N__16878),
            .lcout(\eeprom.n3417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2173_3_lut_LC_19_24_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2173_3_lut_LC_19_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2173_3_lut_LC_19_24_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2173_3_lut_LC_19_24_1  (
            .in0(_gnd_net_),
            .in1(N__17509),
            .in2(N__13847),
            .in3(N__17736),
            .lcout(\eeprom.n3313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_36_LC_19_24_2 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_36_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_36_LC_19_24_2 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \eeprom.i5_4_lut_adj_36_LC_19_24_2  (
            .in0(N__24236),
            .in1(N__14358),
            .in2(N__17456),
            .in3(N__16990),
            .lcout(),
            .ltout(\eeprom.n20_adj_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_adj_40_LC_19_24_3 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_adj_40_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_adj_40_LC_19_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_adj_40_LC_19_24_3  (
            .in0(N__14422),
            .in1(N__14287),
            .in2(N__14273),
            .in3(N__18167),
            .lcout(),
            .ltout(\eeprom.n28_adj_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i14_4_lut_LC_19_24_4 .C_ON=1'b0;
    defparam \eeprom.i14_4_lut_LC_19_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i14_4_lut_LC_19_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i14_4_lut_LC_19_24_4  (
            .in0(N__14270),
            .in1(N__14260),
            .in2(N__14240),
            .in3(N__14237),
            .lcout(\eeprom.n3232 ),
            .ltout(\eeprom.n3232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2166_3_lut_LC_19_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2166_3_lut_LC_19_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2166_3_lut_LC_19_24_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2166_3_lut_LC_19_24_5  (
            .in0(N__14359),
            .in1(_gnd_net_),
            .in2(N__14231),
            .in3(N__14228),
            .lcout(\eeprom.n3306 ),
            .ltout(\eeprom.n3306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_113_LC_19_24_6 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_113_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_113_LC_19_24_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_113_LC_19_24_6  (
            .in0(N__14187),
            .in1(N__17170),
            .in2(N__14171),
            .in3(N__14157),
            .lcout(\eeprom.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4_4_lut_LC_19_25_0 .C_ON=1'b0;
    defparam \eeprom.i4_4_lut_LC_19_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4_4_lut_LC_19_25_0 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \eeprom.i4_4_lut_LC_19_25_0  (
            .in0(N__22412),
            .in1(N__14874),
            .in2(N__17359),
            .in3(N__14135),
            .lcout(),
            .ltout(\eeprom.n18_adj_260_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i12_4_lut_adj_15_LC_19_25_1 .C_ON=1'b0;
    defparam \eeprom.i12_4_lut_adj_15_LC_19_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i12_4_lut_adj_15_LC_19_25_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i12_4_lut_adj_15_LC_19_25_1  (
            .in0(N__15312),
            .in1(N__15270),
            .in2(N__14126),
            .in3(N__14123),
            .lcout(),
            .ltout(\eeprom.n26_adj_262_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i13_4_lut_adj_16_LC_19_25_2 .C_ON=1'b0;
    defparam \eeprom.i13_4_lut_adj_16_LC_19_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i13_4_lut_adj_16_LC_19_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i13_4_lut_adj_16_LC_19_25_2  (
            .in0(N__14117),
            .in1(N__17983),
            .in2(N__14111),
            .in3(N__18033),
            .lcout(\eeprom.n3133 ),
            .ltout(\eeprom.n3133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2103_3_lut_LC_19_25_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2103_3_lut_LC_19_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2103_3_lut_LC_19_25_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i2103_3_lut_LC_19_25_3  (
            .in0(N__18034),
            .in1(_gnd_net_),
            .in2(N__14108),
            .in3(N__15017),
            .lcout(\eeprom.n3211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2097_3_lut_LC_19_25_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2097_3_lut_LC_19_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2097_3_lut_LC_19_25_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2097_3_lut_LC_19_25_4  (
            .in0(_gnd_net_),
            .in1(N__14855),
            .in2(N__17956),
            .in3(N__14875),
            .lcout(\eeprom.n3205 ),
            .ltout(\eeprom.n3205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2164_3_lut_LC_19_25_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2164_3_lut_LC_19_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2164_3_lut_LC_19_25_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2164_3_lut_LC_19_25_5  (
            .in0(_gnd_net_),
            .in1(N__14408),
            .in2(N__14396),
            .in3(N__17762),
            .lcout(\eeprom.n3304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2163_3_lut_LC_19_25_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2163_3_lut_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2163_3_lut_LC_19_25_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2163_3_lut_LC_19_25_6  (
            .in0(_gnd_net_),
            .in1(N__14392),
            .in2(N__17778),
            .in3(N__14378),
            .lcout(\eeprom.n3303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2099_3_lut_LC_19_25_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2099_3_lut_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2099_3_lut_LC_19_25_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2099_3_lut_LC_19_25_7  (
            .in0(_gnd_net_),
            .in1(N__14930),
            .in2(N__14950),
            .in3(N__17941),
            .lcout(\eeprom.n3207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1973_3_lut_LC_19_26_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1973_3_lut_LC_19_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1973_3_lut_LC_19_26_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1973_3_lut_LC_19_26_0  (
            .in0(_gnd_net_),
            .in1(N__18380),
            .in2(N__19478),
            .in3(N__18740),
            .lcout(\eeprom.n3017 ),
            .ltout(\eeprom.n3017_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_77_LC_19_26_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_77_LC_19_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_77_LC_19_26_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_77_LC_19_26_1  (
            .in0(N__14508),
            .in1(N__14442),
            .in2(N__14321),
            .in3(N__18236),
            .lcout(),
            .ltout(\eeprom.n5147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_78_LC_19_26_2 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_78_LC_19_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_78_LC_19_26_2 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \eeprom.i5_4_lut_adj_78_LC_19_26_2  (
            .in0(N__24189),
            .in1(N__14487),
            .in2(N__14318),
            .in3(N__14304),
            .lcout(\eeprom.n18_adj_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2108_3_lut_LC_19_26_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2108_3_lut_LC_19_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2108_3_lut_LC_19_26_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2108_3_lut_LC_19_26_3  (
            .in0(_gnd_net_),
            .in1(N__14744),
            .in2(N__14774),
            .in3(N__17922),
            .lcout(\eeprom.n3216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1965_3_lut_LC_19_26_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1965_3_lut_LC_19_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1965_3_lut_LC_19_26_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1965_3_lut_LC_19_26_4  (
            .in0(_gnd_net_),
            .in1(N__18476),
            .in2(N__18494),
            .in3(N__18741),
            .lcout(\eeprom.n3009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1958_3_lut_LC_19_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1958_3_lut_LC_19_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1958_3_lut_LC_19_26_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1958_3_lut_LC_19_26_5  (
            .in0(_gnd_net_),
            .in1(N__18800),
            .in2(N__18774),
            .in3(N__19718),
            .lcout(\eeprom.n3002 ),
            .ltout(\eeprom.n3002_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_3_lut_LC_19_26_6 .C_ON=1'b0;
    defparam \eeprom.i7_3_lut_LC_19_26_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_3_lut_LC_19_26_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \eeprom.i7_3_lut_LC_19_26_6  (
            .in0(_gnd_net_),
            .in1(N__18013),
            .in2(N__14546),
            .in3(N__18674),
            .lcout(\eeprom.n20_adj_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2034_3_lut_LC_19_27_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2034_3_lut_LC_19_27_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2034_3_lut_LC_19_27_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2034_3_lut_LC_19_27_0  (
            .in0(_gnd_net_),
            .in1(N__18009),
            .in2(N__14528),
            .in3(N__18128),
            .lcout(\eeprom.n3110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1972_3_lut_LC_19_27_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1972_3_lut_LC_19_27_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1972_3_lut_LC_19_27_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1972_3_lut_LC_19_27_1  (
            .in0(N__18364),
            .in1(_gnd_net_),
            .in2(N__18350),
            .in3(N__18745),
            .lcout(\eeprom.n3016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1974_3_lut_LC_19_27_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1974_3_lut_LC_19_27_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1974_3_lut_LC_19_27_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i1974_3_lut_LC_19_27_2  (
            .in0(N__18395),
            .in1(N__22466),
            .in2(N__18775),
            .in3(_gnd_net_),
            .lcout(\eeprom.n3018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1902_3_lut_LC_19_27_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1902_3_lut_LC_19_27_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1902_3_lut_LC_19_27_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1902_3_lut_LC_19_27_3  (
            .in0(_gnd_net_),
            .in1(N__20858),
            .in2(N__19379),
            .in3(N__19670),
            .lcout(\eeprom.n2914 ),
            .ltout(\eeprom.n2914_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_34_LC_19_27_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_34_LC_19_27_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_34_LC_19_27_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_34_LC_19_27_4  (
            .in0(N__18327),
            .in1(N__18363),
            .in2(N__14468),
            .in3(N__18401),
            .lcout(\eeprom.n5301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2029_3_lut_LC_19_27_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2029_3_lut_LC_19_27_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2029_3_lut_LC_19_27_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2029_3_lut_LC_19_27_6  (
            .in0(N__14465),
            .in1(_gnd_net_),
            .in2(N__14690),
            .in3(N__18129),
            .lcout(\eeprom.n3105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1970_3_lut_LC_19_27_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1970_3_lut_LC_19_27_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1970_3_lut_LC_19_27_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1970_3_lut_LC_19_27_7  (
            .in0(_gnd_net_),
            .in1(N__18593),
            .in2(N__18617),
            .in3(N__18746),
            .lcout(\eeprom.n3014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1963_3_lut_LC_19_28_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1963_3_lut_LC_19_28_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1963_3_lut_LC_19_28_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1963_3_lut_LC_19_28_0  (
            .in0(_gnd_net_),
            .in1(N__18884),
            .in2(N__18776),
            .in3(N__18427),
            .lcout(\eeprom.n3007 ),
            .ltout(\eeprom.n3007_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2030_3_lut_LC_19_28_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2030_3_lut_LC_19_28_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2030_3_lut_LC_19_28_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2030_3_lut_LC_19_28_1  (
            .in0(_gnd_net_),
            .in1(N__14705),
            .in2(N__14693),
            .in3(N__18109),
            .lcout(\eeprom.n3106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1962_3_lut_LC_19_28_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1962_3_lut_LC_19_28_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1962_3_lut_LC_19_28_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1962_3_lut_LC_19_28_2  (
            .in0(_gnd_net_),
            .in1(N__18872),
            .in2(N__18778),
            .in3(N__19589),
            .lcout(\eeprom.n3006 ),
            .ltout(\eeprom.n3006_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_85_LC_19_28_3 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_85_LC_19_28_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_85_LC_19_28_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_85_LC_19_28_3  (
            .in0(N__14672),
            .in1(N__14643),
            .in2(N__14666),
            .in3(N__14663),
            .lcout(\eeprom.n24_adj_340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1964_3_lut_LC_19_28_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1964_3_lut_LC_19_28_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1964_3_lut_LC_19_28_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1964_3_lut_LC_19_28_4  (
            .in0(_gnd_net_),
            .in1(N__18440),
            .in2(N__18777),
            .in3(N__18461),
            .lcout(\eeprom.n3008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1961_3_lut_LC_19_28_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1961_3_lut_LC_19_28_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1961_3_lut_LC_19_28_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \eeprom.rem_4_i1961_3_lut_LC_19_28_5  (
            .in0(_gnd_net_),
            .in1(N__18753),
            .in2(N__18860),
            .in3(N__18836),
            .lcout(\eeprom.n3005 ),
            .ltout(\eeprom.n3005_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2028_3_lut_LC_19_28_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2028_3_lut_LC_19_28_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2028_3_lut_LC_19_28_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2028_3_lut_LC_19_28_6  (
            .in0(N__18110),
            .in1(_gnd_net_),
            .in2(N__14603),
            .in3(N__14600),
            .lcout(\eeprom.n3104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2038_3_lut_LC_19_28_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2038_3_lut_LC_19_28_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2038_3_lut_LC_19_28_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i2038_3_lut_LC_19_28_7  (
            .in0(N__18277),
            .in1(N__14588),
            .in2(_gnd_net_),
            .in3(N__18108),
            .lcout(\eeprom.n3114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1966_3_lut_LC_19_29_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1966_3_lut_LC_19_29_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1966_3_lut_LC_19_29_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1966_3_lut_LC_19_29_0  (
            .in0(_gnd_net_),
            .in1(N__18503),
            .in2(N__18784),
            .in3(N__19448),
            .lcout(\eeprom.n3010 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1968_3_lut_LC_19_29_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1968_3_lut_LC_19_29_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1968_3_lut_LC_19_29_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1968_3_lut_LC_19_29_1  (
            .in0(_gnd_net_),
            .in1(N__18545),
            .in2(N__18533),
            .in3(N__18770),
            .lcout(\eeprom.n3012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1959_3_lut_LC_19_29_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1959_3_lut_LC_19_29_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1959_3_lut_LC_19_29_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1959_3_lut_LC_19_29_4  (
            .in0(_gnd_net_),
            .in1(N__18809),
            .in2(N__18783),
            .in3(N__19775),
            .lcout(\eeprom.n3003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2042_3_lut_LC_19_29_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2042_3_lut_LC_19_29_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2042_3_lut_LC_19_29_5 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i2042_3_lut_LC_19_29_5  (
            .in0(N__14801),
            .in1(N__24197),
            .in2(N__18143),
            .in3(_gnd_net_),
            .lcout(\eeprom.n3118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_2_lut_LC_19_30_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_2_lut_LC_19_30_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_2_lut_LC_19_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_2_lut_LC_19_30_0  (
            .in0(_gnd_net_),
            .in1(N__22411),
            .in2(_gnd_net_),
            .in3(N__14780),
            .lcout(\eeprom.n3186 ),
            .ltout(),
            .carryin(bfn_19_30_0_),
            .carryout(\eeprom.n4123 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_3_lut_LC_19_30_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_3_lut_LC_19_30_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_3_lut_LC_19_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_3_lut_LC_19_30_1  (
            .in0(_gnd_net_),
            .in1(N__28562),
            .in2(N__17352),
            .in3(N__14777),
            .lcout(\eeprom.n3185 ),
            .ltout(),
            .carryin(\eeprom.n4123 ),
            .carryout(\eeprom.n4124 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_4_lut_LC_19_30_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_4_lut_LC_19_30_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_4_lut_LC_19_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_4_lut_LC_19_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14773),
            .in3(N__14735),
            .lcout(\eeprom.n3184 ),
            .ltout(),
            .carryin(\eeprom.n4124 ),
            .carryout(\eeprom.n4125 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_5_lut_LC_19_30_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_5_lut_LC_19_30_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_5_lut_LC_19_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_5_lut_LC_19_30_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17446),
            .in3(N__14732),
            .lcout(\eeprom.n3183 ),
            .ltout(),
            .carryin(\eeprom.n4125 ),
            .carryout(\eeprom.n4126 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_6_lut_LC_19_30_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_6_lut_LC_19_30_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_6_lut_LC_19_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_6_lut_LC_19_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17542),
            .in3(N__14729),
            .lcout(\eeprom.n3182 ),
            .ltout(),
            .carryin(\eeprom.n4126 ),
            .carryout(\eeprom.n4127 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_7_lut_LC_19_30_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_7_lut_LC_19_30_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_7_lut_LC_19_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_7_lut_LC_19_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17629),
            .in3(N__14726),
            .lcout(\eeprom.n3181 ),
            .ltout(),
            .carryin(\eeprom.n4127 ),
            .carryout(\eeprom.n4128 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_8_lut_LC_19_30_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_8_lut_LC_19_30_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_8_lut_LC_19_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_8_lut_LC_19_30_6  (
            .in0(_gnd_net_),
            .in1(N__15050),
            .in2(_gnd_net_),
            .in3(N__15020),
            .lcout(\eeprom.n3180 ),
            .ltout(),
            .carryin(\eeprom.n4128 ),
            .carryout(\eeprom.n4129 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_9_lut_LC_19_30_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_9_lut_LC_19_30_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_9_lut_LC_19_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_9_lut_LC_19_30_7  (
            .in0(_gnd_net_),
            .in1(N__28563),
            .in2(N__18041),
            .in3(N__15005),
            .lcout(\eeprom.n3179 ),
            .ltout(),
            .carryin(\eeprom.n4129 ),
            .carryout(\eeprom.n4130 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_10_lut_LC_19_31_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_10_lut_LC_19_31_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_10_lut_LC_19_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_10_lut_LC_19_31_0  (
            .in0(_gnd_net_),
            .in1(N__15002),
            .in2(N__28710),
            .in3(N__14963),
            .lcout(\eeprom.n3178 ),
            .ltout(),
            .carryin(bfn_19_31_0_),
            .carryout(\eeprom.n4131 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_11_lut_LC_19_31_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_11_lut_LC_19_31_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_11_lut_LC_19_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_11_lut_LC_19_31_1  (
            .in0(_gnd_net_),
            .in1(N__17984),
            .in2(N__28713),
            .in3(N__14960),
            .lcout(\eeprom.n3177 ),
            .ltout(),
            .carryin(\eeprom.n4131 ),
            .carryout(\eeprom.n4132 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_12_lut_LC_19_31_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_12_lut_LC_19_31_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_12_lut_LC_19_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_12_lut_LC_19_31_2  (
            .in0(_gnd_net_),
            .in1(N__17299),
            .in2(N__28711),
            .in3(N__14957),
            .lcout(\eeprom.n3176 ),
            .ltout(),
            .carryin(\eeprom.n4132 ),
            .carryout(\eeprom.n4133 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_13_lut_LC_19_31_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_13_lut_LC_19_31_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_13_lut_LC_19_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_13_lut_LC_19_31_3  (
            .in0(_gnd_net_),
            .in1(N__28576),
            .in2(N__14954),
            .in3(N__14918),
            .lcout(\eeprom.n3175 ),
            .ltout(),
            .carryin(\eeprom.n4133 ),
            .carryout(\eeprom.n4134 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_14_lut_LC_19_31_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_14_lut_LC_19_31_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_14_lut_LC_19_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_14_lut_LC_19_31_4  (
            .in0(_gnd_net_),
            .in1(N__14914),
            .in2(N__28712),
            .in3(N__14879),
            .lcout(\eeprom.n3174 ),
            .ltout(),
            .carryin(\eeprom.n4134 ),
            .carryout(\eeprom.n4135 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_15_lut_LC_19_31_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_15_lut_LC_19_31_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_15_lut_LC_19_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_15_lut_LC_19_31_5  (
            .in0(_gnd_net_),
            .in1(N__14876),
            .in2(N__28714),
            .in3(N__14846),
            .lcout(\eeprom.n3173 ),
            .ltout(),
            .carryin(\eeprom.n4135 ),
            .carryout(\eeprom.n4136 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_16_lut_LC_19_31_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_16_lut_LC_19_31_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_16_lut_LC_19_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_16_lut_LC_19_31_6  (
            .in0(_gnd_net_),
            .in1(N__28586),
            .in2(N__15319),
            .in3(N__15278),
            .lcout(\eeprom.n3172 ),
            .ltout(),
            .carryin(\eeprom.n4136 ),
            .carryout(\eeprom.n4137 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_17_lut_LC_19_31_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_17_lut_LC_19_31_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_17_lut_LC_19_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_17_lut_LC_19_31_7  (
            .in0(_gnd_net_),
            .in1(N__15271),
            .in2(N__28715),
            .in3(N__15233),
            .lcout(\eeprom.n3171 ),
            .ltout(),
            .carryin(\eeprom.n4137 ),
            .carryout(\eeprom.n4138 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_18_lut_LC_19_32_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_18_lut_LC_19_32_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_18_lut_LC_19_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_18_lut_LC_19_32_0  (
            .in0(_gnd_net_),
            .in1(N__15225),
            .in2(N__28708),
            .in3(N__15194),
            .lcout(\eeprom.n3170 ),
            .ltout(),
            .carryin(bfn_19_32_0_),
            .carryout(\eeprom.n4139 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_19_lut_LC_19_32_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_19_lut_LC_19_32_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_19_lut_LC_19_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_19_lut_LC_19_32_1  (
            .in0(_gnd_net_),
            .in1(N__15191),
            .in2(N__28716),
            .in3(N__15155),
            .lcout(\eeprom.n3169 ),
            .ltout(),
            .carryin(\eeprom.n4139 ),
            .carryout(\eeprom.n4140 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_20_lut_LC_19_32_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2089_20_lut_LC_19_32_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_20_lut_LC_19_32_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2089_20_lut_LC_19_32_2  (
            .in0(_gnd_net_),
            .in1(N__15152),
            .in2(N__28709),
            .in3(N__15107),
            .lcout(\eeprom.n3168 ),
            .ltout(),
            .carryin(\eeprom.n4140 ),
            .carryout(\eeprom.n4141 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2089_21_lut_LC_19_32_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2089_21_lut_LC_19_32_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2089_21_lut_LC_19_32_3 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2089_21_lut_LC_19_32_3  (
            .in0(N__28593),
            .in1(N__15100),
            .in2(N__17957),
            .in3(N__15086),
            .lcout(\eeprom.n3199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_2_lut_LC_20_17_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_2_lut_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_2_lut_LC_20_17_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_2_lut_LC_20_17_0  (
            .in0(N__25496),
            .in1(N__26708),
            .in2(N__25379),
            .in3(N__15056),
            .lcout(\eeprom.enable_N_60_0 ),
            .ltout(),
            .carryin(bfn_20_17_0_),
            .carryout(\eeprom.n4228 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_3_lut_LC_20_17_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_3_lut_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_3_lut_LC_20_17_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_3_lut_LC_20_17_1  (
            .in0(N__25667),
            .in1(N__23066),
            .in2(N__26737),
            .in3(N__15053),
            .lcout(\eeprom.enable_N_60_1 ),
            .ltout(),
            .carryin(\eeprom.n4228 ),
            .carryout(\eeprom.n4229 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_4_lut_LC_20_17_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_4_lut_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_4_lut_LC_20_17_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_4_lut_LC_20_17_2  (
            .in0(N__24812),
            .in1(N__26712),
            .in2(N__21974),
            .in3(N__15395),
            .lcout(\eeprom.enable_N_60_2 ),
            .ltout(),
            .carryin(\eeprom.n4229 ),
            .carryout(\eeprom.n4230 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_5_lut_LC_20_17_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_5_lut_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_5_lut_LC_20_17_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_5_lut_LC_20_17_3  (
            .in0(N__25772),
            .in1(N__25319),
            .in2(N__26738),
            .in3(N__15392),
            .lcout(\eeprom.enable_N_60_3 ),
            .ltout(),
            .carryin(\eeprom.n4230 ),
            .carryout(\eeprom.n4231 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_6_lut_LC_20_17_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_6_lut_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_6_lut_LC_20_17_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_6_lut_LC_20_17_4  (
            .in0(N__24767),
            .in1(N__26716),
            .in2(N__21593),
            .in3(N__15389),
            .lcout(\eeprom.enable_N_60_4 ),
            .ltout(),
            .carryin(\eeprom.n4231 ),
            .carryout(\eeprom.n4232 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_7_lut_LC_20_17_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_7_lut_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_7_lut_LC_20_17_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_7_lut_LC_20_17_5  (
            .in0(N__25361),
            .in1(N__19001),
            .in2(N__26739),
            .in3(N__15386),
            .lcout(\eeprom.enable_N_60_5 ),
            .ltout(),
            .carryin(\eeprom.n4232 ),
            .carryout(\eeprom.n4233 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_8_lut_LC_20_17_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_8_lut_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_8_lut_LC_20_17_6 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_8_lut_LC_20_17_6  (
            .in0(N__29408),
            .in1(N__26720),
            .in2(N__29369),
            .in3(N__15383),
            .lcout(\eeprom.enable_N_60_6 ),
            .ltout(),
            .carryin(\eeprom.n4233 ),
            .carryout(\eeprom.n4234 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_9_lut_LC_20_17_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_9_lut_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_9_lut_LC_20_17_7 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_9_lut_LC_20_17_7  (
            .in0(N__15380),
            .in1(N__26740),
            .in2(N__15374),
            .in3(N__15365),
            .lcout(\eeprom.enable_N_60_7 ),
            .ltout(),
            .carryin(\eeprom.n4234 ),
            .carryout(\eeprom.n4235 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_10_lut_LC_20_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_10_lut_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_10_lut_LC_20_18_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_10_lut_LC_20_18_0  (
            .in0(N__15362),
            .in1(N__26731),
            .in2(N__15356),
            .in3(N__15347),
            .lcout(\eeprom.enable_N_60_8 ),
            .ltout(),
            .carryin(bfn_20_18_0_),
            .carryout(\eeprom.n4236 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_11_lut_LC_20_18_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_11_lut_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_11_lut_LC_20_18_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_2473_11_lut_LC_20_18_1  (
            .in0(N__15491),
            .in1(N__15500),
            .in2(N__26744),
            .in3(N__15344),
            .lcout(\eeprom.enable_N_60_9 ),
            .ltout(),
            .carryin(\eeprom.n4236 ),
            .carryout(\eeprom.n4237 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_12_lut_LC_20_18_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_12_lut_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_12_lut_LC_20_18_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_12_lut_LC_20_18_2  (
            .in0(N__15341),
            .in1(N__26735),
            .in2(N__15335),
            .in3(N__15326),
            .lcout(\eeprom.enable_N_60_10 ),
            .ltout(),
            .carryin(\eeprom.n4237 ),
            .carryout(\eeprom.n4238 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_13_lut_LC_20_18_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_13_lut_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_13_lut_LC_20_18_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_13_lut_LC_20_18_3  (
            .in0(N__15584),
            .in1(N__26741),
            .in2(N__15578),
            .in3(N__15569),
            .lcout(\eeprom.enable_N_60_11 ),
            .ltout(),
            .carryin(\eeprom.n4238 ),
            .carryout(\eeprom.n4239 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_14_lut_LC_20_18_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_14_lut_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_14_lut_LC_20_18_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_14_lut_LC_20_18_4  (
            .in0(N__15566),
            .in1(N__26736),
            .in2(N__15557),
            .in3(N__15545),
            .lcout(\eeprom.enable_N_60_12 ),
            .ltout(),
            .carryin(\eeprom.n4239 ),
            .carryout(\eeprom.n4240 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_15_lut_LC_20_18_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2473_15_lut_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_15_lut_LC_20_18_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \eeprom.rem_4_add_2473_15_lut_LC_20_18_5  (
            .in0(N__15542),
            .in1(N__26742),
            .in2(N__15536),
            .in3(N__15527),
            .lcout(\eeprom.enable_N_60_13 ),
            .ltout(),
            .carryin(\eeprom.n4240 ),
            .carryout(\eeprom.n4241 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2473_16_lut_LC_20_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2473_16_lut_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2473_16_lut_LC_20_18_6 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \eeprom.rem_4_add_2473_16_lut_LC_20_18_6  (
            .in0(N__26743),
            .in1(N__15524),
            .in2(N__15518),
            .in3(N__15503),
            .lcout(\eeprom.enable_N_60_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4723_1_lut_LC_20_18_7 .C_ON=1'b0;
    defparam \eeprom.i4723_1_lut_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4723_1_lut_LC_20_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.i4723_1_lut_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15499),
            .lcout(\eeprom.n5553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_2_lut_LC_20_19_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_2_lut_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_2_lut_LC_20_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_2_lut_LC_20_19_0  (
            .in0(_gnd_net_),
            .in1(N__29458),
            .in2(_gnd_net_),
            .in3(N__15473),
            .lcout(\eeprom.n3586 ),
            .ltout(),
            .carryin(bfn_20_19_0_),
            .carryout(\eeprom.n4205 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_3_lut_LC_20_19_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_3_lut_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_3_lut_LC_20_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_3_lut_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(N__28504),
            .in2(N__15470),
            .in3(N__15440),
            .lcout(\eeprom.n3585_adj_296 ),
            .ltout(),
            .carryin(\eeprom.n4205 ),
            .carryout(\eeprom.n4206 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_4_lut_LC_20_19_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_4_lut_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_4_lut_LC_20_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_4_lut_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15437),
            .in3(N__15398),
            .lcout(\eeprom.n3584 ),
            .ltout(),
            .carryin(\eeprom.n4206 ),
            .carryout(\eeprom.n4207 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_5_lut_LC_20_19_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_5_lut_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_5_lut_LC_20_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_5_lut_LC_20_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15884),
            .in3(N__15845),
            .lcout(\eeprom.n3583 ),
            .ltout(),
            .carryin(\eeprom.n4207 ),
            .carryout(\eeprom.n4208 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_6_lut_LC_20_19_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_6_lut_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_6_lut_LC_20_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_6_lut_LC_20_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15842),
            .in3(N__15803),
            .lcout(\eeprom.n3582 ),
            .ltout(),
            .carryin(\eeprom.n4208 ),
            .carryout(\eeprom.n4209 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_7_lut_LC_20_19_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_7_lut_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_7_lut_LC_20_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_7_lut_LC_20_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15800),
            .in3(N__15767),
            .lcout(\eeprom.n3581_adj_292 ),
            .ltout(),
            .carryin(\eeprom.n4209 ),
            .carryout(\eeprom.n4210 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_8_lut_LC_20_19_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_8_lut_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_8_lut_LC_20_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_8_lut_LC_20_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15764),
            .in3(N__15734),
            .lcout(\eeprom.n3580 ),
            .ltout(),
            .carryin(\eeprom.n4210 ),
            .carryout(\eeprom.n4211 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_9_lut_LC_20_19_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_9_lut_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_9_lut_LC_20_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_9_lut_LC_20_19_7  (
            .in0(_gnd_net_),
            .in1(N__28505),
            .in2(N__15731),
            .in3(N__15701),
            .lcout(\eeprom.n3579 ),
            .ltout(),
            .carryin(\eeprom.n4211 ),
            .carryout(\eeprom.n4212 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_10_lut_LC_20_20_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_10_lut_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_10_lut_LC_20_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_10_lut_LC_20_20_0  (
            .in0(_gnd_net_),
            .in1(N__28633),
            .in2(N__15698),
            .in3(N__15665),
            .lcout(\eeprom.n3578 ),
            .ltout(),
            .carryin(bfn_20_20_0_),
            .carryout(\eeprom.n4213 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_11_lut_LC_20_20_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_11_lut_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_11_lut_LC_20_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_11_lut_LC_20_20_1  (
            .in0(_gnd_net_),
            .in1(N__28644),
            .in2(N__15662),
            .in3(N__15626),
            .lcout(\eeprom.n3577 ),
            .ltout(),
            .carryin(\eeprom.n4213 ),
            .carryout(\eeprom.n4214 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_12_lut_LC_20_20_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_12_lut_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_12_lut_LC_20_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_12_lut_LC_20_20_2  (
            .in0(_gnd_net_),
            .in1(N__28634),
            .in2(N__15623),
            .in3(N__15587),
            .lcout(\eeprom.n3576 ),
            .ltout(),
            .carryin(\eeprom.n4214 ),
            .carryout(\eeprom.n4215 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_13_lut_LC_20_20_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_13_lut_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_13_lut_LC_20_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_13_lut_LC_20_20_3  (
            .in0(_gnd_net_),
            .in1(N__16128),
            .in2(N__28759),
            .in3(N__16094),
            .lcout(\eeprom.n3575 ),
            .ltout(),
            .carryin(\eeprom.n4215 ),
            .carryout(\eeprom.n4216 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_14_lut_LC_20_20_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_14_lut_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_14_lut_LC_20_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_14_lut_LC_20_20_4  (
            .in0(_gnd_net_),
            .in1(N__16090),
            .in2(N__28762),
            .in3(N__16067),
            .lcout(\eeprom.n3574 ),
            .ltout(),
            .carryin(\eeprom.n4216 ),
            .carryout(\eeprom.n4217 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_15_lut_LC_20_20_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_15_lut_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_15_lut_LC_20_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_15_lut_LC_20_20_5  (
            .in0(_gnd_net_),
            .in1(N__16063),
            .in2(N__28760),
            .in3(N__16034),
            .lcout(\eeprom.n3573 ),
            .ltout(),
            .carryin(\eeprom.n4217 ),
            .carryout(\eeprom.n4218 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_16_lut_LC_20_20_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_16_lut_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_16_lut_LC_20_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_16_lut_LC_20_20_6  (
            .in0(_gnd_net_),
            .in1(N__16030),
            .in2(N__28763),
            .in3(N__16007),
            .lcout(\eeprom.n3572 ),
            .ltout(),
            .carryin(\eeprom.n4218 ),
            .carryout(\eeprom.n4219 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_17_lut_LC_20_20_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_17_lut_LC_20_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_17_lut_LC_20_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_17_lut_LC_20_20_7  (
            .in0(_gnd_net_),
            .in1(N__16004),
            .in2(N__28761),
            .in3(N__15971),
            .lcout(\eeprom.n3571 ),
            .ltout(),
            .carryin(\eeprom.n4219 ),
            .carryout(\eeprom.n4220 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_18_lut_LC_20_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_18_lut_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_18_lut_LC_20_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_18_lut_LC_20_21_0  (
            .in0(_gnd_net_),
            .in1(N__15968),
            .in2(N__28554),
            .in3(N__15938),
            .lcout(\eeprom.n3570 ),
            .ltout(),
            .carryin(bfn_20_21_0_),
            .carryout(\eeprom.n4221 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_19_lut_LC_20_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_19_lut_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_19_lut_LC_20_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_19_lut_LC_20_21_1  (
            .in0(_gnd_net_),
            .in1(N__19074),
            .in2(N__28557),
            .in3(N__15923),
            .lcout(\eeprom.n3569 ),
            .ltout(),
            .carryin(\eeprom.n4221 ),
            .carryout(\eeprom.n4222 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_20_lut_LC_20_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_20_lut_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_20_lut_LC_20_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_20_lut_LC_20_21_2  (
            .in0(_gnd_net_),
            .in1(N__15916),
            .in2(N__28555),
            .in3(N__16490),
            .lcout(\eeprom.n3568 ),
            .ltout(),
            .carryin(\eeprom.n4222 ),
            .carryout(\eeprom.n4223 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_21_lut_LC_20_21_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_21_lut_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_21_lut_LC_20_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_21_lut_LC_20_21_3  (
            .in0(_gnd_net_),
            .in1(N__16485),
            .in2(N__28558),
            .in3(N__16457),
            .lcout(\eeprom.n3567 ),
            .ltout(),
            .carryin(\eeprom.n4223 ),
            .carryout(\eeprom.n4224 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_22_lut_LC_20_21_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_22_lut_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_22_lut_LC_20_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_22_lut_LC_20_21_4  (
            .in0(_gnd_net_),
            .in1(N__28428),
            .in2(N__16454),
            .in3(N__16427),
            .lcout(\eeprom.n3566 ),
            .ltout(),
            .carryin(\eeprom.n4224 ),
            .carryout(\eeprom.n4225 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_23_lut_LC_20_21_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_23_lut_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_23_lut_LC_20_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_23_lut_LC_20_21_5  (
            .in0(_gnd_net_),
            .in1(N__28418),
            .in2(N__16420),
            .in3(N__16394),
            .lcout(\eeprom.n3565 ),
            .ltout(),
            .carryin(\eeprom.n4225 ),
            .carryout(\eeprom.n4226 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_24_lut_LC_20_21_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_2357_24_lut_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_24_lut_LC_20_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_2357_24_lut_LC_20_21_6  (
            .in0(_gnd_net_),
            .in1(N__16391),
            .in2(N__28556),
            .in3(N__16358),
            .lcout(\eeprom.n3564 ),
            .ltout(),
            .carryin(\eeprom.n4226 ),
            .carryout(\eeprom.n4227 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_2357_25_lut_LC_20_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_2357_25_lut_LC_20_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_2357_25_lut_LC_20_21_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_2357_25_lut_LC_20_21_7  (
            .in0(N__28429),
            .in1(N__16355),
            .in2(N__16334),
            .in3(N__16214),
            .lcout(\eeprom.n5355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2242_3_lut_LC_20_22_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2242_3_lut_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2242_3_lut_LC_20_22_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2242_3_lut_LC_20_22_0  (
            .in0(_gnd_net_),
            .in1(N__16199),
            .in2(N__17151),
            .in3(N__17659),
            .lcout(\eeprom.n3414 ),
            .ltout(\eeprom.n3414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_LC_20_22_1 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_LC_20_22_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_LC_20_22_1  (
            .in0(_gnd_net_),
            .in1(N__16155),
            .in2(N__16136),
            .in3(N__16617),
            .lcout(),
            .ltout(\eeprom.n5291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_LC_20_22_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_LC_20_22_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_LC_20_22_2  (
            .in0(N__16656),
            .in1(N__23422),
            .in2(N__16133),
            .in3(N__17201),
            .lcout(),
            .ltout(\eeprom.n4824_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_LC_20_22_3 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_LC_20_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_LC_20_22_3  (
            .in0(N__16737),
            .in1(N__19254),
            .in2(N__16718),
            .in3(N__16714),
            .lcout(\eeprom.n28_adj_261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2246_3_lut_LC_20_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2246_3_lut_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2246_3_lut_LC_20_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i2246_3_lut_LC_20_22_5  (
            .in0(N__22670),
            .in1(N__16676),
            .in2(_gnd_net_),
            .in3(N__17115),
            .lcout(\eeprom.n3418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2244_3_lut_LC_20_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2244_3_lut_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2244_3_lut_LC_20_22_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2244_3_lut_LC_20_22_6  (
            .in0(_gnd_net_),
            .in1(N__16637),
            .in2(N__17150),
            .in3(N__16952),
            .lcout(\eeprom.n3416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2243_3_lut_LC_20_22_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2243_3_lut_LC_20_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2243_3_lut_LC_20_22_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2243_3_lut_LC_20_22_7  (
            .in0(_gnd_net_),
            .in1(N__16906),
            .in2(N__16598),
            .in3(N__17119),
            .lcout(\eeprom.n3415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_108_LC_20_23_1 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_108_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_108_LC_20_23_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_108_LC_20_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17655),
            .in3(N__16572),
            .lcout(\eeprom.n5313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2231_3_lut_LC_20_23_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2231_3_lut_LC_20_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2231_3_lut_LC_20_23_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2231_3_lut_LC_20_23_2  (
            .in0(_gnd_net_),
            .in1(N__16819),
            .in2(N__16556),
            .in3(N__17125),
            .lcout(\eeprom.n3403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2174_3_lut_LC_20_23_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2174_3_lut_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2174_3_lut_LC_20_23_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2174_3_lut_LC_20_23_3  (
            .in0(_gnd_net_),
            .in1(N__17398),
            .in2(N__16541),
            .in3(N__17740),
            .lcout(\eeprom.n3314 ),
            .ltout(\eeprom.n3314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2241_3_lut_LC_20_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2241_3_lut_LC_20_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2241_3_lut_LC_20_23_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2241_3_lut_LC_20_23_4  (
            .in0(_gnd_net_),
            .in1(N__16526),
            .in2(N__16514),
            .in3(N__17123),
            .lcout(\eeprom.n3413 ),
            .ltout(\eeprom.n3413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_12_LC_20_23_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_12_LC_20_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_12_LC_20_23_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_12_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17231),
            .in3(N__17217),
            .lcout(\eeprom.n5289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2170_3_lut_LC_20_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2170_3_lut_LC_20_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2170_3_lut_LC_20_23_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i2170_3_lut_LC_20_23_6  (
            .in0(_gnd_net_),
            .in1(N__17195),
            .in2(N__17773),
            .in3(N__18223),
            .lcout(\eeprom.n3310 ),
            .ltout(\eeprom.n3310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2237_3_lut_LC_20_23_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2237_3_lut_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2237_3_lut_LC_20_23_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_i2237_3_lut_LC_20_23_7  (
            .in0(N__17124),
            .in1(_gnd_net_),
            .in2(N__17048),
            .in3(N__17045),
            .lcout(\eeprom.n3409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2176_3_lut_LC_20_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2176_3_lut_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2176_3_lut_LC_20_24_0 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i2176_3_lut_LC_20_24_0  (
            .in0(N__17006),
            .in1(N__17320),
            .in2(N__17771),
            .in3(_gnd_net_),
            .lcout(\eeprom.n3316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2177_3_lut_LC_20_24_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2177_3_lut_LC_20_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2177_3_lut_LC_20_24_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \eeprom.rem_4_i2177_3_lut_LC_20_24_3  (
            .in0(N__16994),
            .in1(N__17735),
            .in2(_gnd_net_),
            .in3(N__16964),
            .lcout(\eeprom.n3317 ),
            .ltout(\eeprom.n3317_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_109_LC_20_24_4 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_109_LC_20_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_109_LC_20_24_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_109_LC_20_24_4  (
            .in0(_gnd_net_),
            .in1(N__16924),
            .in2(N__16913),
            .in3(N__16905),
            .lcout(),
            .ltout(\eeprom.n5315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_110_LC_20_24_5 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_110_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_110_LC_20_24_5 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_110_LC_20_24_5  (
            .in0(N__22666),
            .in1(N__16879),
            .in2(N__16856),
            .in3(N__16853),
            .lcout(),
            .ltout(\eeprom.n4820_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_112_LC_20_24_6 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_112_LC_20_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_112_LC_20_24_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_112_LC_20_24_6  (
            .in0(N__16836),
            .in1(N__16809),
            .in2(N__16793),
            .in3(N__16789),
            .lcout(\eeprom.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2175_3_lut_LC_20_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2175_3_lut_LC_20_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2175_3_lut_LC_20_24_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2175_3_lut_LC_20_24_7  (
            .in0(_gnd_net_),
            .in1(N__17491),
            .in2(N__17801),
            .in3(N__17731),
            .lcout(\eeprom.n3315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2105_3_lut_LC_20_25_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2105_3_lut_LC_20_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2105_3_lut_LC_20_25_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2105_3_lut_LC_20_25_0  (
            .in0(_gnd_net_),
            .in1(N__17630),
            .in2(N__17600),
            .in3(N__17920),
            .lcout(\eeprom.n3213 ),
            .ltout(\eeprom.n3213_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_31_LC_20_25_1 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_31_LC_20_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_31_LC_20_25_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_31_LC_20_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17561),
            .in3(N__17388),
            .lcout(\eeprom.n5205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2106_3_lut_LC_20_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2106_3_lut_LC_20_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2106_3_lut_LC_20_25_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i2106_3_lut_LC_20_25_2  (
            .in0(_gnd_net_),
            .in1(N__17558),
            .in2(N__17546),
            .in3(N__17919),
            .lcout(\eeprom.n3214 ),
            .ltout(\eeprom.n3214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_32_LC_20_25_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_32_LC_20_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_32_LC_20_25_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_32_LC_20_25_3  (
            .in0(N__17484),
            .in1(N__17319),
            .in2(N__17465),
            .in3(N__17462),
            .lcout(\eeprom.n5209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2107_3_lut_LC_20_25_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2107_3_lut_LC_20_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2107_3_lut_LC_20_25_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2107_3_lut_LC_20_25_4  (
            .in0(_gnd_net_),
            .in1(N__17447),
            .in2(N__17417),
            .in3(N__17915),
            .lcout(\eeprom.n3215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2109_3_lut_LC_20_25_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2109_3_lut_LC_20_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2109_3_lut_LC_20_25_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i2109_3_lut_LC_20_25_5  (
            .in0(N__17372),
            .in1(_gnd_net_),
            .in2(N__17948),
            .in3(N__17360),
            .lcout(\eeprom.n3217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2100_3_lut_LC_20_25_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2100_3_lut_LC_20_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2100_3_lut_LC_20_25_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2100_3_lut_LC_20_25_6  (
            .in0(_gnd_net_),
            .in1(N__17300),
            .in2(N__17267),
            .in3(N__17921),
            .lcout(\eeprom.n3208 ),
            .ltout(\eeprom.n3208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_37_LC_20_25_7 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_37_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_37_LC_20_25_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_37_LC_20_25_7  (
            .in0(N__18216),
            .in1(N__17820),
            .in2(N__18197),
            .in3(N__18193),
            .lcout(\eeprom.n26_adj_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1969_3_lut_LC_20_26_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1969_3_lut_LC_20_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1969_3_lut_LC_20_26_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1969_3_lut_LC_20_26_0  (
            .in0(_gnd_net_),
            .in1(N__18574),
            .in2(N__18560),
            .in3(N__18723),
            .lcout(\eeprom.n3013 ),
            .ltout(\eeprom.n3013_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2036_3_lut_LC_20_26_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2036_3_lut_LC_20_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2036_3_lut_LC_20_26_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i2036_3_lut_LC_20_26_1  (
            .in0(N__18161),
            .in1(_gnd_net_),
            .in2(N__18149),
            .in3(N__18144),
            .lcout(\eeprom.n3112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_2_lut_LC_20_26_2 .C_ON=1'b0;
    defparam \eeprom.i6_2_lut_LC_20_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_2_lut_LC_20_26_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i6_2_lut_LC_20_26_2  (
            .in0(_gnd_net_),
            .in1(N__19434),
            .in2(_gnd_net_),
            .in3(N__19317),
            .lcout(\eeprom.n18_adj_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1967_3_lut_LC_20_26_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1967_3_lut_LC_20_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1967_3_lut_LC_20_26_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1967_3_lut_LC_20_26_3  (
            .in0(N__19318),
            .in1(_gnd_net_),
            .in2(N__18760),
            .in3(N__18518),
            .lcout(\eeprom.n3011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_LC_20_26_4 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_LC_20_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_LC_20_26_4 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \eeprom.i3_4_lut_LC_20_26_4  (
            .in0(N__22465),
            .in1(N__18849),
            .in2(N__19474),
            .in3(N__17990),
            .lcout(\eeprom.n15_adj_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2101_3_lut_LC_20_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2101_3_lut_LC_20_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2101_3_lut_LC_20_26_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i2101_3_lut_LC_20_26_5  (
            .in0(_gnd_net_),
            .in1(N__17979),
            .in2(N__17955),
            .in3(N__17849),
            .lcout(\eeprom.n3209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1904_3_lut_LC_20_27_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1904_3_lut_LC_20_27_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1904_3_lut_LC_20_27_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1904_3_lut_LC_20_27_0  (
            .in0(_gnd_net_),
            .in1(N__20960),
            .in2(N__19400),
            .in3(N__19643),
            .lcout(\eeprom.n2916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1898_3_lut_LC_20_27_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1898_3_lut_LC_20_27_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1898_3_lut_LC_20_27_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1898_3_lut_LC_20_27_1  (
            .in0(_gnd_net_),
            .in1(N__19535),
            .in2(N__19672),
            .in3(N__21365),
            .lcout(\eeprom.n2910 ),
            .ltout(\eeprom.n2910_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_67_LC_20_27_2 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_67_LC_20_27_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_67_LC_20_27_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_67_LC_20_27_2  (
            .in0(N__19588),
            .in1(N__19790),
            .in2(N__18302),
            .in3(N__18299),
            .lcout(),
            .ltout(\eeprom.n22_adj_331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i11_4_lut_adj_68_LC_20_27_3 .C_ON=1'b0;
    defparam \eeprom.i11_4_lut_adj_68_LC_20_27_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i11_4_lut_adj_68_LC_20_27_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i11_4_lut_adj_68_LC_20_27_3  (
            .in0(N__18426),
            .in1(N__18459),
            .in2(N__18293),
            .in3(N__18290),
            .lcout(\eeprom.n2935 ),
            .ltout(\eeprom.n2935_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1971_3_lut_LC_20_27_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1971_3_lut_LC_20_27_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1971_3_lut_LC_20_27_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1971_3_lut_LC_20_27_4  (
            .in0(N__18311),
            .in1(_gnd_net_),
            .in2(N__18284),
            .in3(N__18331),
            .lcout(\eeprom.n3015 ),
            .ltout(\eeprom.n3015_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_76_LC_20_27_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_76_LC_20_27_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_76_LC_20_27_5 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \eeprom.i1_2_lut_adj_76_LC_20_27_5  (
            .in0(_gnd_net_),
            .in1(N__18250),
            .in2(N__18239),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1894_3_lut_LC_20_27_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1894_3_lut_LC_20_27_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1894_3_lut_LC_20_27_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1894_3_lut_LC_20_27_6  (
            .in0(_gnd_net_),
            .in1(N__21163),
            .in2(N__19499),
            .in3(N__19644),
            .lcout(\eeprom.n2906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1896_3_lut_LC_20_27_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1896_3_lut_LC_20_27_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1896_3_lut_LC_20_27_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1896_3_lut_LC_20_27_7  (
            .in0(_gnd_net_),
            .in1(N__19514),
            .in2(N__19673),
            .in3(N__21275),
            .lcout(\eeprom.n2908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_LC_20_28_0 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_LC_20_28_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_LC_20_28_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_LC_20_28_0  (
            .in0(N__21273),
            .in1(N__21210),
            .in2(N__21109),
            .in3(N__21074),
            .lcout(),
            .ltout(\eeprom.n18_adj_290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_adj_29_LC_20_28_1 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_adj_29_LC_20_28_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_adj_29_LC_20_28_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_adj_29_LC_20_28_1  (
            .in0(N__21364),
            .in1(N__21024),
            .in2(N__18230),
            .in3(N__21401),
            .lcout(),
            .ltout(\eeprom.n20_adj_291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i10_4_lut_adj_30_LC_20_28_2 .C_ON=1'b0;
    defparam \eeprom.i10_4_lut_adj_30_LC_20_28_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i10_4_lut_adj_30_LC_20_28_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i10_4_lut_adj_30_LC_20_28_2  (
            .in0(N__19298),
            .in1(N__21310),
            .in2(N__18227),
            .in3(N__21159),
            .lcout(\eeprom.n2836 ),
            .ltout(\eeprom.n2836_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1903_3_lut_LC_20_28_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1903_3_lut_LC_20_28_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1903_3_lut_LC_20_28_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1903_3_lut_LC_20_28_3  (
            .in0(N__19388),
            .in1(_gnd_net_),
            .in2(N__18407),
            .in3(N__20900),
            .lcout(\eeprom.n2915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1897_3_lut_LC_20_28_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1897_3_lut_LC_20_28_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1897_3_lut_LC_20_28_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1897_3_lut_LC_20_28_4  (
            .in0(_gnd_net_),
            .in1(N__21311),
            .in2(N__19526),
            .in3(N__19642),
            .lcout(\eeprom.n2909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1905_3_lut_LC_20_28_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1905_3_lut_LC_20_28_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1905_3_lut_LC_20_28_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \eeprom.rem_4_i1905_3_lut_LC_20_28_5  (
            .in0(N__20990),
            .in1(N__19409),
            .in2(N__19671),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1901_3_lut_LC_20_28_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1901_3_lut_LC_20_28_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1901_3_lut_LC_20_28_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i1901_3_lut_LC_20_28_6  (
            .in0(N__19364),
            .in1(_gnd_net_),
            .in2(N__20819),
            .in3(N__19638),
            .lcout(\eeprom.n2913 ),
            .ltout(\eeprom.n2913_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_33_LC_20_28_7 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_33_LC_20_28_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_33_LC_20_28_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_33_LC_20_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18404),
            .in3(N__18609),
            .lcout(\eeprom.n5297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_2_lut_LC_20_29_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_2_lut_LC_20_29_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_2_lut_LC_20_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_2_lut_LC_20_29_0  (
            .in0(_gnd_net_),
            .in1(N__22464),
            .in2(_gnd_net_),
            .in3(N__18383),
            .lcout(\eeprom.n2986 ),
            .ltout(),
            .carryin(bfn_20_29_0_),
            .carryout(\eeprom.n4088 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_3_lut_LC_20_29_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_3_lut_LC_20_29_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_3_lut_LC_20_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_3_lut_LC_20_29_1  (
            .in0(_gnd_net_),
            .in1(N__19473),
            .in2(N__28559),
            .in3(N__18371),
            .lcout(\eeprom.n2985 ),
            .ltout(),
            .carryin(\eeprom.n4088 ),
            .carryout(\eeprom.n4089 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_4_lut_LC_20_29_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_4_lut_LC_20_29_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_4_lut_LC_20_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_4_lut_LC_20_29_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18368),
            .in3(N__18338),
            .lcout(\eeprom.n2984 ),
            .ltout(),
            .carryin(\eeprom.n4089 ),
            .carryout(\eeprom.n4090 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_5_lut_LC_20_29_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_5_lut_LC_20_29_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_5_lut_LC_20_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_5_lut_LC_20_29_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18335),
            .in3(N__18620),
            .lcout(\eeprom.n2983 ),
            .ltout(),
            .carryin(\eeprom.n4090 ),
            .carryout(\eeprom.n4091 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_6_lut_LC_20_29_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_6_lut_LC_20_29_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_6_lut_LC_20_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_6_lut_LC_20_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18616),
            .in3(N__18581),
            .lcout(\eeprom.n2982 ),
            .ltout(),
            .carryin(\eeprom.n4091 ),
            .carryout(\eeprom.n4092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_7_lut_LC_20_29_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_7_lut_LC_20_29_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_7_lut_LC_20_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_7_lut_LC_20_29_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18578),
            .in3(N__18548),
            .lcout(\eeprom.n2981 ),
            .ltout(),
            .carryin(\eeprom.n4092 ),
            .carryout(\eeprom.n4093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_8_lut_LC_20_29_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_8_lut_LC_20_29_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_8_lut_LC_20_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_8_lut_LC_20_29_6  (
            .in0(_gnd_net_),
            .in1(N__18544),
            .in2(_gnd_net_),
            .in3(N__18521),
            .lcout(\eeprom.n2980 ),
            .ltout(),
            .carryin(\eeprom.n4093 ),
            .carryout(\eeprom.n4094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_9_lut_LC_20_29_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_9_lut_LC_20_29_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_9_lut_LC_20_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_9_lut_LC_20_29_7  (
            .in0(_gnd_net_),
            .in1(N__28433),
            .in2(N__19325),
            .in3(N__18506),
            .lcout(\eeprom.n2979 ),
            .ltout(),
            .carryin(\eeprom.n4094 ),
            .carryout(\eeprom.n4095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_10_lut_LC_20_30_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_10_lut_LC_20_30_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_10_lut_LC_20_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_10_lut_LC_20_30_0  (
            .in0(_gnd_net_),
            .in1(N__19447),
            .in2(N__28919),
            .in3(N__18497),
            .lcout(\eeprom.n2978 ),
            .ltout(),
            .carryin(bfn_20_30_0_),
            .carryout(\eeprom.n4096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_11_lut_LC_20_30_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_11_lut_LC_20_30_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_11_lut_LC_20_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_11_lut_LC_20_30_1  (
            .in0(_gnd_net_),
            .in1(N__18493),
            .in2(N__28923),
            .in3(N__18464),
            .lcout(\eeprom.n2977 ),
            .ltout(),
            .carryin(\eeprom.n4096 ),
            .carryout(\eeprom.n4097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_12_lut_LC_20_30_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_12_lut_LC_20_30_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_12_lut_LC_20_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_12_lut_LC_20_30_2  (
            .in0(_gnd_net_),
            .in1(N__18460),
            .in2(N__28920),
            .in3(N__18431),
            .lcout(\eeprom.n2976 ),
            .ltout(),
            .carryin(\eeprom.n4097 ),
            .carryout(\eeprom.n4098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_13_lut_LC_20_30_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_13_lut_LC_20_30_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_13_lut_LC_20_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_13_lut_LC_20_30_3  (
            .in0(_gnd_net_),
            .in1(N__18428),
            .in2(N__28924),
            .in3(N__18875),
            .lcout(\eeprom.n2975 ),
            .ltout(),
            .carryin(\eeprom.n4098 ),
            .carryout(\eeprom.n4099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_14_lut_LC_20_30_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_14_lut_LC_20_30_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_14_lut_LC_20_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_14_lut_LC_20_30_4  (
            .in0(_gnd_net_),
            .in1(N__19578),
            .in2(N__28921),
            .in3(N__18863),
            .lcout(\eeprom.n2974 ),
            .ltout(),
            .carryin(\eeprom.n4099 ),
            .carryout(\eeprom.n4100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_15_lut_LC_20_30_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_15_lut_LC_20_30_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_15_lut_LC_20_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_15_lut_LC_20_30_5  (
            .in0(_gnd_net_),
            .in1(N__18856),
            .in2(N__28925),
            .in3(N__18827),
            .lcout(\eeprom.n2973 ),
            .ltout(),
            .carryin(\eeprom.n4100 ),
            .carryout(\eeprom.n4101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_16_lut_LC_20_30_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_16_lut_LC_20_30_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_16_lut_LC_20_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_16_lut_LC_20_30_6  (
            .in0(_gnd_net_),
            .in1(N__19741),
            .in2(N__28922),
            .in3(N__18812),
            .lcout(\eeprom.n2972 ),
            .ltout(),
            .carryin(\eeprom.n4101 ),
            .carryout(\eeprom.n4102 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_17_lut_LC_20_30_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_17_lut_LC_20_30_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_17_lut_LC_20_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_17_lut_LC_20_30_7  (
            .in0(_gnd_net_),
            .in1(N__19771),
            .in2(N__28926),
            .in3(N__18803),
            .lcout(\eeprom.n2971 ),
            .ltout(),
            .carryin(\eeprom.n4102 ),
            .carryout(\eeprom.n4103 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_18_lut_LC_20_31_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1955_18_lut_LC_20_31_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_18_lut_LC_20_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1955_18_lut_LC_20_31_0  (
            .in0(_gnd_net_),
            .in1(N__19714),
            .in2(N__28927),
            .in3(N__18788),
            .lcout(\eeprom.n2970 ),
            .ltout(),
            .carryin(bfn_20_31_0_),
            .carryout(\eeprom.n4104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1955_19_lut_LC_20_31_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1955_19_lut_LC_20_31_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1955_19_lut_LC_20_31_1 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1955_19_lut_LC_20_31_1  (
            .in0(N__28440),
            .in1(N__19802),
            .in2(N__18785),
            .in3(N__18677),
            .lcout(\eeprom.n3001 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_41_LC_21_17_0 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_41_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_41_LC_21_17_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \eeprom.i1_3_lut_adj_41_LC_21_17_0  (
            .in0(N__18653),
            .in1(N__18647),
            .in2(_gnd_net_),
            .in3(N__18641),
            .lcout(),
            .ltout(\eeprom.n4847_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_45_LC_21_17_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_45_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_45_LC_21_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_45_LC_21_17_1  (
            .in0(N__18635),
            .in1(N__18626),
            .in2(N__18983),
            .in3(N__18980),
            .lcout(),
            .ltout(\eeprom.n4853_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_46_LC_21_17_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_46_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_46_LC_21_17_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_46_LC_21_17_2  (
            .in0(N__18974),
            .in1(N__18968),
            .in2(N__18962),
            .in3(N__18959),
            .lcout(),
            .ltout(\eeprom.n4859_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_47_LC_21_17_3 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_47_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_47_LC_21_17_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i1_4_lut_adj_47_LC_21_17_3  (
            .in0(N__18953),
            .in1(N__18947),
            .in2(N__18941),
            .in3(N__18938),
            .lcout(\eeprom.n4865 ),
            .ltout(\eeprom.n4865_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4699_4_lut_LC_21_17_4 .C_ON=1'b0;
    defparam \eeprom.i4699_4_lut_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4699_4_lut_LC_21_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \eeprom.i4699_4_lut_LC_21_17_4  (
            .in0(N__18925),
            .in1(N__18904),
            .in2(N__18932),
            .in3(N__18916),
            .lcout(),
            .ltout(\eeprom.enable_N_59_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rw_16_LC_21_17_5 .C_ON=1'b0;
    defparam \eeprom.rw_16_LC_21_17_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.rw_16_LC_21_17_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \eeprom.rw_16_LC_21_17_5  (
            .in0(N__27895),
            .in1(_gnd_net_),
            .in2(N__18929),
            .in3(_gnd_net_),
            .lcout(rw),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29860),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.enable_14_LC_21_17_6 .C_ON=1'b0;
    defparam \eeprom.enable_14_LC_21_17_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.enable_14_LC_21_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \eeprom.enable_14_LC_21_17_6  (
            .in0(N__18926),
            .in1(N__18917),
            .in2(N__18908),
            .in3(N__18893),
            .lcout(\eeprom.enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29860),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1423_3_lut_LC_21_18_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1423_3_lut_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1423_3_lut_LC_21_18_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1423_3_lut_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__22730),
            .in2(N__22700),
            .in3(N__23139),
            .lcout(\eeprom.n2211 ),
            .ltout(\eeprom.n2211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1490_3_lut_LC_21_18_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1490_3_lut_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1490_3_lut_LC_21_18_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1490_3_lut_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__19820),
            .in2(N__18887),
            .in3(N__21734),
            .lcout(\eeprom.n2310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4676_3_lut_LC_21_18_2 .C_ON=1'b0;
    defparam \eeprom.i4676_3_lut_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4676_3_lut_LC_21_18_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.i4676_3_lut_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__22819),
            .in2(N__22844),
            .in3(N__23137),
            .lcout(\eeprom.n2215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1430_3_lut_LC_21_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1430_3_lut_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1430_3_lut_LC_21_18_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1430_3_lut_LC_21_18_6  (
            .in0(N__22373),
            .in1(N__24638),
            .in2(_gnd_net_),
            .in3(N__23138),
            .lcout(\eeprom.n2218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1493_3_lut_LC_21_19_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1493_3_lut_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1493_3_lut_LC_21_19_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1493_3_lut_LC_21_19_1  (
            .in0(_gnd_net_),
            .in1(N__19855),
            .in2(N__19841),
            .in3(N__21722),
            .lcout(\eeprom.n2313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1495_3_lut_LC_21_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1495_3_lut_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1495_3_lut_LC_21_19_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1495_3_lut_LC_21_19_3  (
            .in0(_gnd_net_),
            .in1(N__19889),
            .in2(N__19991),
            .in3(N__21723),
            .lcout(\eeprom.n2315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1426_3_lut_LC_21_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1426_3_lut_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1426_3_lut_LC_21_19_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1426_3_lut_LC_21_19_4  (
            .in0(_gnd_net_),
            .in1(N__22793),
            .in2(N__23315),
            .in3(N__23147),
            .lcout(\eeprom.n2214 ),
            .ltout(\eeprom.n2214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_52_LC_21_19_5 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_52_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_52_LC_21_19_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_52_LC_21_19_5  (
            .in0(N__20226),
            .in1(N__19873),
            .in2(N__19004),
            .in3(N__19983),
            .lcout(\eeprom.n5045 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1497_3_lut_LC_21_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1497_3_lut_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1497_3_lut_LC_21_19_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1497_3_lut_LC_21_19_6  (
            .in0(_gnd_net_),
            .in1(N__19907),
            .in2(N__21738),
            .in3(N__19955),
            .lcout(\eeprom.n2317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i6_3_lut_LC_21_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i6_3_lut_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i6_3_lut_LC_21_19_7 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i6_3_lut_LC_21_19_7  (
            .in0(N__25802),
            .in1(N__29206),
            .in2(_gnd_net_),
            .in3(N__25360),
            .lcout(\eeprom.n3720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_2_lut_LC_21_20_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_2_lut_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_2_lut_LC_21_20_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1553_2_lut_LC_21_20_0  (
            .in0(N__24602),
            .in1(N__24601),
            .in2(N__20319),
            .in3(N__18992),
            .lcout(\eeprom.n2418 ),
            .ltout(),
            .carryin(bfn_21_20_0_),
            .carryout(\eeprom.n4007 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_3_lut_LC_21_20_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_3_lut_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_3_lut_LC_21_20_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1553_3_lut_LC_21_20_1  (
            .in0(N__20108),
            .in1(N__20107),
            .in2(N__20367),
            .in3(N__18989),
            .lcout(\eeprom.n2417 ),
            .ltout(),
            .carryin(\eeprom.n4007 ),
            .carryout(\eeprom.n4008 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_4_lut_LC_21_20_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_4_lut_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_4_lut_LC_21_20_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1553_4_lut_LC_21_20_2  (
            .in0(N__20147),
            .in1(N__20146),
            .in2(N__20320),
            .in3(N__18986),
            .lcout(\eeprom.n2416 ),
            .ltout(),
            .carryin(\eeprom.n4008 ),
            .carryout(\eeprom.n4009 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_5_lut_LC_21_20_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_5_lut_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_5_lut_LC_21_20_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1553_5_lut_LC_21_20_3  (
            .in0(N__20164),
            .in1(N__20165),
            .in2(N__20323),
            .in3(N__19031),
            .lcout(\eeprom.n2415 ),
            .ltout(),
            .carryin(\eeprom.n4009 ),
            .carryout(\eeprom.n4010 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_6_lut_LC_21_20_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_6_lut_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_6_lut_LC_21_20_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1553_6_lut_LC_21_20_4  (
            .in0(N__20062),
            .in1(N__20061),
            .in2(N__20321),
            .in3(N__19028),
            .lcout(\eeprom.n2414 ),
            .ltout(),
            .carryin(\eeprom.n4010 ),
            .carryout(\eeprom.n4011 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_7_lut_LC_21_20_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_7_lut_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_7_lut_LC_21_20_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1553_7_lut_LC_21_20_5  (
            .in0(N__20128),
            .in1(N__20127),
            .in2(N__20324),
            .in3(N__19025),
            .lcout(\eeprom.n2413 ),
            .ltout(),
            .carryin(\eeprom.n4011 ),
            .carryout(\eeprom.n4012 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_8_lut_LC_21_20_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_8_lut_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_8_lut_LC_21_20_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1553_8_lut_LC_21_20_6  (
            .in0(N__20042),
            .in1(N__20041),
            .in2(N__20322),
            .in3(N__19022),
            .lcout(\eeprom.n2412 ),
            .ltout(),
            .carryin(\eeprom.n4012 ),
            .carryout(\eeprom.n4013 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_9_lut_LC_21_20_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_9_lut_LC_21_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_9_lut_LC_21_20_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1553_9_lut_LC_21_20_7  (
            .in0(N__20405),
            .in1(N__20404),
            .in2(N__20368),
            .in3(N__19019),
            .lcout(\eeprom.n2411 ),
            .ltout(),
            .carryin(\eeprom.n4013 ),
            .carryout(\eeprom.n4014 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_10_lut_LC_21_21_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_10_lut_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_10_lut_LC_21_21_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1553_10_lut_LC_21_21_0  (
            .in0(N__20273),
            .in1(N__20272),
            .in2(N__20369),
            .in3(N__19016),
            .lcout(\eeprom.n2410 ),
            .ltout(),
            .carryin(bfn_21_21_0_),
            .carryout(\eeprom.n4015 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_11_lut_LC_21_21_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_11_lut_LC_21_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_11_lut_LC_21_21_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1553_11_lut_LC_21_21_1  (
            .in0(N__20087),
            .in1(N__20086),
            .in2(N__20371),
            .in3(N__19013),
            .lcout(\eeprom.n2409 ),
            .ltout(),
            .carryin(\eeprom.n4015 ),
            .carryout(\eeprom.n4016 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_12_lut_LC_21_21_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1553_12_lut_LC_21_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_12_lut_LC_21_21_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1553_12_lut_LC_21_21_2  (
            .in0(N__20009),
            .in1(N__20008),
            .in2(N__20370),
            .in3(N__19010),
            .lcout(\eeprom.n2408 ),
            .ltout(),
            .carryin(\eeprom.n4016 ),
            .carryout(\eeprom.n4017 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1553_13_lut_LC_21_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1553_13_lut_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1553_13_lut_LC_21_21_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1553_13_lut_LC_21_21_3  (
            .in0(N__20428),
            .in1(N__20429),
            .in2(N__20372),
            .in3(N__19007),
            .lcout(\eeprom.n2407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i2298_3_lut_LC_21_22_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i2298_3_lut_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i2298_3_lut_LC_21_22_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i2298_3_lut_LC_21_22_0  (
            .in0(_gnd_net_),
            .in1(N__19258),
            .in2(N__19238),
            .in3(N__19207),
            .lcout(\eeprom.n3502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1627_3_lut_LC_21_22_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1627_3_lut_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1627_3_lut_LC_21_22_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1627_3_lut_LC_21_22_1  (
            .in0(_gnd_net_),
            .in1(N__20582),
            .in2(N__20558),
            .in3(N__23486),
            .lcout(\eeprom.n2511 ),
            .ltout(\eeprom.n2511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1694_3_lut_LC_21_22_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1694_3_lut_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1694_3_lut_LC_21_22_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1694_3_lut_LC_21_22_2  (
            .in0(_gnd_net_),
            .in1(N__23969),
            .in2(N__19055),
            .in3(N__24434),
            .lcout(\eeprom.n2610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1702_3_lut_LC_21_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1702_3_lut_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1702_3_lut_LC_21_22_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1702_3_lut_LC_21_22_4  (
            .in0(N__23723),
            .in1(N__24320),
            .in2(_gnd_net_),
            .in3(N__24433),
            .lcout(\eeprom.n2618 ),
            .ltout(\eeprom.n2618_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1769_3_lut_LC_21_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1769_3_lut_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1769_3_lut_LC_21_22_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1769_3_lut_LC_21_22_5  (
            .in0(_gnd_net_),
            .in1(N__19046),
            .in2(N__19052),
            .in3(N__22563),
            .lcout(\eeprom.n2717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_2_lut_LC_21_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_2_lut_LC_21_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_2_lut_LC_21_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_2_lut_LC_21_23_0  (
            .in0(_gnd_net_),
            .in1(N__24286),
            .in2(_gnd_net_),
            .in3(N__19049),
            .lcout(\eeprom.n2686 ),
            .ltout(),
            .carryin(bfn_21_23_0_),
            .carryout(\eeprom.n4043 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_3_lut_LC_21_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_3_lut_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_3_lut_LC_21_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_3_lut_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(N__28134),
            .in2(N__22273),
            .in3(N__19040),
            .lcout(\eeprom.n2685 ),
            .ltout(),
            .carryin(\eeprom.n4043 ),
            .carryout(\eeprom.n4044 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_4_lut_LC_21_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_4_lut_LC_21_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_4_lut_LC_21_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_4_lut_LC_21_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23816),
            .in3(N__19037),
            .lcout(\eeprom.n2684 ),
            .ltout(),
            .carryin(\eeprom.n4044 ),
            .carryout(\eeprom.n4045 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_5_lut_LC_21_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_5_lut_LC_21_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_5_lut_LC_21_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_5_lut_LC_21_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23759),
            .in3(N__19034),
            .lcout(\eeprom.n2683 ),
            .ltout(),
            .carryin(\eeprom.n4045 ),
            .carryout(\eeprom.n4046 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_6_lut_LC_21_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_6_lut_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_6_lut_LC_21_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_6_lut_LC_21_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23876),
            .in3(N__19289),
            .lcout(\eeprom.n2682 ),
            .ltout(),
            .carryin(\eeprom.n4046 ),
            .carryout(\eeprom.n4047 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_7_lut_LC_21_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_7_lut_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_7_lut_LC_21_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_7_lut_LC_21_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23789),
            .in3(N__19286),
            .lcout(\eeprom.n2681 ),
            .ltout(),
            .carryin(\eeprom.n4047 ),
            .carryout(\eeprom.n4048 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_8_lut_LC_21_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_8_lut_LC_21_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_8_lut_LC_21_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_8_lut_LC_21_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23846),
            .in3(N__19283),
            .lcout(\eeprom.n2680 ),
            .ltout(),
            .carryin(\eeprom.n4048 ),
            .carryout(\eeprom.n4049 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_9_lut_LC_21_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_9_lut_LC_21_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_9_lut_LC_21_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_9_lut_LC_21_23_7  (
            .in0(_gnd_net_),
            .in1(N__22358),
            .in2(N__28287),
            .in3(N__19280),
            .lcout(\eeprom.n2679 ),
            .ltout(),
            .carryin(\eeprom.n4049 ),
            .carryout(\eeprom.n4050 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_10_lut_LC_21_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_10_lut_LC_21_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_10_lut_LC_21_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_10_lut_LC_21_24_0  (
            .in0(_gnd_net_),
            .in1(N__22342),
            .in2(N__28288),
            .in3(N__19277),
            .lcout(\eeprom.n2678 ),
            .ltout(),
            .carryin(bfn_21_24_0_),
            .carryout(\eeprom.n4051 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_11_lut_LC_21_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_11_lut_LC_21_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_11_lut_LC_21_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_11_lut_LC_21_24_1  (
            .in0(_gnd_net_),
            .in1(N__28141),
            .in2(N__22309),
            .in3(N__19274),
            .lcout(\eeprom.n2677 ),
            .ltout(),
            .carryin(\eeprom.n4051 ),
            .carryout(\eeprom.n4052 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_12_lut_LC_21_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_12_lut_LC_21_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_12_lut_LC_21_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_12_lut_LC_21_24_2  (
            .in0(_gnd_net_),
            .in1(N__22139),
            .in2(N__28289),
            .in3(N__19271),
            .lcout(\eeprom.n2676 ),
            .ltout(),
            .carryin(\eeprom.n4052 ),
            .carryout(\eeprom.n4053 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_13_lut_LC_21_24_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_13_lut_LC_21_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_13_lut_LC_21_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_13_lut_LC_21_24_3  (
            .in0(_gnd_net_),
            .in1(N__22643),
            .in2(N__28290),
            .in3(N__19268),
            .lcout(\eeprom.n2675 ),
            .ltout(),
            .carryin(\eeprom.n4053 ),
            .carryout(\eeprom.n4054 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_14_lut_LC_21_24_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_14_lut_LC_21_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_14_lut_LC_21_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_14_lut_LC_21_24_4  (
            .in0(_gnd_net_),
            .in1(N__28149),
            .in2(N__22622),
            .in3(N__19265),
            .lcout(\eeprom.n2674 ),
            .ltout(),
            .carryin(\eeprom.n4054 ),
            .carryout(\eeprom.n4055 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_15_lut_LC_21_24_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1754_15_lut_LC_21_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_15_lut_LC_21_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1754_15_lut_LC_21_24_5  (
            .in0(_gnd_net_),
            .in1(N__22244),
            .in2(N__28291),
            .in3(N__19355),
            .lcout(\eeprom.n2673 ),
            .ltout(),
            .carryin(\eeprom.n4055 ),
            .carryout(\eeprom.n4056 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1754_16_lut_LC_21_24_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1754_16_lut_LC_21_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1754_16_lut_LC_21_24_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1754_16_lut_LC_21_24_6  (
            .in0(N__28145),
            .in1(N__24335),
            .in2(N__22590),
            .in3(N__19352),
            .lcout(\eeprom.n2704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1761_3_lut_LC_21_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1761_3_lut_LC_21_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1761_3_lut_LC_21_24_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1761_3_lut_LC_21_24_7  (
            .in0(_gnd_net_),
            .in1(N__19349),
            .in2(N__22310),
            .in3(N__22580),
            .lcout(\eeprom.n2709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1762_3_lut_LC_21_25_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1762_3_lut_LC_21_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1762_3_lut_LC_21_25_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1762_3_lut_LC_21_25_1  (
            .in0(_gnd_net_),
            .in1(N__19343),
            .in2(N__22592),
            .in3(N__22343),
            .lcout(\eeprom.n2710 ),
            .ltout(\eeprom.n2710_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_adj_84_LC_21_25_2 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_adj_84_LC_21_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_adj_84_LC_21_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_adj_84_LC_21_25_2  (
            .in0(N__21489),
            .in1(N__21177),
            .in2(N__19337),
            .in3(N__21223),
            .lcout(\eeprom.n17_adj_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1770_3_lut_LC_21_25_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1770_3_lut_LC_21_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1770_3_lut_LC_21_25_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1770_3_lut_LC_21_25_3  (
            .in0(N__19334),
            .in1(_gnd_net_),
            .in2(N__22591),
            .in3(N__24282),
            .lcout(\eeprom.n2718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1900_3_lut_LC_21_25_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1900_3_lut_LC_21_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1900_3_lut_LC_21_25_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1900_3_lut_LC_21_25_5  (
            .in0(_gnd_net_),
            .in1(N__19556),
            .in2(N__20786),
            .in3(N__19681),
            .lcout(\eeprom.n2912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_61_LC_21_26_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_61_LC_21_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_61_LC_21_26_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_61_LC_21_26_0  (
            .in0(N__20889),
            .in1(N__20802),
            .in2(N__20958),
            .in3(N__19484),
            .lcout(),
            .ltout(\eeprom.n5157_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_LC_21_26_1 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_LC_21_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_LC_21_26_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \eeprom.i5_4_lut_LC_21_26_1  (
            .in0(N__24256),
            .in1(N__20982),
            .in2(N__19301),
            .in3(N__20709),
            .lcout(\eeprom.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_60_LC_21_26_2 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_60_LC_21_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_60_LC_21_26_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_60_LC_21_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20847),
            .in3(N__20778),
            .lcout(\eeprom.n5153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1906_3_lut_LC_21_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1906_3_lut_LC_21_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1906_3_lut_LC_21_26_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1906_3_lut_LC_21_26_5  (
            .in0(N__24257),
            .in1(_gnd_net_),
            .in2(N__19421),
            .in3(N__19674),
            .lcout(\eeprom.n2918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1899_3_lut_LC_21_26_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1899_3_lut_LC_21_26_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1899_3_lut_LC_21_26_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1899_3_lut_LC_21_26_6  (
            .in0(N__20710),
            .in1(_gnd_net_),
            .in2(N__19682),
            .in3(N__19544),
            .lcout(\eeprom.n2911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_2_lut_LC_21_27_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_2_lut_LC_21_27_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_2_lut_LC_21_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_2_lut_LC_21_27_0  (
            .in0(_gnd_net_),
            .in1(N__24255),
            .in2(_gnd_net_),
            .in3(N__19412),
            .lcout(\eeprom.n2886 ),
            .ltout(),
            .carryin(bfn_21_27_0_),
            .carryout(\eeprom.n4072 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_3_lut_LC_21_27_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_3_lut_LC_21_27_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_3_lut_LC_21_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_3_lut_LC_21_27_1  (
            .in0(_gnd_net_),
            .in1(N__20986),
            .in2(N__28841),
            .in3(N__19403),
            .lcout(\eeprom.n2885 ),
            .ltout(),
            .carryin(\eeprom.n4072 ),
            .carryout(\eeprom.n4073 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_4_lut_LC_21_27_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_4_lut_LC_21_27_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_4_lut_LC_21_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_4_lut_LC_21_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20959),
            .in3(N__19391),
            .lcout(\eeprom.n2884 ),
            .ltout(),
            .carryin(\eeprom.n4073 ),
            .carryout(\eeprom.n4074 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_5_lut_LC_21_27_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_5_lut_LC_21_27_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_5_lut_LC_21_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_5_lut_LC_21_27_3  (
            .in0(_gnd_net_),
            .in1(N__20896),
            .in2(_gnd_net_),
            .in3(N__19382),
            .lcout(\eeprom.n2883 ),
            .ltout(),
            .carryin(\eeprom.n4074 ),
            .carryout(\eeprom.n4075 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_6_lut_LC_21_27_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_6_lut_LC_21_27_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_6_lut_LC_21_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_6_lut_LC_21_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20854),
            .in3(N__19367),
            .lcout(\eeprom.n2882 ),
            .ltout(),
            .carryin(\eeprom.n4075 ),
            .carryout(\eeprom.n4076 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_7_lut_LC_21_27_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_7_lut_LC_21_27_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_7_lut_LC_21_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_7_lut_LC_21_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20815),
            .in3(N__19358),
            .lcout(\eeprom.n2881 ),
            .ltout(),
            .carryin(\eeprom.n4076 ),
            .carryout(\eeprom.n4077 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_8_lut_LC_21_27_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_8_lut_LC_21_27_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_8_lut_LC_21_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_8_lut_LC_21_27_6  (
            .in0(_gnd_net_),
            .in1(N__20785),
            .in2(_gnd_net_),
            .in3(N__19547),
            .lcout(\eeprom.n2880 ),
            .ltout(),
            .carryin(\eeprom.n4077 ),
            .carryout(\eeprom.n4078 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_9_lut_LC_21_27_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_9_lut_LC_21_27_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_9_lut_LC_21_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_9_lut_LC_21_27_7  (
            .in0(_gnd_net_),
            .in1(N__28721),
            .in2(N__20717),
            .in3(N__19538),
            .lcout(\eeprom.n2879 ),
            .ltout(),
            .carryin(\eeprom.n4078 ),
            .carryout(\eeprom.n4079 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_10_lut_LC_21_28_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_10_lut_LC_21_28_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_10_lut_LC_21_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_10_lut_LC_21_28_0  (
            .in0(_gnd_net_),
            .in1(N__21360),
            .in2(N__28842),
            .in3(N__19529),
            .lcout(\eeprom.n2878 ),
            .ltout(),
            .carryin(bfn_21_28_0_),
            .carryout(\eeprom.n4080 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_11_lut_LC_21_28_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_11_lut_LC_21_28_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_11_lut_LC_21_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_11_lut_LC_21_28_1  (
            .in0(_gnd_net_),
            .in1(N__21304),
            .in2(N__28844),
            .in3(N__19517),
            .lcout(\eeprom.n2877 ),
            .ltout(),
            .carryin(\eeprom.n4080 ),
            .carryout(\eeprom.n4081 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_12_lut_LC_21_28_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_12_lut_LC_21_28_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_12_lut_LC_21_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_12_lut_LC_21_28_2  (
            .in0(_gnd_net_),
            .in1(N__28733),
            .in2(N__21274),
            .in3(N__19505),
            .lcout(\eeprom.n2876 ),
            .ltout(),
            .carryin(\eeprom.n4081 ),
            .carryout(\eeprom.n4082 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_13_lut_LC_21_28_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_13_lut_LC_21_28_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_13_lut_LC_21_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_13_lut_LC_21_28_3  (
            .in0(_gnd_net_),
            .in1(N__21211),
            .in2(N__28845),
            .in3(N__19502),
            .lcout(\eeprom.n2875 ),
            .ltout(),
            .carryin(\eeprom.n4082 ),
            .carryout(\eeprom.n4083 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_14_lut_LC_21_28_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_14_lut_LC_21_28_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_14_lut_LC_21_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_14_lut_LC_21_28_4  (
            .in0(_gnd_net_),
            .in1(N__28737),
            .in2(N__21164),
            .in3(N__19490),
            .lcout(\eeprom.n2874 ),
            .ltout(),
            .carryin(\eeprom.n4083 ),
            .carryout(\eeprom.n4084 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_15_lut_LC_21_28_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_15_lut_LC_21_28_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_15_lut_LC_21_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_15_lut_LC_21_28_5  (
            .in0(_gnd_net_),
            .in1(N__28725),
            .in2(N__21110),
            .in3(N__19487),
            .lcout(\eeprom.n2873 ),
            .ltout(),
            .carryin(\eeprom.n4084 ),
            .carryout(\eeprom.n4085 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_16_lut_LC_21_28_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_16_lut_LC_21_28_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_16_lut_LC_21_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_16_lut_LC_21_28_6  (
            .in0(_gnd_net_),
            .in1(N__21072),
            .in2(N__28843),
            .in3(N__19811),
            .lcout(\eeprom.n2872 ),
            .ltout(),
            .carryin(\eeprom.n4085 ),
            .carryout(\eeprom.n4086 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_17_lut_LC_21_28_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1888_17_lut_LC_21_28_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_17_lut_LC_21_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1888_17_lut_LC_21_28_7  (
            .in0(_gnd_net_),
            .in1(N__28729),
            .in2(N__21029),
            .in3(N__19808),
            .lcout(\eeprom.n2871 ),
            .ltout(),
            .carryin(\eeprom.n4086 ),
            .carryout(\eeprom.n4087 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1888_18_lut_LC_21_29_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1888_18_lut_LC_21_29_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1888_18_lut_LC_21_29_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1888_18_lut_LC_21_29_0  (
            .in0(N__28153),
            .in1(N__21400),
            .in2(N__19680),
            .in3(N__19805),
            .lcout(\eeprom.n2902 ),
            .ltout(\eeprom.n2902_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_adj_62_LC_21_29_1 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_adj_62_LC_21_29_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_adj_62_LC_21_29_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_adj_62_LC_21_29_1  (
            .in0(N__19770),
            .in1(N__19740),
            .in2(N__19793),
            .in3(N__19707),
            .lcout(\eeprom.n19_adj_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1892_3_lut_LC_21_29_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1892_3_lut_LC_21_29_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1892_3_lut_LC_21_29_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1892_3_lut_LC_21_29_2  (
            .in0(N__21073),
            .in1(_gnd_net_),
            .in2(N__19678),
            .in3(N__19781),
            .lcout(\eeprom.n2904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1893_3_lut_LC_21_29_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1893_3_lut_LC_21_29_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1893_3_lut_LC_21_29_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1893_3_lut_LC_21_29_4  (
            .in0(N__21102),
            .in1(_gnd_net_),
            .in2(N__19679),
            .in3(N__19754),
            .lcout(\eeprom.n2905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1891_3_lut_LC_21_29_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1891_3_lut_LC_21_29_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1891_3_lut_LC_21_29_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i1891_3_lut_LC_21_29_5  (
            .in0(N__19724),
            .in1(_gnd_net_),
            .in2(N__21028),
            .in3(N__19656),
            .lcout(\eeprom.n2903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1895_3_lut_LC_21_29_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1895_3_lut_LC_21_29_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1895_3_lut_LC_21_29_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1895_3_lut_LC_21_29_7  (
            .in0(_gnd_net_),
            .in1(N__21212),
            .in2(N__19691),
            .in3(N__19666),
            .lcout(\eeprom.n2907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_2_lut_LC_22_17_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_2_lut_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_2_lut_LC_22_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_2_lut_LC_22_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21998),
            .in3(N__19559),
            .lcout(\eeprom.n2286 ),
            .ltout(),
            .carryin(bfn_22_17_0_),
            .carryout(\eeprom.n3997 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_3_lut_LC_22_17_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_3_lut_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_3_lut_LC_22_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_3_lut_LC_22_17_1  (
            .in0(_gnd_net_),
            .in1(N__28190),
            .in2(N__19954),
            .in3(N__19895),
            .lcout(\eeprom.n2285 ),
            .ltout(),
            .carryin(\eeprom.n3997 ),
            .carryout(\eeprom.n3998 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_4_lut_LC_22_17_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_4_lut_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_4_lut_LC_22_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_4_lut_LC_22_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20231),
            .in3(N__19892),
            .lcout(\eeprom.n2284 ),
            .ltout(),
            .carryin(\eeprom.n3998 ),
            .carryout(\eeprom.n3999 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_5_lut_LC_22_17_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_5_lut_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_5_lut_LC_22_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_5_lut_LC_22_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19990),
            .in3(N__19880),
            .lcout(\eeprom.n2283 ),
            .ltout(),
            .carryin(\eeprom.n3999 ),
            .carryout(\eeprom.n4000 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_6_lut_LC_22_17_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_6_lut_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_6_lut_LC_22_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_6_lut_LC_22_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19877),
            .in3(N__19862),
            .lcout(\eeprom.n2282 ),
            .ltout(),
            .carryin(\eeprom.n4000 ),
            .carryout(\eeprom.n4001 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_7_lut_LC_22_17_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_7_lut_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_7_lut_LC_22_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_7_lut_LC_22_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19859),
            .in3(N__19829),
            .lcout(\eeprom.n2281 ),
            .ltout(),
            .carryin(\eeprom.n4001 ),
            .carryout(\eeprom.n4002 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_8_lut_LC_22_17_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_8_lut_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_8_lut_LC_22_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_8_lut_LC_22_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20189),
            .in3(N__19826),
            .lcout(\eeprom.n2280 ),
            .ltout(),
            .carryin(\eeprom.n4002 ),
            .carryout(\eeprom.n4003 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_9_lut_LC_22_17_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_9_lut_LC_22_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_9_lut_LC_22_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_9_lut_LC_22_17_7  (
            .in0(_gnd_net_),
            .in1(N__21640),
            .in2(N__28352),
            .in3(N__19823),
            .lcout(\eeprom.n2279 ),
            .ltout(),
            .carryin(\eeprom.n4003 ),
            .carryout(\eeprom.n4004 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_10_lut_LC_22_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_10_lut_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_10_lut_LC_22_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_10_lut_LC_22_18_0  (
            .in0(_gnd_net_),
            .in1(N__28264),
            .in2(N__19925),
            .in3(N__19814),
            .lcout(\eeprom.n2278 ),
            .ltout(),
            .carryin(bfn_22_18_0_),
            .carryout(\eeprom.n4005 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_11_lut_LC_22_18_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1486_11_lut_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_11_lut_LC_22_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1486_11_lut_LC_22_18_1  (
            .in0(_gnd_net_),
            .in1(N__21955),
            .in2(N__28411),
            .in3(N__19997),
            .lcout(\eeprom.n2277 ),
            .ltout(),
            .carryin(\eeprom.n4005 ),
            .carryout(\eeprom.n4006 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1486_12_lut_LC_22_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1486_12_lut_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1486_12_lut_LC_22_18_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \eeprom.rem_4_add_1486_12_lut_LC_22_18_2  (
            .in0(N__21737),
            .in1(N__28268),
            .in2(N__23090),
            .in3(N__19994),
            .lcout(\eeprom.n2308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1425_3_lut_LC_22_18_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1425_3_lut_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1425_3_lut_LC_22_18_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1425_3_lut_LC_22_18_3  (
            .in0(_gnd_net_),
            .in1(N__22777),
            .in2(N__23154),
            .in3(N__22757),
            .lcout(\eeprom.n2213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1428_3_lut_LC_22_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1428_3_lut_LC_22_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1428_3_lut_LC_22_18_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1428_3_lut_LC_22_18_4  (
            .in0(_gnd_net_),
            .in1(N__22882),
            .in2(N__22862),
            .in3(N__23140),
            .lcout(\eeprom.n2216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_adj_51_LC_22_18_5 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_adj_51_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_adj_51_LC_22_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i3_4_lut_adj_51_LC_22_18_5  (
            .in0(N__23167),
            .in1(N__23026),
            .in2(N__22726),
            .in3(N__21647),
            .lcout(\eeprom.n2143 ),
            .ltout(\eeprom.n2143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1429_rep_44_3_lut_LC_22_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1429_rep_44_3_lut_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1429_rep_44_3_lut_LC_22_18_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1429_rep_44_3_lut_LC_22_18_6  (
            .in0(_gnd_net_),
            .in1(N__22912),
            .in2(N__19967),
            .in3(N__22898),
            .lcout(\eeprom.n2217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1498_3_lut_LC_22_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1498_3_lut_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1498_3_lut_LC_22_19_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1498_3_lut_LC_22_19_0  (
            .in0(_gnd_net_),
            .in1(N__21993),
            .in2(N__21739),
            .in3(N__19964),
            .lcout(\eeprom.n2318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_54_LC_22_19_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_54_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_54_LC_22_19_1 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_54_LC_22_19_1  (
            .in0(N__20184),
            .in1(N__19950),
            .in2(N__21997),
            .in3(N__19931),
            .lcout(),
            .ltout(\eeprom.n4797_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4_4_lut_adj_55_LC_22_19_2 .C_ON=1'b0;
    defparam \eeprom.i4_4_lut_adj_55_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4_4_lut_adj_55_LC_22_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i4_4_lut_adj_55_LC_22_19_2  (
            .in0(N__21636),
            .in1(N__19921),
            .in2(N__19910),
            .in3(N__21938),
            .lcout(\eeprom.n2242 ),
            .ltout(\eeprom.n2242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1427_rep_42_3_lut_LC_22_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1427_rep_42_3_lut_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1427_rep_42_3_lut_LC_22_19_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1427_rep_42_3_lut_LC_22_19_3  (
            .in0(_gnd_net_),
            .in1(N__20171),
            .in2(N__20246),
            .in3(N__20243),
            .lcout(),
            .ltout(\eeprom.n5400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4677_3_lut_LC_22_19_4 .C_ON=1'b0;
    defparam \eeprom.i4677_3_lut_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4677_3_lut_LC_22_19_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.i4677_3_lut_LC_22_19_4  (
            .in0(_gnd_net_),
            .in1(N__22977),
            .in2(N__20234),
            .in3(N__21680),
            .lcout(\eeprom.n2314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4679_3_lut_LC_22_19_5 .C_ON=1'b0;
    defparam \eeprom.i4679_3_lut_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4679_3_lut_LC_22_19_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.i4679_3_lut_LC_22_19_5  (
            .in0(_gnd_net_),
            .in1(N__20230),
            .in2(N__20210),
            .in3(N__21727),
            .lcout(\eeprom.n2316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1492_3_lut_LC_22_19_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1492_3_lut_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1492_3_lut_LC_22_19_6 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i1492_3_lut_LC_22_19_6  (
            .in0(N__20198),
            .in1(N__20185),
            .in2(N__21740),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1360_rep_47_3_lut_LC_22_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1360_rep_47_3_lut_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1360_rep_47_3_lut_LC_22_19_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1360_rep_47_3_lut_LC_22_19_7  (
            .in0(_gnd_net_),
            .in1(N__22820),
            .in2(N__23155),
            .in3(N__21542),
            .lcout(\eeprom.n5405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_57_LC_22_20_0 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_57_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_57_LC_22_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_57_LC_22_20_0  (
            .in0(N__20163),
            .in1(N__20145),
            .in2(N__20129),
            .in3(N__20024),
            .lcout(),
            .ltout(\eeprom.n5085_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_58_LC_22_20_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_58_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_58_LC_22_20_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \eeprom.i1_4_lut_adj_58_LC_22_20_1  (
            .in0(N__24600),
            .in1(N__20106),
            .in2(N__20090),
            .in3(N__20085),
            .lcout(\eeprom.n7_adj_323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_56_LC_22_20_2 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_56_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_56_LC_22_20_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_56_LC_22_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20063),
            .in3(N__20040),
            .lcout(\eeprom.n5081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1489_3_lut_LC_22_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1489_3_lut_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1489_3_lut_LC_22_20_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1489_3_lut_LC_22_20_3  (
            .in0(_gnd_net_),
            .in1(N__20018),
            .in2(N__21959),
            .in3(N__21736),
            .lcout(\eeprom.n2309 ),
            .ltout(\eeprom.n2309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2_2_lut_LC_22_20_4 .C_ON=1'b0;
    defparam \eeprom.i2_2_lut_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_2_lut_LC_22_20_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i2_2_lut_LC_22_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20432),
            .in3(N__20271),
            .lcout(),
            .ltout(\eeprom.n8_adj_322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_59_LC_22_20_5 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_59_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_59_LC_22_20_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_adj_59_LC_22_20_5  (
            .in0(N__20421),
            .in1(N__20392),
            .in2(N__20381),
            .in3(N__20378),
            .lcout(\eeprom.n2341 ),
            .ltout(\eeprom.n2341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4746_1_lut_LC_22_20_6 .C_ON=1'b0;
    defparam \eeprom.i4746_1_lut_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4746_1_lut_LC_22_20_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4746_1_lut_LC_22_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20327),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1491_3_lut_LC_22_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1491_3_lut_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1491_3_lut_LC_22_20_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1491_3_lut_LC_22_20_7  (
            .in0(_gnd_net_),
            .in1(N__20282),
            .in2(N__21641),
            .in3(N__21735),
            .lcout(\eeprom.n2311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_26_LC_22_21_0 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_26_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_26_LC_22_21_0 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_26_LC_22_21_0  (
            .in0(_gnd_net_),
            .in1(N__20454),
            .in2(N__21921),
            .in3(N__20607),
            .lcout(),
            .ltout(\eeprom.n5073_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_27_LC_22_21_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_27_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_27_LC_22_21_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_27_LC_22_21_1  (
            .in0(N__21876),
            .in1(N__22441),
            .in2(N__20255),
            .in3(N__20483),
            .lcout(),
            .ltout(\eeprom.n4782_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_28_LC_22_21_2 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_28_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_28_LC_22_21_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_adj_28_LC_22_21_2  (
            .in0(N__23526),
            .in1(N__20535),
            .in2(N__20252),
            .in3(N__21837),
            .lcout(),
            .ltout(\eeprom.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_4_lut_LC_22_21_3 .C_ON=1'b0;
    defparam \eeprom.i6_4_lut_LC_22_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_4_lut_LC_22_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i6_4_lut_LC_22_21_3  (
            .in0(N__20577),
            .in1(N__21813),
            .in2(N__20249),
            .in3(N__20500),
            .lcout(\eeprom.n2440 ),
            .ltout(\eeprom.n2440_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1629_3_lut_LC_22_21_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1629_3_lut_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1629_3_lut_LC_22_21_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1629_3_lut_LC_22_21_4  (
            .in0(_gnd_net_),
            .in1(N__20455),
            .in2(N__20486),
            .in3(N__20441),
            .lcout(\eeprom.n2513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_25_LC_22_21_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_25_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_25_LC_22_21_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_25_LC_22_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21765),
            .in3(N__22095),
            .lcout(\eeprom.n5071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1628_3_lut_LC_22_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1628_3_lut_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1628_3_lut_LC_22_21_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1628_3_lut_LC_22_21_6  (
            .in0(_gnd_net_),
            .in1(N__20608),
            .in2(N__20594),
            .in3(N__23479),
            .lcout(\eeprom.n2512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1624_3_lut_LC_22_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1624_3_lut_LC_22_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1624_3_lut_LC_22_21_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \eeprom.rem_4_i1624_3_lut_LC_22_21_7  (
            .in0(N__20536),
            .in1(N__20522),
            .in2(N__23493),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_2_lut_LC_22_22_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_2_lut_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_2_lut_LC_22_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_2_lut_LC_22_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22440),
            .in3(N__20477),
            .lcout(\eeprom.n2486 ),
            .ltout(),
            .carryin(bfn_22_22_0_),
            .carryout(\eeprom.n4018 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_3_lut_LC_22_22_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_3_lut_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_3_lut_LC_22_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_3_lut_LC_22_22_1  (
            .in0(_gnd_net_),
            .in1(N__21880),
            .in2(N__28549),
            .in3(N__20474),
            .lcout(\eeprom.n2485 ),
            .ltout(),
            .carryin(\eeprom.n4018 ),
            .carryout(\eeprom.n4019 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_4_lut_LC_22_22_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_4_lut_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_4_lut_LC_22_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_4_lut_LC_22_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21772),
            .in3(N__20471),
            .lcout(\eeprom.n2484 ),
            .ltout(),
            .carryin(\eeprom.n4019 ),
            .carryout(\eeprom.n4020 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_5_lut_LC_22_22_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_5_lut_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_5_lut_LC_22_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_5_lut_LC_22_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21925),
            .in3(N__20468),
            .lcout(\eeprom.n2483 ),
            .ltout(),
            .carryin(\eeprom.n4020 ),
            .carryout(\eeprom.n4021 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_6_lut_LC_22_22_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_6_lut_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_6_lut_LC_22_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_6_lut_LC_22_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22108),
            .in3(N__20465),
            .lcout(\eeprom.n2482 ),
            .ltout(),
            .carryin(\eeprom.n4021 ),
            .carryout(\eeprom.n4022 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_7_lut_LC_22_22_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_7_lut_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_7_lut_LC_22_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_7_lut_LC_22_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20462),
            .in3(N__20435),
            .lcout(\eeprom.n2481 ),
            .ltout(),
            .carryin(\eeprom.n4022 ),
            .carryout(\eeprom.n4023 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_8_lut_LC_22_22_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_8_lut_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_8_lut_LC_22_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_8_lut_LC_22_22_6  (
            .in0(_gnd_net_),
            .in1(N__20612),
            .in2(_gnd_net_),
            .in3(N__20585),
            .lcout(\eeprom.n2480 ),
            .ltout(),
            .carryin(\eeprom.n4023 ),
            .carryout(\eeprom.n4024 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_9_lut_LC_22_22_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_9_lut_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_9_lut_LC_22_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_9_lut_LC_22_22_7  (
            .in0(_gnd_net_),
            .in1(N__20581),
            .in2(N__28550),
            .in3(N__20549),
            .lcout(\eeprom.n2479 ),
            .ltout(),
            .carryin(\eeprom.n4024 ),
            .carryout(\eeprom.n4025 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_10_lut_LC_22_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_10_lut_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_10_lut_LC_22_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_10_lut_LC_22_23_0  (
            .in0(_gnd_net_),
            .in1(N__28400),
            .in2(N__23539),
            .in3(N__20546),
            .lcout(\eeprom.n2478 ),
            .ltout(),
            .carryin(bfn_22_23_0_),
            .carryout(\eeprom.n4026 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_11_lut_LC_22_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_11_lut_LC_22_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_11_lut_LC_22_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_11_lut_LC_22_23_1  (
            .in0(_gnd_net_),
            .in1(N__21844),
            .in2(N__28551),
            .in3(N__20543),
            .lcout(\eeprom.n2477 ),
            .ltout(),
            .carryin(\eeprom.n4026 ),
            .carryout(\eeprom.n4027 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_12_lut_LC_22_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_12_lut_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_12_lut_LC_22_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_12_lut_LC_22_23_2  (
            .in0(_gnd_net_),
            .in1(N__20540),
            .in2(N__28553),
            .in3(N__20513),
            .lcout(\eeprom.n2476 ),
            .ltout(),
            .carryin(\eeprom.n4027 ),
            .carryout(\eeprom.n4028 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_13_lut_LC_22_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1620_13_lut_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_13_lut_LC_22_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1620_13_lut_LC_22_23_3  (
            .in0(_gnd_net_),
            .in1(N__21820),
            .in2(N__28552),
            .in3(N__20510),
            .lcout(\eeprom.n2475 ),
            .ltout(),
            .carryin(\eeprom.n4028 ),
            .carryout(\eeprom.n4029 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1620_14_lut_LC_22_23_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1620_14_lut_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1620_14_lut_LC_22_23_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \eeprom.rem_4_add_1620_14_lut_LC_22_23_4  (
            .in0(N__23495),
            .in1(N__28407),
            .in2(N__20507),
            .in3(N__20489),
            .lcout(\eeprom.n2506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i8_4_lut_adj_75_LC_22_23_5 .C_ON=1'b0;
    defparam \eeprom.i8_4_lut_adj_75_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i8_4_lut_adj_75_LC_22_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i8_4_lut_adj_75_LC_22_23_5  (
            .in0(N__22638),
            .in1(N__22615),
            .in2(N__22253),
            .in3(N__22280),
            .lcout(\eeprom.n2638 ),
            .ltout(\eeprom.n2638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1768_3_lut_LC_22_23_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1768_3_lut_LC_22_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1768_3_lut_LC_22_23_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1768_3_lut_LC_22_23_6  (
            .in0(_gnd_net_),
            .in1(N__23809),
            .in2(N__20675),
            .in3(N__20672),
            .lcout(\eeprom.n2716 ),
            .ltout(\eeprom.n2716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_81_LC_22_23_7 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_81_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_81_LC_22_23_7 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \eeprom.i1_3_lut_adj_81_LC_22_23_7  (
            .in0(N__22155),
            .in1(N__20916),
            .in2(N__20666),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1764_3_lut_LC_22_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1764_3_lut_LC_22_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1764_3_lut_LC_22_24_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1764_3_lut_LC_22_24_0  (
            .in0(_gnd_net_),
            .in1(N__23842),
            .in2(N__20663),
            .in3(N__22575),
            .lcout(\eeprom.n2712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1763_3_lut_LC_22_24_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1763_3_lut_LC_22_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1763_3_lut_LC_22_24_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \eeprom.rem_4_i1763_3_lut_LC_22_24_1  (
            .in0(N__20654),
            .in1(N__22357),
            .in2(N__22588),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1760_3_lut_LC_22_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1760_3_lut_LC_22_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1760_3_lut_LC_22_24_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \eeprom.rem_4_i1760_3_lut_LC_22_24_2  (
            .in0(N__22138),
            .in1(_gnd_net_),
            .in2(N__20648),
            .in3(N__22568),
            .lcout(\eeprom.n2708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1759_3_lut_LC_22_24_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1759_3_lut_LC_22_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1759_3_lut_LC_22_24_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1759_3_lut_LC_22_24_3  (
            .in0(_gnd_net_),
            .in1(N__20639),
            .in2(N__22589),
            .in3(N__22642),
            .lcout(\eeprom.n2707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1757_3_lut_LC_22_24_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1757_3_lut_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1757_3_lut_LC_22_24_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1757_3_lut_LC_22_24_4  (
            .in0(_gnd_net_),
            .in1(N__22243),
            .in2(N__20633),
            .in3(N__22576),
            .lcout(\eeprom.n2705 ),
            .ltout(\eeprom.n2705_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_4_lut_adj_83_LC_22_24_5 .C_ON=1'b0;
    defparam \eeprom.i6_4_lut_adj_83_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_4_lut_adj_83_LC_22_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i6_4_lut_adj_83_LC_22_24_5  (
            .in0(N__21324),
            .in1(N__22500),
            .in2(N__20624),
            .in3(N__22175),
            .lcout(),
            .ltout(\eeprom.n16_adj_338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i9_4_lut_adj_86_LC_22_24_6 .C_ON=1'b0;
    defparam \eeprom.i9_4_lut_adj_86_LC_22_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i9_4_lut_adj_86_LC_22_24_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i9_4_lut_adj_86_LC_22_24_6  (
            .in0(N__21126),
            .in1(N__20621),
            .in2(N__20615),
            .in3(N__20691),
            .lcout(\eeprom.n2737 ),
            .ltout(\eeprom.n2737_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4745_1_lut_LC_22_24_7 .C_ON=1'b0;
    defparam \eeprom.i4745_1_lut_LC_22_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4745_1_lut_LC_22_24_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.i4745_1_lut_LC_22_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20993),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_2_lut_LC_22_25_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_2_lut_LC_22_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_2_lut_LC_22_25_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1821_2_lut_LC_22_25_0  (
            .in0(N__22485),
            .in1(N__22487),
            .in2(N__20754),
            .in3(N__20963),
            .lcout(\eeprom.n2818 ),
            .ltout(),
            .carryin(bfn_22_25_0_),
            .carryout(\eeprom.n4057 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_3_lut_LC_22_25_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_3_lut_LC_22_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_3_lut_LC_22_25_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_3_lut_LC_22_25_1  (
            .in0(N__22209),
            .in1(N__22213),
            .in2(N__21443),
            .in3(N__20930),
            .lcout(\eeprom.n2817 ),
            .ltout(),
            .carryin(\eeprom.n4057 ),
            .carryout(\eeprom.n4058 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_4_lut_LC_22_25_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_4_lut_LC_22_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_4_lut_LC_22_25_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1821_4_lut_LC_22_25_2  (
            .in0(N__20926),
            .in1(N__20927),
            .in2(N__20755),
            .in3(N__20876),
            .lcout(\eeprom.n2816 ),
            .ltout(),
            .carryin(\eeprom.n4058 ),
            .carryout(\eeprom.n4059 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_5_lut_LC_22_25_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_5_lut_LC_22_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_5_lut_LC_22_25_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1821_5_lut_LC_22_25_3  (
            .in0(N__20873),
            .in1(N__20872),
            .in2(N__20758),
            .in3(N__20822),
            .lcout(\eeprom.n2815 ),
            .ltout(),
            .carryin(\eeprom.n4059 ),
            .carryout(\eeprom.n4060 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_6_lut_LC_22_25_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_6_lut_LC_22_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_6_lut_LC_22_25_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1821_6_lut_LC_22_25_4  (
            .in0(N__22025),
            .in1(N__22024),
            .in2(N__20756),
            .in3(N__20789),
            .lcout(\eeprom.n2814 ),
            .ltout(),
            .carryin(\eeprom.n4060 ),
            .carryout(\eeprom.n4061 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_7_lut_LC_22_25_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_7_lut_LC_22_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_7_lut_LC_22_25_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1821_7_lut_LC_22_25_5  (
            .in0(N__22157),
            .in1(N__22156),
            .in2(N__20759),
            .in3(N__20762),
            .lcout(\eeprom.n2813 ),
            .ltout(),
            .carryin(\eeprom.n4061 ),
            .carryout(\eeprom.n4062 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_8_lut_LC_22_25_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_8_lut_LC_22_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_8_lut_LC_22_25_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \eeprom.rem_4_add_1821_8_lut_LC_22_25_6  (
            .in0(N__22046),
            .in1(N__22042),
            .in2(N__20757),
            .in3(N__20696),
            .lcout(\eeprom.n2812 ),
            .ltout(),
            .carryin(\eeprom.n4062 ),
            .carryout(\eeprom.n4063 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_9_lut_LC_22_25_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_9_lut_LC_22_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_9_lut_LC_22_25_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_9_lut_LC_22_25_7  (
            .in0(N__20693),
            .in1(N__20692),
            .in2(N__21444),
            .in3(N__21335),
            .lcout(\eeprom.n2811 ),
            .ltout(),
            .carryin(\eeprom.n4063 ),
            .carryout(\eeprom.n4064 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_10_lut_LC_22_26_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_10_lut_LC_22_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_10_lut_LC_22_26_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_10_lut_LC_22_26_0  (
            .in0(N__21332),
            .in1(N__21331),
            .in2(N__21469),
            .in3(N__21290),
            .lcout(\eeprom.n2810 ),
            .ltout(),
            .carryin(bfn_22_26_0_),
            .carryout(\eeprom.n4065 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_11_lut_LC_22_26_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_11_lut_LC_22_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_11_lut_LC_22_26_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_11_lut_LC_22_26_1  (
            .in0(N__21287),
            .in1(N__21286),
            .in2(N__21473),
            .in3(N__21239),
            .lcout(\eeprom.n2809 ),
            .ltout(),
            .carryin(\eeprom.n4065 ),
            .carryout(\eeprom.n4066 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_12_lut_LC_22_26_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_12_lut_LC_22_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_12_lut_LC_22_26_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_12_lut_LC_22_26_2  (
            .in0(N__21236),
            .in1(N__21235),
            .in2(N__21470),
            .in3(N__21188),
            .lcout(\eeprom.n2808 ),
            .ltout(),
            .carryin(\eeprom.n4066 ),
            .carryout(\eeprom.n4067 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_13_lut_LC_22_26_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_13_lut_LC_22_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_13_lut_LC_22_26_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_13_lut_LC_22_26_3  (
            .in0(N__21185),
            .in1(N__21184),
            .in2(N__21474),
            .in3(N__21137),
            .lcout(\eeprom.n2807 ),
            .ltout(),
            .carryin(\eeprom.n4067 ),
            .carryout(\eeprom.n4068 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_14_lut_LC_22_26_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_14_lut_LC_22_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_14_lut_LC_22_26_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_14_lut_LC_22_26_4  (
            .in0(N__21134),
            .in1(N__21133),
            .in2(N__21471),
            .in3(N__21077),
            .lcout(\eeprom.n2806 ),
            .ltout(),
            .carryin(\eeprom.n4068 ),
            .carryout(\eeprom.n4069 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_15_lut_LC_22_26_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_15_lut_LC_22_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_15_lut_LC_22_26_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_15_lut_LC_22_26_5  (
            .in0(N__22510),
            .in1(N__22511),
            .in2(N__21475),
            .in3(N__21047),
            .lcout(\eeprom.n2805 ),
            .ltout(),
            .carryin(\eeprom.n4069 ),
            .carryout(\eeprom.n4070 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_16_lut_LC_22_26_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1821_16_lut_LC_22_26_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_16_lut_LC_22_26_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_16_lut_LC_22_26_6  (
            .in0(N__21044),
            .in1(N__21043),
            .in2(N__21472),
            .in3(N__20996),
            .lcout(\eeprom.n2804 ),
            .ltout(),
            .carryin(\eeprom.n4070 ),
            .carryout(\eeprom.n4071 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1821_17_lut_LC_22_26_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1821_17_lut_LC_22_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1821_17_lut_LC_22_26_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \eeprom.rem_4_add_1821_17_lut_LC_22_26_7  (
            .in0(N__21496),
            .in1(N__21497),
            .in2(N__21476),
            .in3(N__21404),
            .lcout(\eeprom.n2803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_105_LC_23_17_0 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_105_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_105_LC_23_17_0 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_105_LC_23_17_0  (
            .in0(_gnd_net_),
            .in1(N__23049),
            .in2(N__22978),
            .in3(N__23392),
            .lcout(),
            .ltout(\eeprom.n5005_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_106_LC_23_17_1 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_106_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_106_LC_23_17_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \eeprom.i1_4_lut_adj_106_LC_23_17_1  (
            .in0(N__22941),
            .in1(N__21617),
            .in2(N__21380),
            .in3(N__22998),
            .lcout(),
            .ltout(\eeprom.n5009_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_107_LC_23_17_2 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_107_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_107_LC_23_17_2 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \eeprom.i1_4_lut_adj_107_LC_23_17_2  (
            .in0(N__23231),
            .in1(N__23257),
            .in2(N__21377),
            .in3(N__23561),
            .lcout(\eeprom.n2044 ),
            .ltout(\eeprom.n2044_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1358_3_lut_LC_23_17_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1358_3_lut_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1358_3_lut_LC_23_17_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1358_3_lut_LC_23_17_3  (
            .in0(N__23050),
            .in1(_gnd_net_),
            .in2(N__21374),
            .in3(N__21524),
            .lcout(\eeprom.n2114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1360_3_lut_LC_23_17_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1360_3_lut_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1360_3_lut_LC_23_17_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1360_3_lut_LC_23_17_4  (
            .in0(_gnd_net_),
            .in1(N__21541),
            .in2(N__22979),
            .in3(N__23341),
            .lcout(\eeprom.n2116 ),
            .ltout(\eeprom.n2116_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_49_LC_23_17_5 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_49_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_49_LC_23_17_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_3_lut_adj_49_LC_23_17_5  (
            .in0(_gnd_net_),
            .in1(N__22773),
            .in2(N__21371),
            .in3(N__22878),
            .lcout(\eeprom.n5061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1361_3_lut_LC_23_17_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1361_3_lut_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1361_3_lut_LC_23_17_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1361_3_lut_LC_23_17_6  (
            .in0(_gnd_net_),
            .in1(N__21551),
            .in2(N__23003),
            .in3(N__23340),
            .lcout(\eeprom.n2117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1356_3_lut_LC_23_17_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1356_3_lut_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1356_3_lut_LC_23_17_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1356_3_lut_LC_23_17_7  (
            .in0(N__21512),
            .in1(_gnd_net_),
            .in2(N__23358),
            .in3(N__23258),
            .lcout(\eeprom.n2112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_2_lut_LC_23_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_2_lut_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_2_lut_LC_23_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_2_lut_LC_23_18_0  (
            .in0(_gnd_net_),
            .in1(N__21616),
            .in2(_gnd_net_),
            .in3(N__21368),
            .lcout(\eeprom.n2086 ),
            .ltout(),
            .carryin(bfn_23_18_0_),
            .carryout(\eeprom.n3980 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_3_lut_LC_23_18_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_3_lut_LC_23_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_3_lut_LC_23_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_3_lut_LC_23_18_1  (
            .in0(_gnd_net_),
            .in1(N__28242),
            .in2(N__23002),
            .in3(N__21545),
            .lcout(\eeprom.n2085 ),
            .ltout(),
            .carryin(\eeprom.n3980 ),
            .carryout(\eeprom.n3981 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_4_lut_LC_23_18_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_4_lut_LC_23_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_4_lut_LC_23_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_4_lut_LC_23_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22976),
            .in3(N__21530),
            .lcout(\eeprom.n2084 ),
            .ltout(),
            .carryin(\eeprom.n3981 ),
            .carryout(\eeprom.n3982 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_5_lut_LC_23_18_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_5_lut_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_5_lut_LC_23_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_5_lut_LC_23_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23393),
            .in3(N__21527),
            .lcout(\eeprom.n2083 ),
            .ltout(),
            .carryin(\eeprom.n3982 ),
            .carryout(\eeprom.n3983 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_6_lut_LC_23_18_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_6_lut_LC_23_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_6_lut_LC_23_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_6_lut_LC_23_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23054),
            .in3(N__21518),
            .lcout(\eeprom.n2082 ),
            .ltout(),
            .carryin(\eeprom.n3983 ),
            .carryout(\eeprom.n3984 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_7_lut_LC_23_18_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_7_lut_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_7_lut_LC_23_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_7_lut_LC_23_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22942),
            .in3(N__21515),
            .lcout(\eeprom.n2081 ),
            .ltout(),
            .carryin(\eeprom.n3984 ),
            .carryout(\eeprom.n3985 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_8_lut_LC_23_18_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_8_lut_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_8_lut_LC_23_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_8_lut_LC_23_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23256),
            .in3(N__21506),
            .lcout(\eeprom.n2080 ),
            .ltout(),
            .carryin(\eeprom.n3985 ),
            .carryout(\eeprom.n3986 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_9_lut_LC_23_18_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1352_9_lut_LC_23_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_9_lut_LC_23_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1352_9_lut_LC_23_18_7  (
            .in0(_gnd_net_),
            .in1(N__23229),
            .in2(N__28393),
            .in3(N__21503),
            .lcout(\eeprom.n2079 ),
            .ltout(),
            .carryin(\eeprom.n3986 ),
            .carryout(\eeprom.n3987 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1352_10_lut_LC_23_19_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1352_10_lut_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1352_10_lut_LC_23_19_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \eeprom.rem_4_add_1352_10_lut_LC_23_19_0  (
            .in0(N__28243),
            .in1(N__23363),
            .in2(N__23560),
            .in3(N__21500),
            .lcout(\eeprom.n2110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4671_3_lut_LC_23_19_1 .C_ON=1'b0;
    defparam \eeprom.i4671_3_lut_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4671_3_lut_LC_23_19_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \eeprom.i4671_3_lut_LC_23_19_1  (
            .in0(N__23364),
            .in1(N__23146),
            .in2(_gnd_net_),
            .in3(N__21721),
            .lcout(\eeprom.n5501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1422_3_lut_LC_23_19_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1422_3_lut_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1422_3_lut_LC_23_19_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \eeprom.rem_4_i1422_3_lut_LC_23_19_2  (
            .in0(N__23144),
            .in1(N__23025),
            .in2(N__22682),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1357_3_lut_LC_23_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1357_3_lut_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1357_3_lut_LC_23_19_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1357_3_lut_LC_23_19_4  (
            .in0(_gnd_net_),
            .in1(N__21674),
            .in2(N__22943),
            .in3(N__23359),
            .lcout(\eeprom.n2113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1362_3_lut_LC_23_19_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1362_3_lut_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1362_3_lut_LC_23_19_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1362_3_lut_LC_23_19_5  (
            .in0(N__21615),
            .in1(_gnd_net_),
            .in2(N__23366),
            .in3(N__21668),
            .lcout(\eeprom.n2118 ),
            .ltout(\eeprom.n2118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_50_LC_23_19_6 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_50_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_50_LC_23_19_6 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_50_LC_23_19_6  (
            .in0(N__24634),
            .in1(N__21659),
            .in2(N__21650),
            .in3(N__23264),
            .lcout(\eeprom.n4788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1424_3_lut_LC_23_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1424_3_lut_LC_23_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1424_3_lut_LC_23_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1424_3_lut_LC_23_19_7  (
            .in0(N__22742),
            .in1(N__23284),
            .in2(_gnd_net_),
            .in3(N__23145),
            .lcout(\eeprom.n2212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i24_3_lut_LC_23_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i24_3_lut_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i24_3_lut_LC_23_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i24_3_lut_LC_23_20_0  (
            .in0(N__26429),
            .in1(N__29208),
            .in2(_gnd_net_),
            .in3(N__24983),
            .lcout(\eeprom.n2019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i5_3_lut_LC_23_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i5_3_lut_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i5_3_lut_LC_23_20_1 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \eeprom.rem_4_mux_3_i5_3_lut_LC_23_20_1  (
            .in0(N__29212),
            .in1(_gnd_net_),
            .in2(N__25835),
            .in3(N__24763),
            .lcout(\eeprom.n3721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i8_3_lut_LC_23_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i8_3_lut_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i8_3_lut_LC_23_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i8_3_lut_LC_23_20_2  (
            .in0(N__26096),
            .in1(N__29210),
            .in2(_gnd_net_),
            .in3(N__25544),
            .lcout(\eeprom.n3619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i22_3_lut_LC_23_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i22_3_lut_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i22_3_lut_LC_23_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i22_3_lut_LC_23_20_3  (
            .in0(N__29209),
            .in1(N__26150),
            .in2(_gnd_net_),
            .in3(N__25025),
            .lcout(\eeprom.n2219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i3_3_lut_LC_23_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i3_3_lut_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i3_3_lut_LC_23_20_4 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i3_3_lut_LC_23_20_4  (
            .in0(N__25883),
            .in1(N__29211),
            .in2(_gnd_net_),
            .in3(N__24808),
            .lcout(\eeprom.n3723 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_53_LC_23_20_6 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_53_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_53_LC_23_20_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_adj_53_LC_23_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23089),
            .in3(N__21954),
            .lcout(\eeprom.n6_adj_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1631_3_lut_LC_23_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1631_3_lut_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1631_3_lut_LC_23_21_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1631_3_lut_LC_23_21_0  (
            .in0(_gnd_net_),
            .in1(N__21932),
            .in2(N__23490),
            .in3(N__21926),
            .lcout(\eeprom.n2515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1633_3_lut_LC_23_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1633_3_lut_LC_23_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1633_3_lut_LC_23_21_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1633_3_lut_LC_23_21_1  (
            .in0(_gnd_net_),
            .in1(N__21893),
            .in2(N__21887),
            .in3(N__23467),
            .lcout(\eeprom.n2517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1625_3_lut_LC_23_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1625_3_lut_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1625_3_lut_LC_23_21_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1625_3_lut_LC_23_21_3  (
            .in0(_gnd_net_),
            .in1(N__21857),
            .in2(N__21848),
            .in3(N__23475),
            .lcout(\eeprom.n2509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1623_3_lut_LC_23_21_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1623_3_lut_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1623_3_lut_LC_23_21_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1623_3_lut_LC_23_21_4  (
            .in0(_gnd_net_),
            .in1(N__21821),
            .in2(N__23492),
            .in3(N__21797),
            .lcout(\eeprom.n2507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1634_3_lut_LC_23_21_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1634_3_lut_LC_23_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1634_3_lut_LC_23_21_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_i1634_3_lut_LC_23_21_5  (
            .in0(N__22442),
            .in1(N__21788),
            .in2(_gnd_net_),
            .in3(N__23466),
            .lcout(\eeprom.n2518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1632_3_lut_LC_23_21_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1632_3_lut_LC_23_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1632_3_lut_LC_23_21_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1632_3_lut_LC_23_21_6  (
            .in0(_gnd_net_),
            .in1(N__21779),
            .in2(N__23491),
            .in3(N__21773),
            .lcout(\eeprom.n2516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1630_3_lut_LC_23_21_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1630_3_lut_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1630_3_lut_LC_23_21_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1630_3_lut_LC_23_21_7  (
            .in0(_gnd_net_),
            .in1(N__22118),
            .in2(N__22112),
            .in3(N__23474),
            .lcout(\eeprom.n2514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1695_3_lut_LC_23_22_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1695_3_lut_LC_23_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1695_3_lut_LC_23_22_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1695_3_lut_LC_23_22_0  (
            .in0(N__24019),
            .in1(_gnd_net_),
            .in2(N__24432),
            .in3(N__24002),
            .lcout(\eeprom.n2611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1701_3_lut_LC_23_22_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1701_3_lut_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1701_3_lut_LC_23_22_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1701_3_lut_LC_23_22_1  (
            .in0(_gnd_net_),
            .in1(N__23681),
            .in2(N__23707),
            .in3(N__24408),
            .lcout(\eeprom.n2617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_66_LC_23_22_2 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_66_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_66_LC_23_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_adj_66_LC_23_22_2  (
            .in0(N__24493),
            .in1(N__23907),
            .in2(N__24355),
            .in3(N__24462),
            .lcout(),
            .ltout(\eeprom.n13_adj_329_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_adj_69_LC_23_22_3 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_adj_69_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_adj_69_LC_23_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_adj_69_LC_23_22_3  (
            .in0(N__23989),
            .in1(N__24018),
            .in2(N__22079),
            .in3(N__23882),
            .lcout(\eeprom.n2539 ),
            .ltout(\eeprom.n2539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1697_3_lut_LC_23_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1697_3_lut_LC_23_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1697_3_lut_LC_23_22_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1697_3_lut_LC_23_22_4  (
            .in0(_gnd_net_),
            .in1(N__24094),
            .in2(N__22076),
            .in3(N__24074),
            .lcout(\eeprom.n2613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1767_3_lut_LC_23_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1767_3_lut_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1767_3_lut_LC_23_22_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1767_3_lut_LC_23_22_5  (
            .in0(_gnd_net_),
            .in1(N__23752),
            .in2(N__22073),
            .in3(N__22564),
            .lcout(\eeprom.n2715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1765_3_lut_LC_23_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1765_3_lut_LC_23_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1765_3_lut_LC_23_22_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1765_3_lut_LC_23_22_6  (
            .in0(_gnd_net_),
            .in1(N__23782),
            .in2(N__22587),
            .in3(N__22058),
            .lcout(\eeprom.n2713 ),
            .ltout(\eeprom.n2713_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_80_LC_23_22_7 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_80_LC_23_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_80_LC_23_22_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_80_LC_23_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22028),
            .in3(N__22011),
            .lcout(\eeprom.n5213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1696_3_lut_LC_23_23_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1696_3_lut_LC_23_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1696_3_lut_LC_23_23_0 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \eeprom.rem_4_i1696_3_lut_LC_23_23_0  (
            .in0(N__24061),
            .in1(N__24035),
            .in2(N__24436),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2612 ),
            .ltout(\eeprom.n2612_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i7_4_lut_adj_74_LC_23_23_1 .C_ON=1'b0;
    defparam \eeprom.i7_4_lut_adj_74_LC_23_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i7_4_lut_adj_74_LC_23_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i7_4_lut_adj_74_LC_23_23_1  (
            .in0(N__22329),
            .in1(N__22220),
            .in2(N__22313),
            .in3(N__22308),
            .lcout(\eeprom.n16_adj_334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_23_23_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_23_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_23_23_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_23_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24920),
            .in3(_gnd_net_),
            .lcout(\eeprom.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_adj_73_LC_23_23_4 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_adj_73_LC_23_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_adj_73_LC_23_23_4 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \eeprom.i3_4_lut_adj_73_LC_23_23_4  (
            .in0(N__24287),
            .in1(N__22134),
            .in2(N__23732),
            .in3(N__22274),
            .lcout(\eeprom.n12_adj_333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1690_3_lut_LC_23_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1690_3_lut_LC_23_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1690_3_lut_LC_23_23_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1690_3_lut_LC_23_23_5  (
            .in0(_gnd_net_),
            .in1(N__24470),
            .in2(N__24449),
            .in3(N__24422),
            .lcout(\eeprom.n2606 ),
            .ltout(\eeprom.n2606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_72_LC_23_23_6 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_72_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_72_LC_23_23_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \eeprom.i1_2_lut_adj_72_LC_23_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22223),
            .in3(N__24331),
            .lcout(\eeprom.n10_adj_332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_82_LC_23_23_7 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_82_LC_23_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_82_LC_23_23_7 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_82_LC_23_23_7  (
            .in0(N__22486),
            .in1(N__22214),
            .in2(N__22190),
            .in3(N__22181),
            .lcout(\eeprom.n4830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1766_3_lut_LC_23_24_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1766_3_lut_LC_23_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1766_3_lut_LC_23_24_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1766_3_lut_LC_23_24_1  (
            .in0(_gnd_net_),
            .in1(N__22169),
            .in2(N__23875),
            .in3(N__22561),
            .lcout(\eeprom.n2714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1693_3_lut_LC_23_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1693_3_lut_LC_23_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1693_3_lut_LC_23_24_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1693_3_lut_LC_23_24_2  (
            .in0(_gnd_net_),
            .in1(N__23927),
            .in2(N__23954),
            .in3(N__24427),
            .lcout(\eeprom.n2609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i11_3_lut_LC_23_24_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i11_3_lut_LC_23_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i11_3_lut_LC_23_24_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i11_3_lut_LC_23_24_4  (
            .in0(N__26051),
            .in1(N__29204),
            .in2(_gnd_net_),
            .in3(N__25625),
            .lcout(\eeprom.n3319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1692_3_lut_LC_23_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1692_3_lut_LC_23_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1692_3_lut_LC_23_24_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1692_3_lut_LC_23_24_5  (
            .in0(N__23917),
            .in1(_gnd_net_),
            .in2(N__24437),
            .in3(N__23894),
            .lcout(\eeprom.n2608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1691_3_lut_LC_23_24_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1691_3_lut_LC_23_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1691_3_lut_LC_23_24_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1691_3_lut_LC_23_24_6  (
            .in0(_gnd_net_),
            .in1(N__24508),
            .in2(N__24482),
            .in3(N__24431),
            .lcout(\eeprom.n2607 ),
            .ltout(\eeprom.n2607_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1758_3_lut_LC_23_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1758_3_lut_LC_23_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1758_3_lut_LC_23_24_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i1758_3_lut_LC_23_24_7  (
            .in0(N__22604),
            .in1(_gnd_net_),
            .in2(N__22595),
            .in3(N__22562),
            .lcout(\eeprom.n2706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i17_3_lut_LC_23_25_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i17_3_lut_LC_23_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i17_3_lut_LC_23_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i17_3_lut_LC_23_25_1  (
            .in0(N__29176),
            .in1(N__26258),
            .in2(_gnd_net_),
            .in3(N__24956),
            .lcout(\eeprom.n2719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i15_3_lut_LC_23_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i15_3_lut_LC_23_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i15_3_lut_LC_23_25_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i15_3_lut_LC_23_25_2  (
            .in0(N__25967),
            .in1(N__29177),
            .in2(_gnd_net_),
            .in3(N__27581),
            .lcout(\eeprom.n2919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i20_3_lut_LC_23_25_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i20_3_lut_LC_23_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i20_3_lut_LC_23_25_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i20_3_lut_LC_23_25_4  (
            .in0(N__26201),
            .in1(N__29175),
            .in2(_gnd_net_),
            .in3(N__29348),
            .lcout(\eeprom.n2419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i13_3_lut_LC_23_26_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i13_3_lut_LC_23_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i13_3_lut_LC_23_26_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i13_3_lut_LC_23_26_1  (
            .in0(N__26012),
            .in1(N__29207),
            .in2(_gnd_net_),
            .in3(N__25691),
            .lcout(\eeprom.n3119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_2_lut_LC_24_17_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_2_lut_LC_24_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_2_lut_LC_24_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_2_lut_LC_24_17_0  (
            .in0(_gnd_net_),
            .in1(N__24633),
            .in2(_gnd_net_),
            .in3(N__22361),
            .lcout(\eeprom.n2186 ),
            .ltout(),
            .carryin(bfn_24_17_0_),
            .carryout(\eeprom.n3988 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_3_lut_LC_24_17_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_3_lut_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_3_lut_LC_24_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_3_lut_LC_24_17_1  (
            .in0(_gnd_net_),
            .in1(N__28031),
            .in2(N__22916),
            .in3(N__22886),
            .lcout(\eeprom.n2185 ),
            .ltout(),
            .carryin(\eeprom.n3988 ),
            .carryout(\eeprom.n3989 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_4_lut_LC_24_17_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_4_lut_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_4_lut_LC_24_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_4_lut_LC_24_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22883),
            .in3(N__22847),
            .lcout(\eeprom.n2184 ),
            .ltout(),
            .carryin(\eeprom.n3989 ),
            .carryout(\eeprom.n3990 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_5_lut_LC_24_17_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_5_lut_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_5_lut_LC_24_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_5_lut_LC_24_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22837),
            .in3(N__22796),
            .lcout(\eeprom.n2183 ),
            .ltout(),
            .carryin(\eeprom.n3990 ),
            .carryout(\eeprom.n3991 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_6_lut_LC_24_17_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_6_lut_LC_24_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_6_lut_LC_24_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_6_lut_LC_24_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23314),
            .in3(N__22781),
            .lcout(\eeprom.n2182 ),
            .ltout(),
            .carryin(\eeprom.n3991 ),
            .carryout(\eeprom.n3992 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_7_lut_LC_24_17_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_7_lut_LC_24_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_7_lut_LC_24_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_7_lut_LC_24_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22778),
            .in3(N__22745),
            .lcout(\eeprom.n2181 ),
            .ltout(),
            .carryin(\eeprom.n3992 ),
            .carryout(\eeprom.n3993 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_8_lut_LC_24_17_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_8_lut_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_8_lut_LC_24_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_8_lut_LC_24_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23288),
            .in3(N__22733),
            .lcout(\eeprom.n2180 ),
            .ltout(),
            .carryin(\eeprom.n3993 ),
            .carryout(\eeprom.n3994 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_9_lut_LC_24_17_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_9_lut_LC_24_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_9_lut_LC_24_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_9_lut_LC_24_17_7  (
            .in0(_gnd_net_),
            .in1(N__28032),
            .in2(N__22725),
            .in3(N__22685),
            .lcout(\eeprom.n2179 ),
            .ltout(),
            .carryin(\eeprom.n3994 ),
            .carryout(\eeprom.n3995 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_10_lut_LC_24_18_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1419_10_lut_LC_24_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_10_lut_LC_24_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1419_10_lut_LC_24_18_0  (
            .in0(_gnd_net_),
            .in1(N__28318),
            .in2(N__23027),
            .in3(N__22673),
            .lcout(\eeprom.n2178 ),
            .ltout(),
            .carryin(bfn_24_18_0_),
            .carryout(\eeprom.n3996 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1419_11_lut_LC_24_18_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1419_11_lut_LC_24_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1419_11_lut_LC_24_18_1 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1419_11_lut_LC_24_18_1  (
            .in0(N__28319),
            .in1(N__23168),
            .in2(N__23156),
            .in3(N__23093),
            .lcout(\eeprom.n2209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i2_3_lut_LC_24_18_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i2_3_lut_LC_24_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i2_3_lut_LC_24_18_2 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i2_3_lut_LC_24_18_2  (
            .in0(N__25916),
            .in1(N__29213),
            .in2(_gnd_net_),
            .in3(N__25663),
            .lcout(\eeprom.n3724 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1291_3_lut_LC_24_18_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1291_3_lut_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1291_3_lut_LC_24_18_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1291_3_lut_LC_24_18_4  (
            .in0(_gnd_net_),
            .in1(N__23180),
            .in2(N__25739),
            .in3(N__23596),
            .lcout(\eeprom.n2015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1355_3_lut_LC_24_18_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1355_3_lut_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1355_3_lut_LC_24_18_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \eeprom.rem_4_i1355_3_lut_LC_24_18_6  (
            .in0(N__23357),
            .in1(N__23230),
            .in2(N__23036),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1294_3_lut_LC_24_18_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1294_3_lut_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1294_3_lut_LC_24_18_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1294_3_lut_LC_24_18_7  (
            .in0(N__25145),
            .in1(_gnd_net_),
            .in2(N__23605),
            .in3(N__23210),
            .lcout(\eeprom.n2018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3487_4_lut_LC_24_19_0 .C_ON=1'b0;
    defparam \eeprom.i3487_4_lut_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3487_4_lut_LC_24_19_0 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \eeprom.i3487_4_lut_LC_24_19_0  (
            .in0(N__25144),
            .in1(N__25459),
            .in2(N__25520),
            .in3(N__25703),
            .lcout(\eeprom.n1945 ),
            .ltout(\eeprom.n1945_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1293_3_lut_LC_24_19_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1293_3_lut_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1293_3_lut_LC_24_19_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.rem_4_i1293_3_lut_LC_24_19_1  (
            .in0(N__23198),
            .in1(_gnd_net_),
            .in2(N__22982),
            .in3(N__25519),
            .lcout(\eeprom.n2017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1290_3_lut_LC_24_19_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1290_3_lut_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1290_3_lut_LC_24_19_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \eeprom.rem_4_i1290_3_lut_LC_24_19_2  (
            .in0(N__27808),
            .in1(_gnd_net_),
            .in2(N__23603),
            .in3(N__23636),
            .lcout(\eeprom.n2014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1292_3_lut_LC_24_19_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1292_3_lut_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1292_3_lut_LC_24_19_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1292_3_lut_LC_24_19_3  (
            .in0(_gnd_net_),
            .in1(N__23189),
            .in2(N__27701),
            .in3(N__23588),
            .lcout(\eeprom.n2016 ),
            .ltout(\eeprom.n2016_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1359_3_lut_LC_24_19_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1359_3_lut_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1359_3_lut_LC_24_19_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.rem_4_i1359_3_lut_LC_24_19_4  (
            .in0(_gnd_net_),
            .in1(N__23375),
            .in2(N__23369),
            .in3(N__23365),
            .lcout(\eeprom.n2115 ),
            .ltout(\eeprom.n2115_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_48_LC_24_19_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_48_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_48_LC_24_19_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_48_LC_24_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23291),
            .in3(N__23280),
            .lcout(\eeprom.n5059 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4674_3_lut_LC_24_19_6 .C_ON=1'b0;
    defparam \eeprom.i4674_3_lut_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4674_3_lut_LC_24_19_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \eeprom.i4674_3_lut_LC_24_19_6  (
            .in0(N__23627),
            .in1(_gnd_net_),
            .in2(N__23604),
            .in3(N__27613),
            .lcout(\eeprom.n2013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1288_3_lut_LC_24_19_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1288_3_lut_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1288_3_lut_LC_24_19_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1288_3_lut_LC_24_19_7  (
            .in0(_gnd_net_),
            .in1(N__25568),
            .in2(N__23618),
            .in3(N__23592),
            .lcout(\eeprom.n2012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_2_lut_LC_24_20_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_2_lut_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_2_lut_LC_24_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_2_lut_LC_24_20_0  (
            .in0(_gnd_net_),
            .in1(N__25143),
            .in2(_gnd_net_),
            .in3(N__23201),
            .lcout(\eeprom.n1986 ),
            .ltout(),
            .carryin(bfn_24_20_0_),
            .carryout(\eeprom.n3973 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_3_lut_LC_24_20_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_3_lut_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_3_lut_LC_24_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_3_lut_LC_24_20_1  (
            .in0(_gnd_net_),
            .in1(N__25515),
            .in2(N__28594),
            .in3(N__23192),
            .lcout(\eeprom.n1985 ),
            .ltout(),
            .carryin(\eeprom.n3973 ),
            .carryout(\eeprom.n3974 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_4_lut_LC_24_20_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_4_lut_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_4_lut_LC_24_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_4_lut_LC_24_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27700),
            .in3(N__23183),
            .lcout(\eeprom.n1984 ),
            .ltout(),
            .carryin(\eeprom.n3974 ),
            .carryout(\eeprom.n3975 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_5_lut_LC_24_20_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_5_lut_LC_24_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_5_lut_LC_24_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_5_lut_LC_24_20_3  (
            .in0(_gnd_net_),
            .in1(N__25735),
            .in2(_gnd_net_),
            .in3(N__23171),
            .lcout(\eeprom.n1983 ),
            .ltout(),
            .carryin(\eeprom.n3975 ),
            .carryout(\eeprom.n3976 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_6_lut_LC_24_20_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_6_lut_LC_24_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_6_lut_LC_24_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_6_lut_LC_24_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27809),
            .in3(N__23630),
            .lcout(\eeprom.n1982 ),
            .ltout(),
            .carryin(\eeprom.n3976 ),
            .carryout(\eeprom.n3977 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_7_lut_LC_24_20_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_7_lut_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_7_lut_LC_24_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_7_lut_LC_24_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27614),
            .in3(N__23621),
            .lcout(\eeprom.n1981 ),
            .ltout(),
            .carryin(\eeprom.n3977 ),
            .carryout(\eeprom.n3978 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_8_lut_LC_24_20_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1285_8_lut_LC_24_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_8_lut_LC_24_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1285_8_lut_LC_24_20_6  (
            .in0(_gnd_net_),
            .in1(N__25564),
            .in2(_gnd_net_),
            .in3(N__23609),
            .lcout(\eeprom.n1980 ),
            .ltout(),
            .carryin(\eeprom.n3978 ),
            .carryout(\eeprom.n3979 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1285_9_lut_LC_24_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1285_9_lut_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1285_9_lut_LC_24_20_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \eeprom.rem_4_add_1285_9_lut_LC_24_20_7  (
            .in0(N__28477),
            .in1(N__25460),
            .in2(N__23606),
            .in3(N__23564),
            .lcout(\eeprom.n2011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1626_3_lut_LC_24_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1626_3_lut_LC_24_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1626_3_lut_LC_24_21_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1626_3_lut_LC_24_21_0  (
            .in0(_gnd_net_),
            .in1(N__23540),
            .in2(N__23510),
            .in3(N__23494),
            .lcout(\eeprom.n2510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i10_3_lut_LC_24_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i10_3_lut_LC_24_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i10_3_lut_LC_24_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \eeprom.rem_4_mux_3_i10_3_lut_LC_24_21_3  (
            .in0(N__29738),
            .in1(N__26078),
            .in2(_gnd_net_),
            .in3(N__29199),
            .lcout(\eeprom.n3419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_63_LC_24_21_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_63_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_63_LC_24_21_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_63_LC_24_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24130),
            .in3(N__24057),
            .lcout(),
            .ltout(\eeprom.n5169_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_64_LC_24_21_6 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_64_LC_24_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_64_LC_24_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_64_LC_24_21_6  (
            .in0(N__24093),
            .in1(N__23664),
            .in2(N__23396),
            .in3(N__24162),
            .lcout(),
            .ltout(\eeprom.n5173_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i3_4_lut_adj_65_LC_24_21_7 .C_ON=1'b0;
    defparam \eeprom.i3_4_lut_adj_65_LC_24_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i3_4_lut_adj_65_LC_24_21_7 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \eeprom.i3_4_lut_adj_65_LC_24_21_7  (
            .in0(N__24319),
            .in1(N__23940),
            .in2(N__23885),
            .in3(N__23700),
            .lcout(\eeprom.n11_adj_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1700_3_lut_LC_24_22_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1700_3_lut_LC_24_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1700_3_lut_LC_24_22_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \eeprom.rem_4_i1700_3_lut_LC_24_22_2  (
            .in0(N__24418),
            .in1(N__23645),
            .in2(N__23671),
            .in3(_gnd_net_),
            .lcout(\eeprom.n2616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1698_3_lut_LC_24_22_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1698_3_lut_LC_24_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1698_3_lut_LC_24_22_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \eeprom.rem_4_i1698_3_lut_LC_24_22_3  (
            .in0(N__24107),
            .in1(N__24129),
            .in2(_gnd_net_),
            .in3(N__24417),
            .lcout(\eeprom.n2614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1699_3_lut_LC_24_22_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1699_3_lut_LC_24_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1699_3_lut_LC_24_22_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1699_3_lut_LC_24_22_4  (
            .in0(_gnd_net_),
            .in1(N__24163),
            .in2(N__24435),
            .in3(N__24143),
            .lcout(\eeprom.n2615 ),
            .ltout(\eeprom.n2615_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_70_LC_24_22_5 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_70_LC_24_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_70_LC_24_22_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_70_LC_24_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23849),
            .in3(N__23832),
            .lcout(),
            .ltout(\eeprom.n5101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_71_LC_24_22_6 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_71_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_71_LC_24_22_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_71_LC_24_22_6  (
            .in0(N__23805),
            .in1(N__23778),
            .in2(N__23762),
            .in3(N__23748),
            .lcout(\eeprom.n5105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_2_lut_LC_24_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_2_lut_LC_24_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_2_lut_LC_24_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_2_lut_LC_24_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24312),
            .in3(N__23711),
            .lcout(\eeprom.n2586 ),
            .ltout(),
            .carryin(bfn_24_23_0_),
            .carryout(\eeprom.n4030 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_3_lut_LC_24_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_3_lut_LC_24_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_3_lut_LC_24_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_3_lut_LC_24_23_1  (
            .in0(_gnd_net_),
            .in1(N__28478),
            .in2(N__23708),
            .in3(N__23675),
            .lcout(\eeprom.n2585 ),
            .ltout(),
            .carryin(\eeprom.n4030 ),
            .carryout(\eeprom.n4031 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_4_lut_LC_24_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_4_lut_LC_24_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_4_lut_LC_24_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_4_lut_LC_24_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23672),
            .in3(N__23639),
            .lcout(\eeprom.n2584 ),
            .ltout(),
            .carryin(\eeprom.n4031 ),
            .carryout(\eeprom.n4032 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_5_lut_LC_24_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_5_lut_LC_24_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_5_lut_LC_24_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_5_lut_LC_24_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24167),
            .in3(N__24137),
            .lcout(\eeprom.n2583 ),
            .ltout(),
            .carryin(\eeprom.n4032 ),
            .carryout(\eeprom.n4033 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_6_lut_LC_24_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_6_lut_LC_24_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_6_lut_LC_24_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_6_lut_LC_24_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24134),
            .in3(N__24101),
            .lcout(\eeprom.n2582 ),
            .ltout(),
            .carryin(\eeprom.n4033 ),
            .carryout(\eeprom.n4034 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_7_lut_LC_24_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_7_lut_LC_24_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_7_lut_LC_24_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_7_lut_LC_24_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24098),
            .in3(N__24068),
            .lcout(\eeprom.n2581 ),
            .ltout(),
            .carryin(\eeprom.n4034 ),
            .carryout(\eeprom.n4035 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_8_lut_LC_24_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_8_lut_LC_24_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_8_lut_LC_24_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_8_lut_LC_24_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24065),
            .in3(N__24029),
            .lcout(\eeprom.n2580 ),
            .ltout(),
            .carryin(\eeprom.n4035 ),
            .carryout(\eeprom.n4036 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_9_lut_LC_24_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_9_lut_LC_24_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_9_lut_LC_24_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_9_lut_LC_24_23_7  (
            .in0(_gnd_net_),
            .in1(N__28479),
            .in2(N__24026),
            .in3(N__23996),
            .lcout(\eeprom.n2579 ),
            .ltout(),
            .carryin(\eeprom.n4036 ),
            .carryout(\eeprom.n4037 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_10_lut_LC_24_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_10_lut_LC_24_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_10_lut_LC_24_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_10_lut_LC_24_24_0  (
            .in0(_gnd_net_),
            .in1(N__28595),
            .in2(N__23993),
            .in3(N__23957),
            .lcout(\eeprom.n2578 ),
            .ltout(),
            .carryin(bfn_24_24_0_),
            .carryout(\eeprom.n4038 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_11_lut_LC_24_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_11_lut_LC_24_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_11_lut_LC_24_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_11_lut_LC_24_24_1  (
            .in0(_gnd_net_),
            .in1(N__23947),
            .in2(N__28717),
            .in3(N__23921),
            .lcout(\eeprom.n2577 ),
            .ltout(),
            .carryin(\eeprom.n4038 ),
            .carryout(\eeprom.n4039 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_12_lut_LC_24_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_12_lut_LC_24_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_12_lut_LC_24_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_12_lut_LC_24_24_2  (
            .in0(_gnd_net_),
            .in1(N__28599),
            .in2(N__23918),
            .in3(N__23888),
            .lcout(\eeprom.n2576 ),
            .ltout(),
            .carryin(\eeprom.n4039 ),
            .carryout(\eeprom.n4040 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_13_lut_LC_24_24_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_13_lut_LC_24_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_13_lut_LC_24_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_13_lut_LC_24_24_3  (
            .in0(_gnd_net_),
            .in1(N__28500),
            .in2(N__24509),
            .in3(N__24473),
            .lcout(\eeprom.n2575 ),
            .ltout(),
            .carryin(\eeprom.n4040 ),
            .carryout(\eeprom.n4041 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_14_lut_LC_24_24_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_add_1687_14_lut_LC_24_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_14_lut_LC_24_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_add_1687_14_lut_LC_24_24_4  (
            .in0(_gnd_net_),
            .in1(N__24469),
            .in2(N__28632),
            .in3(N__24440),
            .lcout(\eeprom.n2574 ),
            .ltout(),
            .carryin(\eeprom.n4041 ),
            .carryout(\eeprom.n4042 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_add_1687_15_lut_LC_24_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_add_1687_15_lut_LC_24_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_add_1687_15_lut_LC_24_24_5 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \eeprom.rem_4_add_1687_15_lut_LC_24_24_5  (
            .in0(N__28600),
            .in1(N__24426),
            .in2(N__24362),
            .in3(N__24338),
            .lcout(\eeprom.n2605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i19_3_lut_LC_24_24_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i19_3_lut_LC_24_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i19_3_lut_LC_24_24_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i19_3_lut_LC_24_24_7  (
            .in0(N__26216),
            .in1(N__29198),
            .in2(_gnd_net_),
            .in3(N__25103),
            .lcout(\eeprom.n2519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i18_3_lut_LC_24_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i18_3_lut_LC_24_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i18_3_lut_LC_24_25_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i18_3_lut_LC_24_25_2  (
            .in0(N__26237),
            .in1(N__29178),
            .in2(_gnd_net_),
            .in3(N__25076),
            .lcout(\eeprom.n2619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i16_3_lut_LC_24_25_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i16_3_lut_LC_24_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i16_3_lut_LC_24_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i16_3_lut_LC_24_25_3  (
            .in0(N__29179),
            .in1(N__26282),
            .in2(_gnd_net_),
            .in3(N__29984),
            .lcout(\eeprom.n2819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i12_3_lut_LC_24_25_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i12_3_lut_LC_24_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i12_3_lut_LC_24_25_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i12_3_lut_LC_24_25_4  (
            .in0(N__26039),
            .in1(N__29180),
            .in2(_gnd_net_),
            .in3(N__29549),
            .lcout(\eeprom.n3219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i14_3_lut_LC_24_26_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i14_3_lut_LC_24_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i14_3_lut_LC_24_26_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i14_3_lut_LC_24_26_5  (
            .in0(N__25982),
            .in1(N__29203),
            .in2(_gnd_net_),
            .in3(N__24860),
            .lcout(\eeprom.n3019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_9_LC_26_17_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_9_LC_26_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_9_LC_26_17_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_adj_9_LC_26_17_0  (
            .in0(N__27423),
            .in1(N__27143),
            .in2(_gnd_net_),
            .in3(N__26886),
            .lcout(\eeprom.i2c.n534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3200_2_lut_LC_26_17_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i3200_2_lut_LC_26_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3200_2_lut_LC_26_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i3200_2_lut_LC_26_17_1  (
            .in0(_gnd_net_),
            .in1(N__26986),
            .in2(_gnd_net_),
            .in3(N__27028),
            .lcout(n3585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_10_LC_26_17_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_10_LC_26_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_10_LC_26_17_2 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_adj_10_LC_26_17_2  (
            .in0(N__25245),
            .in1(N__25168),
            .in2(_gnd_net_),
            .in3(N__26948),
            .lcout(n1805),
            .ltout(n1805_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i1_LC_26_17_3 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i1_LC_26_17_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i1_LC_26_17_3 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \eeprom.i2c.data_out_i0_i1_LC_26_17_3  (
            .in0(N__24542),
            .in1(N__26560),
            .in2(N__24545),
            .in3(N__26521),
            .lcout(n170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29694),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_26_17_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_26_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_26_17_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_26_17_4  (
            .in0(N__25246),
            .in1(N__25169),
            .in2(_gnd_net_),
            .in3(N__26949),
            .lcout(n1800),
            .ltout(n1800_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i4_LC_26_17_5 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i4_LC_26_17_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i4_LC_26_17_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \eeprom.i2c.data_out_i0_i4_LC_26_17_5  (
            .in0(N__24533),
            .in1(N__24527),
            .in2(N__24536),
            .in3(N__26522),
            .lcout(n164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29694),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_36_i4_2_lut_LC_26_17_6 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_36_i4_2_lut_LC_26_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_36_i4_2_lut_LC_26_17_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \eeprom.i2c.equal_36_i4_2_lut_LC_26_17_6  (
            .in0(N__26987),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27032),
            .lcout(n4_adj_361),
            .ltout(n4_adj_361_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i5_LC_26_17_7 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i5_LC_26_17_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i5_LC_26_17_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \eeprom.i2c.data_out_i0_i5_LC_26_17_7  (
            .in0(N__24705),
            .in1(N__24518),
            .in2(N__24521),
            .in3(N__26523),
            .lcout(n162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29694),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4589_3_lut_4_lut_4_lut_LC_26_18_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i4589_3_lut_4_lut_4_lut_LC_26_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4589_3_lut_4_lut_4_lut_LC_26_18_0 .LUT_INIT=16'b1110110111111111;
    LogicCell40 \eeprom.i2c.i4589_3_lut_4_lut_4_lut_LC_26_18_0  (
            .in0(N__27152),
            .in1(N__27516),
            .in2(N__26897),
            .in3(N__27419),
            .lcout(),
            .ltout(n5361_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_26_18_1.C_ON=1'b0;
    defparam i3_4_lut_LC_26_18_1.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_26_18_1.LUT_INIT=16'b1110000011110000;
    LogicCell40 i3_4_lut_LC_26_18_1 (
            .in0(N__26498),
            .in1(N__25183),
            .in2(N__24512),
            .in3(N__27884),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i0_LC_26_18_3 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i0_LC_26_18_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i0_LC_26_18_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \eeprom.i2c.data_out_i0_i0_LC_26_18_3  (
            .in0(N__26499),
            .in1(N__24670),
            .in2(N__26564),
            .in3(N__24581),
            .lcout(n172),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29688),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_26_18_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_26_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_26_18_4 .LUT_INIT=16'b1111011100110011;
    LogicCell40 \eeprom.i2c.i1_4_lut_4_lut_LC_26_18_4  (
            .in0(N__29785),
            .in1(N__27515),
            .in2(N__26519),
            .in3(N__27418),
            .lcout(),
            .ltout(n22_adj_367_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_26_18_5.C_ON=1'b0;
    defparam i1_4_lut_LC_26_18_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_26_18_5.LUT_INIT=16'b0010001011110010;
    LogicCell40 i1_4_lut_LC_26_18_5 (
            .in0(N__26497),
            .in1(N__25182),
            .in2(N__24575),
            .in3(N__25166),
            .lcout(),
            .ltout(n4_adj_369_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2_3_lut_4_lut_LC_26_18_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i2_3_lut_4_lut_LC_26_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i2_3_lut_4_lut_LC_26_18_6 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \eeprom.i2c.i2_3_lut_4_lut_LC_26_18_6  (
            .in0(N__27153),
            .in1(N__26891),
            .in2(N__24572),
            .in3(N__25247),
            .lcout(n4733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_26_18_7 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_26_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_26_18_7 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_26_18_7  (
            .in0(N__27514),
            .in1(N__27151),
            .in2(N__27424),
            .in3(N__26887),
            .lcout(n11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_38_i4_2_lut_LC_26_19_0 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_38_i4_2_lut_LC_26_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_38_i4_2_lut_LC_26_19_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \eeprom.i2c.equal_38_i4_2_lut_LC_26_19_0  (
            .in0(N__27037),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26993),
            .lcout(n4),
            .ltout(n4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i3_LC_26_19_1 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i3_LC_26_19_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i3_LC_26_19_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \eeprom.i2c.data_out_i0_i3_LC_26_19_1  (
            .in0(N__24566),
            .in1(N__24712),
            .in2(N__24569),
            .in3(N__26514),
            .lcout(n166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29695),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_26_19_2 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_26_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_26_19_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_26_19_2  (
            .in0(_gnd_net_),
            .in1(N__27144),
            .in2(_gnd_net_),
            .in3(N__26893),
            .lcout(n10_adj_360),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i2_LC_26_19_3 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i2_LC_26_19_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i2_LC_26_19_3 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \eeprom.i2c.data_out_i0_i2_LC_26_19_3  (
            .in0(N__24551),
            .in1(N__24676),
            .in2(N__24560),
            .in3(N__26513),
            .lcout(n168),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29695),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i7_LC_26_19_4 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i7_LC_26_19_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i7_LC_26_19_4 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \eeprom.i2c.data_out_i0_i7_LC_26_19_4  (
            .in0(N__24692),
            .in1(N__24658),
            .in2(N__26524),
            .in3(N__24713),
            .lcout(n158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29695),
            .ce(),
            .sr(_gnd_net_));
    defparam i4649_3_lut_4_lut_LC_26_19_5.C_ON=1'b0;
    defparam i4649_3_lut_4_lut_LC_26_19_5.SEQ_MODE=4'b0000;
    defparam i4649_3_lut_4_lut_LC_26_19_5.LUT_INIT=16'b1111111011111011;
    LogicCell40 i4649_3_lut_4_lut_LC_26_19_5 (
            .in0(N__26894),
            .in1(N__27425),
            .in2(N__27160),
            .in3(N__27520),
            .lcout(),
            .ltout(n5461_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i1_LC_26_19_6 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i1_LC_26_19_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i1_LC_26_19_6 .LUT_INIT=16'b1010101000111111;
    LogicCell40 \eeprom.i2c.state_i0_i1_LC_26_19_6  (
            .in0(N__27521),
            .in1(N__24686),
            .in2(N__24680),
            .in3(N__27176),
            .lcout(state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29695),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i6_LC_26_19_7 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i6_LC_26_19_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i6_LC_26_19_7 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \eeprom.i2c.data_out_i0_i6_LC_26_19_7  (
            .in0(N__24644),
            .in1(N__24677),
            .in2(N__24659),
            .in3(N__26515),
            .lcout(n160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29695),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i23_3_lut_LC_26_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i23_3_lut_LC_26_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i23_3_lut_LC_26_20_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i23_3_lut_LC_26_20_1  (
            .in0(N__26123),
            .in1(N__29173),
            .in2(_gnd_net_),
            .in3(N__25049),
            .lcout(\eeprom.n2119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_26_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_26_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_26_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_26_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24749),
            .lcout(\eeprom.n29_adj_278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_26_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_26_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_26_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_26_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24856),
            .lcout(\eeprom.n20_adj_259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i21_3_lut_LC_26_20_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i21_3_lut_LC_26_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i21_3_lut_LC_26_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i21_3_lut_LC_26_20_4  (
            .in0(N__29174),
            .in1(N__26174),
            .in2(_gnd_net_),
            .in3(N__24919),
            .lcout(\eeprom.n2319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_26_20_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_26_20_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_26_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_26_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24794),
            .lcout(\eeprom.n31_adj_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i0_LC_26_21_0 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i0_LC_26_21_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i0_LC_26_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i0_LC_26_21_0  (
            .in0(_gnd_net_),
            .in1(N__25485),
            .in2(_gnd_net_),
            .in3(N__24818),
            .lcout(\eeprom.eeprom_counter_0 ),
            .ltout(),
            .carryin(bfn_26_21_0_),
            .carryout(\eeprom.n3931 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i1_LC_26_21_1 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i1_LC_26_21_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i1_LC_26_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i1_LC_26_21_1  (
            .in0(_gnd_net_),
            .in1(N__25653),
            .in2(_gnd_net_),
            .in3(N__24815),
            .lcout(\eeprom.eeprom_counter_1 ),
            .ltout(),
            .carryin(\eeprom.n3931 ),
            .carryout(\eeprom.n3932 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i2_LC_26_21_2 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i2_LC_26_21_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i2_LC_26_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i2_LC_26_21_2  (
            .in0(_gnd_net_),
            .in1(N__24798),
            .in2(_gnd_net_),
            .in3(N__24773),
            .lcout(\eeprom.eeprom_counter_2 ),
            .ltout(),
            .carryin(\eeprom.n3932 ),
            .carryout(\eeprom.n3933 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i3_LC_26_21_3 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i3_LC_26_21_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i3_LC_26_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i3_LC_26_21_3  (
            .in0(_gnd_net_),
            .in1(N__25762),
            .in2(_gnd_net_),
            .in3(N__24770),
            .lcout(\eeprom.eeprom_counter_3 ),
            .ltout(),
            .carryin(\eeprom.n3933 ),
            .carryout(\eeprom.n3934 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i4_LC_26_21_4 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i4_LC_26_21_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i4_LC_26_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i4_LC_26_21_4  (
            .in0(_gnd_net_),
            .in1(N__24753),
            .in2(_gnd_net_),
            .in3(N__24728),
            .lcout(\eeprom.eeprom_counter_4 ),
            .ltout(),
            .carryin(\eeprom.n3934 ),
            .carryout(\eeprom.n3935 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i5_LC_26_21_5 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i5_LC_26_21_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i5_LC_26_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i5_LC_26_21_5  (
            .in0(_gnd_net_),
            .in1(N__25344),
            .in2(_gnd_net_),
            .in3(N__24725),
            .lcout(\eeprom.eeprom_counter_5 ),
            .ltout(),
            .carryin(\eeprom.n3935 ),
            .carryout(\eeprom.n3936 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i6_LC_26_21_6 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i6_LC_26_21_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i6_LC_26_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i6_LC_26_21_6  (
            .in0(_gnd_net_),
            .in1(N__29394),
            .in2(_gnd_net_),
            .in3(N__24722),
            .lcout(\eeprom.eeprom_counter_6 ),
            .ltout(),
            .carryin(\eeprom.n3936 ),
            .carryout(\eeprom.n3937 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i7_LC_26_21_7 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i7_LC_26_21_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i7_LC_26_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i7_LC_26_21_7  (
            .in0(_gnd_net_),
            .in1(N__25540),
            .in2(_gnd_net_),
            .in3(N__24719),
            .lcout(\eeprom.eeprom_counter_7 ),
            .ltout(),
            .carryin(\eeprom.n3937 ),
            .carryout(\eeprom.n3938 ),
            .clk(N__29861),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i8_LC_26_22_0 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i8_LC_26_22_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i8_LC_26_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i8_LC_26_22_0  (
            .in0(_gnd_net_),
            .in1(N__29244),
            .in2(_gnd_net_),
            .in3(N__24716),
            .lcout(\eeprom.eeprom_counter_8 ),
            .ltout(),
            .carryin(bfn_26_22_0_),
            .carryout(\eeprom.n3939 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i9_LC_26_22_1 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i9_LC_26_22_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i9_LC_26_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i9_LC_26_22_1  (
            .in0(_gnd_net_),
            .in1(N__29730),
            .in2(_gnd_net_),
            .in3(N__24872),
            .lcout(\eeprom.eeprom_counter_9 ),
            .ltout(),
            .carryin(\eeprom.n3939 ),
            .carryout(\eeprom.n3940 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i10_LC_26_22_2 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i10_LC_26_22_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i10_LC_26_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i10_LC_26_22_2  (
            .in0(_gnd_net_),
            .in1(N__25621),
            .in2(_gnd_net_),
            .in3(N__24869),
            .lcout(\eeprom.eeprom_counter_10 ),
            .ltout(),
            .carryin(\eeprom.n3940 ),
            .carryout(\eeprom.n3941 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i11_LC_26_22_3 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i11_LC_26_22_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i11_LC_26_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i11_LC_26_22_3  (
            .in0(_gnd_net_),
            .in1(N__29544),
            .in2(_gnd_net_),
            .in3(N__24866),
            .lcout(\eeprom.eeprom_counter_11 ),
            .ltout(),
            .carryin(\eeprom.n3941 ),
            .carryout(\eeprom.n3942 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i12_LC_26_22_4 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i12_LC_26_22_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i12_LC_26_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i12_LC_26_22_4  (
            .in0(_gnd_net_),
            .in1(N__25687),
            .in2(_gnd_net_),
            .in3(N__24863),
            .lcout(\eeprom.eeprom_counter_12 ),
            .ltout(),
            .carryin(\eeprom.n3942 ),
            .carryout(\eeprom.n3943 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i13_LC_26_22_5 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i13_LC_26_22_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i13_LC_26_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i13_LC_26_22_5  (
            .in0(_gnd_net_),
            .in1(N__24855),
            .in2(_gnd_net_),
            .in3(N__24833),
            .lcout(\eeprom.eeprom_counter_13 ),
            .ltout(),
            .carryin(\eeprom.n3943 ),
            .carryout(\eeprom.n3944 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i14_LC_26_22_6 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i14_LC_26_22_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i14_LC_26_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i14_LC_26_22_6  (
            .in0(_gnd_net_),
            .in1(N__27573),
            .in2(_gnd_net_),
            .in3(N__24830),
            .lcout(\eeprom.eeprom_counter_14 ),
            .ltout(),
            .carryin(\eeprom.n3944 ),
            .carryout(\eeprom.n3945 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i15_LC_26_22_7 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i15_LC_26_22_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i15_LC_26_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i15_LC_26_22_7  (
            .in0(_gnd_net_),
            .in1(N__29976),
            .in2(_gnd_net_),
            .in3(N__24827),
            .lcout(\eeprom.eeprom_counter_15 ),
            .ltout(),
            .carryin(\eeprom.n3945 ),
            .carryout(\eeprom.n3946 ),
            .clk(N__29863),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i16_LC_26_23_0 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i16_LC_26_23_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i16_LC_26_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i16_LC_26_23_0  (
            .in0(_gnd_net_),
            .in1(N__24948),
            .in2(_gnd_net_),
            .in3(N__24824),
            .lcout(\eeprom.eeprom_counter_16 ),
            .ltout(),
            .carryin(bfn_26_23_0_),
            .carryout(\eeprom.n3947 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i17_LC_26_23_1 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i17_LC_26_23_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i17_LC_26_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i17_LC_26_23_1  (
            .in0(_gnd_net_),
            .in1(N__25071),
            .in2(_gnd_net_),
            .in3(N__24821),
            .lcout(\eeprom.eeprom_counter_17 ),
            .ltout(),
            .carryin(\eeprom.n3947 ),
            .carryout(\eeprom.n3948 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i18_LC_26_23_2 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i18_LC_26_23_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i18_LC_26_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i18_LC_26_23_2  (
            .in0(_gnd_net_),
            .in1(N__25102),
            .in2(_gnd_net_),
            .in3(N__24926),
            .lcout(\eeprom.eeprom_counter_18 ),
            .ltout(),
            .carryin(\eeprom.n3948 ),
            .carryout(\eeprom.n3949 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i19_LC_26_23_3 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i19_LC_26_23_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i19_LC_26_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i19_LC_26_23_3  (
            .in0(_gnd_net_),
            .in1(N__29340),
            .in2(_gnd_net_),
            .in3(N__24923),
            .lcout(\eeprom.eeprom_counter_19 ),
            .ltout(),
            .carryin(\eeprom.n3949 ),
            .carryout(\eeprom.n3950 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i20_LC_26_23_4 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i20_LC_26_23_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i20_LC_26_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i20_LC_26_23_4  (
            .in0(_gnd_net_),
            .in1(N__24915),
            .in2(_gnd_net_),
            .in3(N__24893),
            .lcout(\eeprom.eeprom_counter_20 ),
            .ltout(),
            .carryin(\eeprom.n3950 ),
            .carryout(\eeprom.n3951 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i21_LC_26_23_5 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i21_LC_26_23_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i21_LC_26_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i21_LC_26_23_5  (
            .in0(_gnd_net_),
            .in1(N__25020),
            .in2(_gnd_net_),
            .in3(N__24890),
            .lcout(\eeprom.eeprom_counter_21 ),
            .ltout(),
            .carryin(\eeprom.n3951 ),
            .carryout(\eeprom.n3952 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i22_LC_26_23_6 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i22_LC_26_23_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i22_LC_26_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i22_LC_26_23_6  (
            .in0(_gnd_net_),
            .in1(N__25044),
            .in2(_gnd_net_),
            .in3(N__24887),
            .lcout(\eeprom.eeprom_counter_22 ),
            .ltout(),
            .carryin(\eeprom.n3952 ),
            .carryout(\eeprom.n3953 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i23_LC_26_23_7 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i23_LC_26_23_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i23_LC_26_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i23_LC_26_23_7  (
            .in0(_gnd_net_),
            .in1(N__24978),
            .in2(_gnd_net_),
            .in3(N__24884),
            .lcout(\eeprom.eeprom_counter_23 ),
            .ltout(),
            .carryin(\eeprom.n3953 ),
            .carryout(\eeprom.n3954 ),
            .clk(N__29865),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i24_LC_26_24_0 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i24_LC_26_24_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i24_LC_26_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i24_LC_26_24_0  (
            .in0(_gnd_net_),
            .in1(N__25120),
            .in2(_gnd_net_),
            .in3(N__24881),
            .lcout(\eeprom.eeprom_counter_24 ),
            .ltout(),
            .carryin(bfn_26_24_0_),
            .carryout(\eeprom.n3955 ),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i25_LC_26_24_1 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i25_LC_26_24_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i25_LC_26_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i25_LC_26_24_1  (
            .in0(_gnd_net_),
            .in1(N__29496),
            .in2(_gnd_net_),
            .in3(N__24878),
            .lcout(\eeprom.eeprom_counter_25 ),
            .ltout(),
            .carryin(\eeprom.n3955 ),
            .carryout(\eeprom.n3956 ),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i26_LC_26_24_2 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i26_LC_26_24_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i26_LC_26_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i26_LC_26_24_2  (
            .in0(_gnd_net_),
            .in1(N__29312),
            .in2(_gnd_net_),
            .in3(N__24875),
            .lcout(\eeprom.eeprom_counter_26 ),
            .ltout(),
            .carryin(\eeprom.n3956 ),
            .carryout(\eeprom.n3957 ),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i27_LC_26_24_3 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i27_LC_26_24_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i27_LC_26_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i27_LC_26_24_3  (
            .in0(_gnd_net_),
            .in1(N__25438),
            .in2(_gnd_net_),
            .in3(N__24998),
            .lcout(\eeprom.eeprom_counter_27 ),
            .ltout(),
            .carryin(\eeprom.n3957 ),
            .carryout(\eeprom.n3958 ),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i28_LC_26_24_4 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i28_LC_26_24_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i28_LC_26_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i28_LC_26_24_4  (
            .in0(_gnd_net_),
            .in1(N__25593),
            .in2(_gnd_net_),
            .in3(N__24995),
            .lcout(\eeprom.eeprom_counter_28 ),
            .ltout(),
            .carryin(\eeprom.n3958 ),
            .carryout(\eeprom.n3959 ),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i29_LC_26_24_5 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i29_LC_26_24_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i29_LC_26_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i29_LC_26_24_5  (
            .in0(_gnd_net_),
            .in1(N__27778),
            .in2(_gnd_net_),
            .in3(N__24992),
            .lcout(\eeprom.eeprom_counter_29 ),
            .ltout(),
            .carryin(\eeprom.n3959 ),
            .carryout(\eeprom.n3960 ),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i30_LC_26_24_6 .C_ON=1'b1;
    defparam \eeprom.eeprom_counter_228__i30_LC_26_24_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i30_LC_26_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i30_LC_26_24_6  (
            .in0(_gnd_net_),
            .in1(N__25300),
            .in2(_gnd_net_),
            .in3(N__24989),
            .lcout(\eeprom.eeprom_counter_30 ),
            .ltout(),
            .carryin(\eeprom.n3960 ),
            .carryout(\eeprom.n3961 ),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.eeprom_counter_228__i31_LC_26_24_7 .C_ON=1'b0;
    defparam \eeprom.eeprom_counter_228__i31_LC_26_24_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.eeprom_counter_228__i31_LC_26_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.eeprom_counter_228__i31_LC_26_24_7  (
            .in0(_gnd_net_),
            .in1(N__29094),
            .in2(_gnd_net_),
            .in3(N__24986),
            .lcout(\eeprom.eeprom_counter_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29866),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_26_25_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_26_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_26_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_26_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27774),
            .lcout(\eeprom.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_26_25_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_26_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_26_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_26_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29304),
            .lcout(\eeprom.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_26_25_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_26_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_26_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_26_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24979),
            .lcout(\eeprom.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_26_25_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_26_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_26_25_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_26_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24955),
            .in3(_gnd_net_),
            .lcout(\eeprom.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_26_25_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_26_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_26_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_26_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25434),
            .lcout(\eeprom.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_26_25_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_26_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_26_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_26_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25296),
            .lcout(\eeprom.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i25_3_lut_LC_26_25_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i25_3_lut_LC_26_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i25_3_lut_LC_26_25_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \eeprom.rem_4_mux_3_i25_3_lut_LC_26_25_6  (
            .in0(_gnd_net_),
            .in1(N__29090),
            .in2(N__26405),
            .in3(N__25119),
            .lcout(\eeprom.n1919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_26_25_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_26_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_26_25_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_26_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25121),
            .in3(_gnd_net_),
            .lcout(\eeprom.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_26_26_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_26_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_26_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_26_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25098),
            .lcout(\eeprom.n15_adj_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_26_26_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_26_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_26_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_26_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25072),
            .lcout(\eeprom.n16_adj_294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_26_26_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_26_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_26_26_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_26_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25045),
            .lcout(\eeprom.n11_adj_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_26_26_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_26_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_26_26_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_26_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25600),
            .in3(_gnd_net_),
            .lcout(\eeprom.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_26_26_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_26_26_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_26_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_26_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29095),
            .lcout(\eeprom.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_26_26_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_26_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_26_26_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_26_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25021),
            .lcout(\eeprom.n12_adj_298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.counter_i0_LC_27_17_0 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i0_LC_27_17_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i0_LC_27_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i0_LC_27_17_0  (
            .in0(_gnd_net_),
            .in1(N__26947),
            .in2(_gnd_net_),
            .in3(N__25208),
            .lcout(\eeprom.i2c.counter_0 ),
            .ltout(),
            .carryin(bfn_27_17_0_),
            .carryout(\eeprom.i2c.n3899 ),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.counter_i1_LC_27_17_1 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i1_LC_27_17_1 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i1_LC_27_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i1_LC_27_17_1  (
            .in0(_gnd_net_),
            .in1(N__28003),
            .in2(N__27038),
            .in3(N__25205),
            .lcout(\eeprom.i2c.counter_1 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3899 ),
            .carryout(\eeprom.i2c.n3900 ),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.counter_i2_LC_27_17_2 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i2_LC_27_17_2 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i2_LC_27_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i2_LC_27_17_2  (
            .in0(_gnd_net_),
            .in1(N__26988),
            .in2(N__28103),
            .in3(N__25202),
            .lcout(\eeprom.i2c.counter_2 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3900 ),
            .carryout(\eeprom.i2c.n3901 ),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.counter_i3_LC_27_17_3 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i3_LC_27_17_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i3_LC_27_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i3_LC_27_17_3  (
            .in0(_gnd_net_),
            .in1(N__28007),
            .in2(N__26645),
            .in3(N__25199),
            .lcout(\eeprom.i2c.counter_3 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3901 ),
            .carryout(\eeprom.i2c.n3902 ),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.counter_i4_LC_27_17_4 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i4_LC_27_17_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i4_LC_27_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i4_LC_27_17_4  (
            .in0(_gnd_net_),
            .in1(N__26615),
            .in2(N__28104),
            .in3(N__25196),
            .lcout(\eeprom.i2c.counter_4 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3902 ),
            .carryout(\eeprom.i2c.n3903 ),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.counter_i5_LC_27_17_5 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i5_LC_27_17_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i5_LC_27_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i5_LC_27_17_5  (
            .in0(_gnd_net_),
            .in1(N__28011),
            .in2(N__26630),
            .in3(N__25193),
            .lcout(\eeprom.i2c.counter_5 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3903 ),
            .carryout(\eeprom.i2c.n3904 ),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.counter_i6_LC_27_17_6 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i6_LC_27_17_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i6_LC_27_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i6_LC_27_17_6  (
            .in0(_gnd_net_),
            .in1(N__26591),
            .in2(N__28105),
            .in3(N__25190),
            .lcout(\eeprom.i2c.counter_6 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3904 ),
            .carryout(\eeprom.i2c.n3905 ),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.counter_i7_LC_27_17_7 .C_ON=1'b0;
    defparam \eeprom.i2c.counter_i7_LC_27_17_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i7_LC_27_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \eeprom.i2c.counter_i7_LC_27_17_7  (
            .in0(N__26603),
            .in1(N__28015),
            .in2(_gnd_net_),
            .in3(N__25187),
            .lcout(\eeprom.i2c.counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29693),
            .ce(N__25256),
            .sr(N__25274));
    defparam \eeprom.i2c.i4657_3_lut_4_lut_LC_27_18_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i4657_3_lut_4_lut_LC_27_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4657_3_lut_4_lut_LC_27_18_0 .LUT_INIT=16'b1111101011001000;
    LogicCell40 \eeprom.i2c.i4657_3_lut_4_lut_LC_27_18_0  (
            .in0(N__25184),
            .in1(N__25167),
            .in2(N__26520),
            .in3(N__25244),
            .lcout(n5458),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i56_3_lut_LC_27_18_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i56_3_lut_LC_27_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i56_3_lut_LC_27_18_1 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \eeprom.i2c.i56_3_lut_LC_27_18_1  (
            .in0(N__27367),
            .in1(N__27129),
            .in2(_gnd_net_),
            .in3(N__26815),
            .lcout(\eeprom.i2c.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i3_LC_27_18_2 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i3_LC_27_18_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i3_LC_27_18_2 .LUT_INIT=16'b1010111110101000;
    LogicCell40 \eeprom.i2c.state_i0_i3_LC_27_18_2  (
            .in0(N__27132),
            .in1(N__26753),
            .in2(N__25223),
            .in3(N__25280),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29689),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3794_2_lut_4_lut_LC_27_18_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i3794_2_lut_4_lut_LC_27_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3794_2_lut_4_lut_LC_27_18_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \eeprom.i2c.i3794_2_lut_4_lut_LC_27_18_3  (
            .in0(N__27369),
            .in1(N__27130),
            .in2(N__26895),
            .in3(N__26446),
            .lcout(\eeprom.i2c.n1913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i20_4_lut_LC_27_18_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i20_4_lut_LC_27_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i20_4_lut_LC_27_18_4 .LUT_INIT=16'b0111010001000100;
    LogicCell40 \eeprom.i2c.i20_4_lut_LC_27_18_4  (
            .in0(N__26447),
            .in1(N__25262),
            .in2(N__26576),
            .in3(N__25415),
            .lcout(\eeprom.i2c.n1829 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_144_i9_2_lut_LC_27_18_5 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_144_i9_2_lut_LC_27_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_144_i9_2_lut_LC_27_18_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \eeprom.i2c.state_7__I_0_144_i9_2_lut_LC_27_18_5  (
            .in0(N__27368),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27513),
            .lcout(\eeprom.i2c.n9 ),
            .ltout(\eeprom.i2c.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_4_lut_LC_27_18_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_4_lut_LC_27_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_4_lut_LC_27_18_6 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \eeprom.i2c.i1_3_lut_4_lut_LC_27_18_6  (
            .in0(N__26572),
            .in1(N__27065),
            .in2(N__25226),
            .in3(N__27055),
            .lcout(n1814),
            .ltout(n1814_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_LC_27_18_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_LC_27_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_LC_27_18_7 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \eeprom.i2c.i1_3_lut_LC_27_18_7  (
            .in0(N__26752),
            .in1(_gnd_net_),
            .in2(N__25211),
            .in3(N__27131),
            .lcout(n471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_adj_8_LC_27_19_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_adj_8_LC_27_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_adj_8_LC_27_19_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \eeprom.i2c.i1_3_lut_adj_8_LC_27_19_0  (
            .in0(N__25400),
            .in1(N__25414),
            .in2(_gnd_net_),
            .in3(N__27526),
            .lcout(\eeprom.i2c.n1901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i321_2_lut_LC_27_19_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i321_2_lut_LC_27_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i321_2_lut_LC_27_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i321_2_lut_LC_27_19_1  (
            .in0(_gnd_net_),
            .in1(N__27301),
            .in2(_gnd_net_),
            .in3(N__26912),
            .lcout(state_7_N_162_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_4_lut_LC_27_19_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_4_lut_LC_27_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_4_lut_LC_27_19_2 .LUT_INIT=16'b0001000100110010;
    LogicCell40 \eeprom.i2c.i1_4_lut_LC_27_19_2  (
            .in0(N__27385),
            .in1(N__27138),
            .in2(N__27522),
            .in3(N__26816),
            .lcout(\eeprom.i2c.n37 ),
            .ltout(\eeprom.i2c.n37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_adj_7_LC_27_19_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_adj_7_LC_27_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_adj_7_LC_27_19_3 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \eeprom.i2c.i1_3_lut_adj_7_LC_27_19_3  (
            .in0(_gnd_net_),
            .in1(N__27493),
            .in2(N__25403),
            .in3(N__25399),
            .lcout(\eeprom.i2c.n39 ),
            .ltout(\eeprom.i2c.n39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4684_4_lut_LC_27_19_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i4684_4_lut_LC_27_19_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4684_4_lut_LC_27_19_4 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \eeprom.i2c.i4684_4_lut_LC_27_19_4  (
            .in0(N__26819),
            .in1(N__27527),
            .in2(N__25391),
            .in3(N__25550),
            .lcout(\eeprom.i2c.n4513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3_4_lut_4_lut_LC_27_19_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i3_4_lut_4_lut_LC_27_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3_4_lut_4_lut_LC_27_19_5 .LUT_INIT=16'b0000010000010100;
    LogicCell40 \eeprom.i2c.i3_4_lut_4_lut_LC_27_19_5  (
            .in0(N__26817),
            .in1(N__27386),
            .in2(N__27159),
            .in3(N__27494),
            .lcout(\eeprom.i2c.n407 ),
            .ltout(\eeprom.i2c.n407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4692_4_lut_LC_27_19_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i4692_4_lut_LC_27_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4692_4_lut_LC_27_19_6 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \eeprom.i2c.i4692_4_lut_LC_27_19_6  (
            .in0(N__27495),
            .in1(N__25388),
            .in2(N__25382),
            .in3(N__26818),
            .lcout(\eeprom.i2c.n524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i1_3_lut_LC_27_20_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i1_3_lut_LC_27_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i1_3_lut_LC_27_20_0 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i1_3_lut_LC_27_20_0  (
            .in0(N__25937),
            .in1(N__29171),
            .in2(_gnd_net_),
            .in3(N__25484),
            .lcout(\eeprom.n917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_27_20_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_27_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_27_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_27_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25340),
            .lcout(\eeprom.n28_adj_279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i4_3_lut_LC_27_20_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i4_3_lut_LC_27_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i4_3_lut_LC_27_20_2 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \eeprom.rem_4_mux_3_i4_3_lut_LC_27_20_2  (
            .in0(N__25761),
            .in1(N__29172),
            .in2(_gnd_net_),
            .in3(N__25859),
            .lcout(\eeprom.n3722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i31_3_lut_LC_27_20_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i31_3_lut_LC_27_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i31_3_lut_LC_27_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \eeprom.rem_4_mux_3_i31_3_lut_LC_27_20_3  (
            .in0(N__29170),
            .in1(N__25304),
            .in2(_gnd_net_),
            .in3(N__26297),
            .lcout(\eeprom.n1256 ),
            .ltout(\eeprom.n1256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4559_2_lut_LC_27_20_4 .C_ON=1'b0;
    defparam \eeprom.i4559_2_lut_LC_27_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4559_2_lut_LC_27_20_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i4559_2_lut_LC_27_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25571),
            .in3(N__27208),
            .lcout(\eeprom.n1913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_3_lut_LC_27_20_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_3_lut_LC_27_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_3_lut_LC_27_20_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \eeprom.i2c.i1_3_lut_3_lut_LC_27_20_5  (
            .in0(N__27406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27157),
            .lcout(\eeprom.i2c.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_27_20_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_27_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_27_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_27_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25536),
            .lcout(\eeprom.n26_adj_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_27_20_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_27_20_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_27_20_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \eeprom.i2c.i2c_scl_enable_124_LC_27_20_7  (
            .in0(N__27407),
            .in1(N__26892),
            .in2(N__27538),
            .in3(N__27158),
            .lcout(scl_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.i2c_scl_enable_124C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1226_3_lut_LC_27_21_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1226_3_lut_LC_27_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1226_3_lut_LC_27_21_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \eeprom.rem_4_i1226_3_lut_LC_27_21_0  (
            .in0(_gnd_net_),
            .in1(N__27268),
            .in2(N__27254),
            .in3(N__27636),
            .lcout(\eeprom.n1918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_27_21_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_27_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_27_21_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_27_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25489),
            .in3(_gnd_net_),
            .lcout(\eeprom.n33_adj_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1220_3_lut_4_lut_LC_27_21_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1220_3_lut_4_lut_LC_27_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1220_3_lut_4_lut_LC_27_21_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \eeprom.rem_4_i1220_3_lut_4_lut_LC_27_21_2  (
            .in0(N__29169),
            .in1(N__27854),
            .in2(N__28985),
            .in3(N__27637),
            .lcout(\eeprom.n1912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i28_3_lut_LC_27_21_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i28_3_lut_LC_27_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i28_3_lut_LC_27_21_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \eeprom.rem_4_mux_3_i28_3_lut_LC_27_21_3  (
            .in0(N__29168),
            .in1(N__25442),
            .in2(_gnd_net_),
            .in3(N__26357),
            .lcout(\eeprom.n1139 ),
            .ltout(\eeprom.n1139_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1224_3_lut_LC_27_21_4 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1224_3_lut_LC_27_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1224_3_lut_LC_27_21_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \eeprom.rem_4_i1224_3_lut_LC_27_21_4  (
            .in0(N__27230),
            .in1(_gnd_net_),
            .in2(N__25418),
            .in3(N__27635),
            .lcout(\eeprom.n1916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_27_21_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_27_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_27_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_27_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25760),
            .lcout(\eeprom.n30_adj_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_3_lut_LC_27_21_6 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_3_lut_LC_27_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_3_lut_LC_27_21_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \eeprom.i1_2_lut_3_lut_LC_27_21_6  (
            .in0(_gnd_net_),
            .in1(N__27843),
            .in2(N__27209),
            .in3(N__27793),
            .lcout(),
            .ltout(\eeprom.n5035_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_87_LC_27_21_7 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_87_LC_27_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_87_LC_27_21_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_87_LC_27_21_7  (
            .in0(N__27681),
            .in1(N__25722),
            .in2(N__25706),
            .in3(N__27597),
            .lcout(\eeprom.n5039 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_27_22_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_27_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_27_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_27_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25683),
            .lcout(\eeprom.n21_adj_264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_27_22_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_27_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_27_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_27_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29390),
            .lcout(\eeprom.n27_adj_280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_27_22_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_27_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_27_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_27_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25649),
            .lcout(\eeprom.n32_adj_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i26_3_lut_LC_27_22_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i26_3_lut_LC_27_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i26_3_lut_LC_27_22_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \eeprom.rem_4_mux_3_i26_3_lut_LC_27_22_3  (
            .in0(N__29096),
            .in1(_gnd_net_),
            .in2(N__29507),
            .in3(N__26393),
            .lcout(\eeprom.n892 ),
            .ltout(\eeprom.n892_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_42_LC_27_22_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_42_LC_27_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_42_LC_27_22_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_42_LC_27_22_4  (
            .in0(N__29291),
            .in1(N__29098),
            .in2(N__25628),
            .in3(N__26356),
            .lcout(\eeprom.n4977 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_27_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_27_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_27_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_27_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25617),
            .lcout(\eeprom.n23_adj_268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i29_3_lut_LC_27_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i29_3_lut_LC_27_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i29_3_lut_LC_27_22_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \eeprom.rem_4_mux_3_i29_3_lut_LC_27_22_6  (
            .in0(_gnd_net_),
            .in1(N__29097),
            .in2(N__25601),
            .in3(N__26330),
            .lcout(\eeprom.n1138 ),
            .ltout(\eeprom.n1138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4557_1_lut_4_lut_LC_27_22_7 .C_ON=1'b0;
    defparam \eeprom.i4557_1_lut_4_lut_LC_27_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4557_1_lut_4_lut_LC_27_22_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \eeprom.i4557_1_lut_4_lut_LC_27_22_7  (
            .in0(N__27654),
            .in1(N__28981),
            .in2(N__25952),
            .in3(N__27725),
            .lcout(\eeprom.n5327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_27_23_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_27_23_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_27_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_27_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25949),
            .in3(N__25928),
            .lcout(\eeprom.n33 ),
            .ltout(),
            .carryin(bfn_27_23_0_),
            .carryout(\eeprom.n4242 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_27_23_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_27_23_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_27_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_27_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25925),
            .in3(N__25901),
            .lcout(\eeprom.n32_adj_287 ),
            .ltout(),
            .carryin(\eeprom.n4242 ),
            .carryout(\eeprom.n4243 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_27_23_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_27_23_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_27_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_27_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25898),
            .in3(N__25871),
            .lcout(\eeprom.n31_adj_285 ),
            .ltout(),
            .carryin(\eeprom.n4243 ),
            .carryout(\eeprom.n4244 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_27_23_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_27_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_27_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_27_23_3  (
            .in0(_gnd_net_),
            .in1(N__25868),
            .in2(_gnd_net_),
            .in3(N__25850),
            .lcout(\eeprom.n30_adj_284 ),
            .ltout(),
            .carryin(\eeprom.n4244 ),
            .carryout(\eeprom.n4245 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_27_23_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_27_23_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_27_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_27_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25847),
            .in3(N__25820),
            .lcout(\eeprom.n29_adj_283 ),
            .ltout(),
            .carryin(\eeprom.n4245 ),
            .carryout(\eeprom.n4246 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_27_23_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_27_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_27_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_27_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25817),
            .in3(N__25787),
            .lcout(\eeprom.n28_adj_282 ),
            .ltout(),
            .carryin(\eeprom.n4246 ),
            .carryout(\eeprom.n4247 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_27_23_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_27_23_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_27_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_27_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25784),
            .in3(N__25775),
            .lcout(\eeprom.n27_adj_281 ),
            .ltout(),
            .carryin(\eeprom.n4247 ),
            .carryout(\eeprom.n4248 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_27_23_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_27_23_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_27_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_27_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26108),
            .in3(N__26084),
            .lcout(\eeprom.n26_adj_275 ),
            .ltout(),
            .carryin(\eeprom.n4248 ),
            .carryout(\eeprom.n4249 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_27_24_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_27_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_27_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_27_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29222),
            .in3(N__26081),
            .lcout(\eeprom.n25_adj_271 ),
            .ltout(),
            .carryin(bfn_27_24_0_),
            .carryout(\eeprom.n4250 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_27_24_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_27_24_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_27_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_27_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29711),
            .in3(N__26066),
            .lcout(\eeprom.n24_adj_269 ),
            .ltout(),
            .carryin(\eeprom.n4250 ),
            .carryout(\eeprom.n4251 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_27_24_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_27_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_27_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_27_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26063),
            .in3(N__26042),
            .lcout(\eeprom.n23 ),
            .ltout(),
            .carryin(\eeprom.n4251 ),
            .carryout(\eeprom.n4252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_27_24_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_27_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_27_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_27_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29522),
            .in3(N__26027),
            .lcout(\eeprom.n22_adj_265 ),
            .ltout(),
            .carryin(\eeprom.n4252 ),
            .carryout(\eeprom.n4253 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_27_24_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_27_24_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_27_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_27_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26024),
            .in3(N__26000),
            .lcout(\eeprom.n21 ),
            .ltout(),
            .carryin(\eeprom.n4253 ),
            .carryout(\eeprom.n4254 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_27_24_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_27_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_27_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_27_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25997),
            .in3(N__25970),
            .lcout(\eeprom.n20 ),
            .ltout(),
            .carryin(\eeprom.n4254 ),
            .carryout(\eeprom.n4255 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_27_24_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_27_24_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_27_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_27_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27551),
            .in3(N__25955),
            .lcout(\eeprom.n19_adj_320 ),
            .ltout(),
            .carryin(\eeprom.n4255 ),
            .carryout(\eeprom.n4256 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_27_24_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_27_24_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_27_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_27_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29957),
            .in3(N__26270),
            .lcout(\eeprom.n18_adj_326 ),
            .ltout(),
            .carryin(\eeprom.n4256 ),
            .carryout(\eeprom.n4257 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_27_25_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_27_25_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_27_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_27_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26267),
            .in3(N__26249),
            .lcout(\eeprom.n17_adj_324 ),
            .ltout(),
            .carryin(bfn_27_25_0_),
            .carryout(\eeprom.n4258 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_27_25_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_27_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_27_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_27_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26246),
            .in3(N__26228),
            .lcout(\eeprom.n16_adj_325 ),
            .ltout(),
            .carryin(\eeprom.n4258 ),
            .carryout(\eeprom.n4259 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_27_25_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_27_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_27_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_27_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26225),
            .in3(N__26204),
            .lcout(\eeprom.n15 ),
            .ltout(),
            .carryin(\eeprom.n4259 ),
            .carryout(\eeprom.n4260 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_27_25_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_27_25_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_27_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_27_25_3  (
            .in0(_gnd_net_),
            .in1(N__29318),
            .in2(_gnd_net_),
            .in3(N__26192),
            .lcout(\eeprom.n14 ),
            .ltout(),
            .carryin(\eeprom.n4260 ),
            .carryout(\eeprom.n4261 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_27_25_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_27_25_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_27_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_27_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26189),
            .in3(N__26162),
            .lcout(\eeprom.n13_adj_318 ),
            .ltout(),
            .carryin(\eeprom.n4261 ),
            .carryout(\eeprom.n4262 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_27_25_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_27_25_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_27_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_27_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26159),
            .in3(N__26135),
            .lcout(\eeprom.n12_adj_319 ),
            .ltout(),
            .carryin(\eeprom.n4262 ),
            .carryout(\eeprom.n4263 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_27_25_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_27_25_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_27_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_27_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26132),
            .in3(N__26111),
            .lcout(\eeprom.n11 ),
            .ltout(),
            .carryin(\eeprom.n4263 ),
            .carryout(\eeprom.n4264 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_27_25_7 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_27_25_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_27_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_27_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26438),
            .in3(N__26417),
            .lcout(\eeprom.n10_adj_343 ),
            .ltout(),
            .carryin(\eeprom.n4264 ),
            .carryout(\eeprom.n4265 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_27_26_0 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_27_26_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_27_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_27_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26414),
            .in3(N__26396),
            .lcout(\eeprom.n9_adj_308 ),
            .ltout(),
            .carryin(bfn_27_26_0_),
            .carryout(\eeprom.n4266 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_27_26_1 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_27_26_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_27_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_27_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29480),
            .in3(N__26381),
            .lcout(\eeprom.n8_adj_311 ),
            .ltout(),
            .carryin(\eeprom.n4266 ),
            .carryout(\eeprom.n4267 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_27_26_2 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_27_26_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_27_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_27_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26378),
            .in3(N__26369),
            .lcout(\eeprom.n7_adj_309 ),
            .ltout(),
            .carryin(\eeprom.n4267 ),
            .carryout(\eeprom.n4268 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_27_26_3 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_27_26_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_27_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_27_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26366),
            .in3(N__26342),
            .lcout(\eeprom.n6_adj_306 ),
            .ltout(),
            .carryin(\eeprom.n4268 ),
            .carryout(\eeprom.n4269 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_27_26_4 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_27_26_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_27_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_27_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26339),
            .in3(N__26321),
            .lcout(\eeprom.n5_adj_317 ),
            .ltout(),
            .carryin(\eeprom.n4269 ),
            .carryout(\eeprom.n4270 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_27_26_5 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_27_26_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_27_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_27_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26318),
            .in3(N__26309),
            .lcout(\eeprom.n4_adj_310 ),
            .ltout(),
            .carryin(\eeprom.n4270 ),
            .carryout(\eeprom.n4271 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_27_26_6 .C_ON=1'b1;
    defparam \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_27_26_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_27_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_27_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26306),
            .in3(N__26285),
            .lcout(\eeprom.n3_adj_312 ),
            .ltout(),
            .carryin(\eeprom.n4271 ),
            .carryout(\eeprom.n4272 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_27_26_7 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_27_26_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_27_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_27_26_7  (
            .in0(_gnd_net_),
            .in1(N__26659),
            .in2(_gnd_net_),
            .in3(N__26648),
            .lcout(\eeprom.n2_adj_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4695_2_lut_3_lut_4_lut_LC_28_17_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i4695_2_lut_3_lut_4_lut_LC_28_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4695_2_lut_3_lut_4_lut_LC_28_17_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \eeprom.i2c.i4695_2_lut_3_lut_4_lut_LC_28_17_1  (
            .in0(N__27405),
            .in1(N__26853),
            .in2(N__27161),
            .in3(N__27542),
            .lcout(n174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i5_4_lut_LC_28_17_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i5_4_lut_LC_28_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i5_4_lut_LC_28_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2c.i5_4_lut_LC_28_17_5  (
            .in0(N__26641),
            .in1(N__26626),
            .in2(N__26951),
            .in3(N__26614),
            .lcout(),
            .ltout(\eeprom.i2c.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i6_4_lut_LC_28_17_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i6_4_lut_LC_28_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i6_4_lut_LC_28_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2c.i6_4_lut_LC_28_17_6  (
            .in0(N__26602),
            .in1(N__26590),
            .in2(N__26579),
            .in3(N__26550),
            .lcout(\eeprom.i2c.n464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_41_i4_2_lut_LC_28_17_7 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_41_i4_2_lut_LC_28_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_41_i4_2_lut_LC_28_17_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \eeprom.i2c.equal_41_i4_2_lut_LC_28_17_7  (
            .in0(N__27027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26982),
            .lcout(n4_adj_358),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_142_i11_2_lut_3_lut_4_lut_LC_28_18_0 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_142_i11_2_lut_3_lut_4_lut_LC_28_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_142_i11_2_lut_3_lut_4_lut_LC_28_18_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \eeprom.i2c.state_7__I_0_142_i11_2_lut_3_lut_4_lut_LC_28_18_0  (
            .in0(N__27541),
            .in1(N__27402),
            .in2(N__26877),
            .in3(N__27149),
            .lcout(n11_adj_359),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_137_i10_2_lut_LC_28_18_1 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_137_i10_2_lut_LC_28_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_137_i10_2_lut_LC_28_18_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i2c.state_7__I_0_137_i10_2_lut_LC_28_18_1  (
            .in0(_gnd_net_),
            .in1(N__27142),
            .in2(_gnd_net_),
            .in3(N__26839),
            .lcout(n10),
            .ltout(n10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3809_3_lut_4_lut_LC_28_18_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i3809_3_lut_4_lut_LC_28_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3809_3_lut_4_lut_LC_28_18_2 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \eeprom.i2c.i3809_3_lut_4_lut_LC_28_18_2  (
            .in0(N__27539),
            .in1(N__27400),
            .in2(N__26534),
            .in3(N__26493),
            .lcout(\eeprom.i2c.n4579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i2_LC_28_18_3 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i2_LC_28_18_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i2_LC_28_18_3 .LUT_INIT=16'b1111000001110111;
    LogicCell40 \eeprom.i2c.state_i0_i2_LC_28_18_3  (
            .in0(N__27191),
            .in1(N__27185),
            .in2(N__26896),
            .in3(N__27175),
            .lcout(state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29687),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2_2_lut_3_lut_4_lut_LC_28_18_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i2_2_lut_3_lut_4_lut_LC_28_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i2_2_lut_3_lut_4_lut_LC_28_18_4 .LUT_INIT=16'b1111101111111101;
    LogicCell40 \eeprom.i2c.i2_2_lut_3_lut_4_lut_LC_28_18_4  (
            .in0(N__27540),
            .in1(N__27403),
            .in2(N__26878),
            .in3(N__27150),
            .lcout(),
            .ltout(n6_adj_365_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i0_LC_28_18_5 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i0_LC_28_18_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i0_LC_28_18_5 .LUT_INIT=16'b1010101000111111;
    LogicCell40 \eeprom.i2c.state_i0_i0_LC_28_18_5  (
            .in0(N__27404),
            .in1(N__27044),
            .in2(N__27179),
            .in3(N__27174),
            .lcout(state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29687),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3258_2_lut_3_lut_LC_28_18_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i3258_2_lut_3_lut_LC_28_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3258_2_lut_3_lut_LC_28_18_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \eeprom.i2c.i3258_2_lut_3_lut_LC_28_18_6  (
            .in0(N__26840),
            .in1(N__27401),
            .in2(_gnd_net_),
            .in3(N__27148),
            .lcout(n3587),
            .ltout(n3587_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4641_4_lut_LC_28_18_7.C_ON=1'b0;
    defparam i4641_4_lut_LC_28_18_7.SEQ_MODE=4'b0000;
    defparam i4641_4_lut_LC_28_18_7.LUT_INIT=16'b1111000011010000;
    LogicCell40 i4641_4_lut_LC_28_18_7 (
            .in0(N__29798),
            .in1(N__27443),
            .in2(N__27059),
            .in3(N__27056),
            .lcout(n5454),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4645_2_lut_LC_28_19_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i4645_2_lut_LC_28_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4645_2_lut_LC_28_19_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \eeprom.i2c.i4645_2_lut_LC_28_19_0  (
            .in0(_gnd_net_),
            .in1(N__27880),
            .in2(_gnd_net_),
            .in3(N__27036),
            .lcout(),
            .ltout(\eeprom.i2c.n5464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4644_4_lut_LC_28_19_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i4644_4_lut_LC_28_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4644_4_lut_LC_28_19_1 .LUT_INIT=16'b1001100000000000;
    LogicCell40 \eeprom.i2c.i4644_4_lut_LC_28_19_1  (
            .in0(N__26989),
            .in1(N__26950),
            .in2(N__26918),
            .in3(N__27523),
            .lcout(),
            .ltout(\eeprom.i2c.n5451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.sda_out_133_LC_28_19_2 .C_ON=1'b0;
    defparam \eeprom.i2c.sda_out_133_LC_28_19_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.sda_out_133_LC_28_19_2 .LUT_INIT=16'b0001000010111010;
    LogicCell40 \eeprom.i2c.sda_out_133_LC_28_19_2  (
            .in0(N__27437),
            .in1(N__26854),
            .in2(N__26915),
            .in3(N__27408),
            .lcout(\eeprom.i2c.sda_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.sda_out_133C_net ),
            .ce(N__26906),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3210_2_lut_3_lut_LC_28_19_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i3210_2_lut_3_lut_LC_28_19_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3210_2_lut_3_lut_LC_28_19_3 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \eeprom.i2c.i3210_2_lut_3_lut_LC_28_19_3  (
            .in0(N__27410),
            .in1(N__27525),
            .in2(N__26885),
            .in3(_gnd_net_),
            .lcout(n3595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3196_2_lut_LC_28_19_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i3196_2_lut_LC_28_19_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3196_2_lut_LC_28_19_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \eeprom.i2c.i3196_2_lut_LC_28_19_6  (
            .in0(N__27524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27409),
            .lcout(n3581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.write_enable_132_LC_28_20_0 .C_ON=1'b0;
    defparam \eeprom.i2c.write_enable_132_LC_28_20_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.write_enable_132_LC_28_20_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \eeprom.i2c.write_enable_132_LC_28_20_0  (
            .in0(_gnd_net_),
            .in1(N__27436),
            .in2(_gnd_net_),
            .in3(N__27411),
            .lcout(sda_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.write_enable_132C_net ),
            .ce(N__27290),
            .sr(N__27278));
    defparam \eeprom.add_822_2_lut_LC_28_21_0 .C_ON=1'b1;
    defparam \eeprom.add_822_2_lut_LC_28_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_822_2_lut_LC_28_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_822_2_lut_LC_28_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27269),
            .in3(N__27245),
            .lcout(\eeprom.n1198 ),
            .ltout(),
            .carryin(bfn_28_21_0_),
            .carryout(\eeprom.n4273 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_822_3_lut_LC_28_21_1 .C_ON=1'b1;
    defparam \eeprom.add_822_3_lut_LC_28_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_822_3_lut_LC_28_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_822_3_lut_LC_28_21_1  (
            .in0(_gnd_net_),
            .in1(N__28169),
            .in2(N__29273),
            .in3(N__27242),
            .lcout(\eeprom.n1197 ),
            .ltout(),
            .carryin(\eeprom.n4273 ),
            .carryout(\eeprom.n4274 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_822_4_lut_LC_28_21_2 .C_ON=1'b1;
    defparam \eeprom.add_822_4_lut_LC_28_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_822_4_lut_LC_28_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_822_4_lut_LC_28_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27239),
            .in3(N__27224),
            .lcout(\eeprom.n1196 ),
            .ltout(),
            .carryin(\eeprom.n4274 ),
            .carryout(\eeprom.n4275 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_822_5_lut_LC_28_21_3 .C_ON=1'b1;
    defparam \eeprom.add_822_5_lut_LC_28_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_822_5_lut_LC_28_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_822_5_lut_LC_28_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27746),
            .in3(N__27221),
            .lcout(\eeprom.n1195 ),
            .ltout(),
            .carryin(\eeprom.n4275 ),
            .carryout(\eeprom.n4276 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_822_6_lut_LC_28_21_4 .C_ON=1'b1;
    defparam \eeprom.add_822_6_lut_LC_28_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_822_6_lut_LC_28_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_822_6_lut_LC_28_21_4  (
            .in0(_gnd_net_),
            .in1(N__27655),
            .in2(_gnd_net_),
            .in3(N__27218),
            .lcout(\eeprom.n1194 ),
            .ltout(),
            .carryin(\eeprom.n4276 ),
            .carryout(\eeprom.n4277 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_822_7_lut_LC_28_21_5 .C_ON=1'b1;
    defparam \eeprom.add_822_7_lut_LC_28_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_822_7_lut_LC_28_21_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \eeprom.add_822_7_lut_LC_28_21_5  (
            .in0(N__27215),
            .in1(_gnd_net_),
            .in2(N__27844),
            .in3(N__27194),
            .lcout(\eeprom.n5328 ),
            .ltout(),
            .carryin(\eeprom.n4277 ),
            .carryout(\eeprom.n4278 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_822_8_lut_LC_28_21_6 .C_ON=1'b0;
    defparam \eeprom.add_822_8_lut_LC_28_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_822_8_lut_LC_28_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_822_8_lut_LC_28_21_6  (
            .in0(_gnd_net_),
            .in1(N__28946),
            .in2(_gnd_net_),
            .in3(N__27857),
            .lcout(\eeprom.n1192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_2_lut_adj_44_LC_28_22_1 .C_ON=1'b0;
    defparam \eeprom.i1_2_lut_adj_44_LC_28_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_2_lut_adj_44_LC_28_22_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \eeprom.i1_2_lut_adj_44_LC_28_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27845),
            .in3(N__27713),
            .lcout(\eeprom.n1843 ),
            .ltout(\eeprom.n1843_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1223_3_lut_LC_28_22_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1223_3_lut_LC_28_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1223_3_lut_LC_28_22_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_i1223_3_lut_LC_28_22_2  (
            .in0(_gnd_net_),
            .in1(N__27742),
            .in2(N__27818),
            .in3(N__27815),
            .lcout(\eeprom.n1915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i30_3_lut_LC_28_22_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i30_3_lut_LC_28_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i30_3_lut_LC_28_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \eeprom.rem_4_mux_3_i30_3_lut_LC_28_22_3  (
            .in0(N__29185),
            .in1(N__27782),
            .in2(_gnd_net_),
            .in3(N__27758),
            .lcout(\eeprom.n1137 ),
            .ltout(\eeprom.n1137_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_4_lut_adj_43_LC_28_22_4 .C_ON=1'b0;
    defparam \eeprom.i1_4_lut_adj_43_LC_28_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_4_lut_adj_43_LC_28_22_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i1_4_lut_adj_43_LC_28_22_4  (
            .in0(N__28980),
            .in1(N__27741),
            .in2(N__27728),
            .in3(N__27724),
            .lcout(\eeprom.n4983 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_i1225_3_lut_LC_28_22_6 .C_ON=1'b0;
    defparam \eeprom.rem_4_i1225_3_lut_LC_28_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_i1225_3_lut_LC_28_22_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \eeprom.rem_4_i1225_3_lut_LC_28_22_6  (
            .in0(_gnd_net_),
            .in1(N__27707),
            .in2(N__27638),
            .in3(N__29272),
            .lcout(\eeprom.n1917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i4673_3_lut_LC_28_22_7 .C_ON=1'b0;
    defparam \eeprom.i4673_3_lut_LC_28_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i4673_3_lut_LC_28_22_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \eeprom.i4673_3_lut_LC_28_22_7  (
            .in0(_gnd_net_),
            .in1(N__27665),
            .in2(N__27659),
            .in3(N__27631),
            .lcout(\eeprom.n1914 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_28_23_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_28_23_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_28_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_28_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27580),
            .lcout(\eeprom.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i9_3_lut_LC_28_23_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i9_3_lut_LC_28_23_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i9_3_lut_LC_28_23_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \eeprom.rem_4_mux_3_i9_3_lut_LC_28_23_5  (
            .in0(N__29465),
            .in1(N__29205),
            .in2(_gnd_net_),
            .in3(N__29252),
            .lcout(\eeprom.n3519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i7_3_lut_LC_28_24_0 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i7_3_lut_LC_28_24_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i7_3_lut_LC_28_24_0 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \eeprom.rem_4_mux_3_i7_3_lut_LC_28_24_0  (
            .in0(N__29414),
            .in1(N__29137),
            .in2(_gnd_net_),
            .in3(N__29404),
            .lcout(\eeprom.n3719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_28_24_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_28_24_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_28_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_28_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29347),
            .lcout(\eeprom.n14_adj_297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_mux_3_i27_3_lut_LC_28_24_3 .C_ON=1'b0;
    defparam \eeprom.rem_4_mux_3_i27_3_lut_LC_28_24_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_mux_3_i27_3_lut_LC_28_24_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \eeprom.rem_4_mux_3_i27_3_lut_LC_28_24_3  (
            .in0(_gnd_net_),
            .in1(N__29311),
            .in2(N__29184),
            .in3(N__29287),
            .lcout(\eeprom.n1140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_28_24_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_28_24_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_28_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_28_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29251),
            .lcout(\eeprom.n25_adj_272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i401_2_lut_LC_28_25_2 .C_ON=1'b0;
    defparam \eeprom.i401_2_lut_LC_28_25_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i401_2_lut_LC_28_25_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \eeprom.i401_2_lut_LC_28_25_2  (
            .in0(N__29186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28967),
            .lcout(\eeprom.n1135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_29_17_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_29_17_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_29_17_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_29_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.saved_addr__i1_LC_29_17_5 .C_ON=1'b0;
    defparam \eeprom.i2c.saved_addr__i1_LC_29_17_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.saved_addr__i1_LC_29_17_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \eeprom.i2c.saved_addr__i1_LC_29_17_5  (
            .in0(N__29797),
            .in1(N__27908),
            .in2(N__27902),
            .in3(N__27879),
            .lcout(saved_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29658),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.enable_slow_121_LC_29_18_3 .C_ON=1'b0;
    defparam \eeprom.i2c.enable_slow_121_LC_29_18_3 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.enable_slow_121_LC_29_18_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \eeprom.i2c.enable_slow_121_LC_29_18_3  (
            .in0(N__29632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29824),
            .lcout(state_7_N_146_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29862),
            .ce(N__29753),
            .sr(N__29786));
    defparam \eeprom.i2c.i2c_clk_122_LC_29_19_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i2c_clk_122_LC_29_19_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.i2c_clk_122_LC_29_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \eeprom.i2c.i2c_clk_122_LC_29_19_4  (
            .in0(N__29817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29625),
            .lcout(\eeprom.i2c.i2c_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29864),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_29_19_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_29_19_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_29_19_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_LC_29_19_5  (
            .in0(N__29624),
            .in1(N__29781),
            .in2(_gnd_net_),
            .in3(N__29816),
            .lcout(\eeprom.i2c.n1832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_LC_29_20_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_LC_29_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_LC_29_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i1_2_lut_LC_29_20_1  (
            .in0(_gnd_net_),
            .in1(N__29896),
            .in2(_gnd_net_),
            .in3(N__29941),
            .lcout(),
            .ltout(\eeprom.i2c.n6_adj_255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4_4_lut_LC_29_20_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i4_4_lut_LC_29_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4_4_lut_LC_29_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i2c.i4_4_lut_LC_29_20_2  (
            .in0(N__29911),
            .in1(N__29878),
            .in2(N__29741),
            .in3(N__29926),
            .lcout(\eeprom.i2c.counter2_7__N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_29_21_2 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_29_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_29_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_29_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29737),
            .lcout(\eeprom.n24_adj_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i3188_2_lut_LC_29_21_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i3188_2_lut_LC_29_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i3188_2_lut_LC_29_21_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \eeprom.i2c.i3188_2_lut_LC_29_21_5  (
            .in0(N__29657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29578),
            .lcout(scl_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_29_22_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_29_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_29_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_29_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29545),
            .lcout(\eeprom.n22_adj_266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_29_22_5 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_29_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_29_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_29_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29503),
            .lcout(\eeprom.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_29_25_1 .C_ON=1'b0;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_29_25_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_29_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_29_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29983),
            .lcout(\eeprom.n18_adj_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.counter2_229_230__i1_LC_30_20_0 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_229_230__i1_LC_30_20_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_229_230__i1_LC_30_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_229_230__i1_LC_30_20_0  (
            .in0(_gnd_net_),
            .in1(N__29942),
            .in2(_gnd_net_),
            .in3(N__29930),
            .lcout(\eeprom.i2c.counter2_0 ),
            .ltout(),
            .carryin(bfn_30_20_0_),
            .carryout(\eeprom.i2c.n3962 ),
            .clk(N__29867),
            .ce(),
            .sr(N__29825));
    defparam \eeprom.i2c.counter2_229_230__i2_LC_30_20_1 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_229_230__i2_LC_30_20_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_229_230__i2_LC_30_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_229_230__i2_LC_30_20_1  (
            .in0(_gnd_net_),
            .in1(N__29927),
            .in2(_gnd_net_),
            .in3(N__29915),
            .lcout(\eeprom.i2c.counter2_1 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3962 ),
            .carryout(\eeprom.i2c.n3963 ),
            .clk(N__29867),
            .ce(),
            .sr(N__29825));
    defparam \eeprom.i2c.counter2_229_230__i3_LC_30_20_2 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_229_230__i3_LC_30_20_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_229_230__i3_LC_30_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_229_230__i3_LC_30_20_2  (
            .in0(_gnd_net_),
            .in1(N__29912),
            .in2(_gnd_net_),
            .in3(N__29900),
            .lcout(\eeprom.i2c.counter2_2 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3963 ),
            .carryout(\eeprom.i2c.n3964 ),
            .clk(N__29867),
            .ce(),
            .sr(N__29825));
    defparam \eeprom.i2c.counter2_229_230__i4_LC_30_20_3 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_229_230__i4_LC_30_20_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_229_230__i4_LC_30_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_229_230__i4_LC_30_20_3  (
            .in0(_gnd_net_),
            .in1(N__29897),
            .in2(_gnd_net_),
            .in3(N__29885),
            .lcout(\eeprom.i2c.counter2_3 ),
            .ltout(),
            .carryin(\eeprom.i2c.n3964 ),
            .carryout(\eeprom.i2c.n3965 ),
            .clk(N__29867),
            .ce(),
            .sr(N__29825));
    defparam \eeprom.i2c.counter2_229_230__i5_LC_30_20_4 .C_ON=1'b0;
    defparam \eeprom.i2c.counter2_229_230__i5_LC_30_20_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_229_230__i5_LC_30_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_229_230__i5_LC_30_20_4  (
            .in0(_gnd_net_),
            .in1(N__29879),
            .in2(_gnd_net_),
            .in3(N__29882),
            .lcout(\eeprom.i2c.counter2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29867),
            .ce(),
            .sr(N__29825));
endmodule // TinyFPGA_B
