// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Feb 4 2020 22:10:19

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    output USBPU;
    output TX;
    input SDA;
    input SCL;
    input RX;
    output NEOPXL;
    output LED;
    output INLC;
    output INLB;
    output INLA;
    output INHC;
    output INHB;
    output INHA;
    input HALL3;
    input HALL2;
    input HALL1;
    input FAULT_N;
    input ENCODER1_B;
    input ENCODER1_A;
    input ENCODER0_B;
    input ENCODER0_A;
    output DE;
    input CS_MISO;
    output CS_CLK;
    output CS;
    input CLK;

    wire N__56344;
    wire N__56343;
    wire N__56342;
    wire N__56335;
    wire N__56334;
    wire N__56333;
    wire N__56326;
    wire N__56325;
    wire N__56324;
    wire N__56317;
    wire N__56316;
    wire N__56315;
    wire N__56308;
    wire N__56307;
    wire N__56306;
    wire N__56299;
    wire N__56298;
    wire N__56297;
    wire N__56290;
    wire N__56289;
    wire N__56288;
    wire N__56281;
    wire N__56280;
    wire N__56279;
    wire N__56272;
    wire N__56271;
    wire N__56270;
    wire N__56263;
    wire N__56262;
    wire N__56261;
    wire N__56254;
    wire N__56253;
    wire N__56252;
    wire N__56245;
    wire N__56244;
    wire N__56243;
    wire N__56236;
    wire N__56235;
    wire N__56234;
    wire N__56227;
    wire N__56226;
    wire N__56225;
    wire N__56218;
    wire N__56217;
    wire N__56216;
    wire N__56209;
    wire N__56208;
    wire N__56207;
    wire N__56200;
    wire N__56199;
    wire N__56198;
    wire N__56191;
    wire N__56190;
    wire N__56189;
    wire N__56182;
    wire N__56181;
    wire N__56180;
    wire N__56163;
    wire N__56160;
    wire N__56157;
    wire N__56154;
    wire N__56151;
    wire N__56148;
    wire N__56147;
    wire N__56146;
    wire N__56145;
    wire N__56144;
    wire N__56143;
    wire N__56140;
    wire N__56137;
    wire N__56132;
    wire N__56127;
    wire N__56126;
    wire N__56125;
    wire N__56124;
    wire N__56119;
    wire N__56118;
    wire N__56113;
    wire N__56112;
    wire N__56111;
    wire N__56110;
    wire N__56107;
    wire N__56102;
    wire N__56101;
    wire N__56100;
    wire N__56099;
    wire N__56096;
    wire N__56093;
    wire N__56090;
    wire N__56083;
    wire N__56080;
    wire N__56077;
    wire N__56074;
    wire N__56069;
    wire N__56064;
    wire N__56055;
    wire N__56046;
    wire N__56045;
    wire N__56044;
    wire N__56043;
    wire N__56040;
    wire N__56037;
    wire N__56036;
    wire N__56031;
    wire N__56030;
    wire N__56029;
    wire N__56024;
    wire N__56021;
    wire N__56018;
    wire N__56017;
    wire N__56014;
    wire N__56013;
    wire N__56010;
    wire N__56003;
    wire N__56002;
    wire N__55999;
    wire N__55996;
    wire N__55993;
    wire N__55990;
    wire N__55987;
    wire N__55982;
    wire N__55977;
    wire N__55968;
    wire N__55965;
    wire N__55964;
    wire N__55963;
    wire N__55962;
    wire N__55961;
    wire N__55960;
    wire N__55957;
    wire N__55952;
    wire N__55951;
    wire N__55950;
    wire N__55947;
    wire N__55944;
    wire N__55941;
    wire N__55936;
    wire N__55933;
    wire N__55930;
    wire N__55927;
    wire N__55922;
    wire N__55921;
    wire N__55920;
    wire N__55915;
    wire N__55912;
    wire N__55907;
    wire N__55902;
    wire N__55899;
    wire N__55890;
    wire N__55889;
    wire N__55884;
    wire N__55883;
    wire N__55882;
    wire N__55881;
    wire N__55878;
    wire N__55873;
    wire N__55872;
    wire N__55869;
    wire N__55864;
    wire N__55861;
    wire N__55854;
    wire N__55851;
    wire N__55848;
    wire N__55845;
    wire N__55842;
    wire N__55839;
    wire N__55836;
    wire N__55835;
    wire N__55834;
    wire N__55833;
    wire N__55832;
    wire N__55831;
    wire N__55830;
    wire N__55829;
    wire N__55828;
    wire N__55827;
    wire N__55826;
    wire N__55825;
    wire N__55824;
    wire N__55823;
    wire N__55822;
    wire N__55821;
    wire N__55820;
    wire N__55819;
    wire N__55818;
    wire N__55817;
    wire N__55816;
    wire N__55815;
    wire N__55814;
    wire N__55813;
    wire N__55812;
    wire N__55811;
    wire N__55810;
    wire N__55809;
    wire N__55808;
    wire N__55807;
    wire N__55806;
    wire N__55805;
    wire N__55804;
    wire N__55803;
    wire N__55802;
    wire N__55801;
    wire N__55800;
    wire N__55799;
    wire N__55798;
    wire N__55797;
    wire N__55796;
    wire N__55795;
    wire N__55794;
    wire N__55793;
    wire N__55792;
    wire N__55791;
    wire N__55790;
    wire N__55789;
    wire N__55788;
    wire N__55787;
    wire N__55786;
    wire N__55785;
    wire N__55784;
    wire N__55783;
    wire N__55782;
    wire N__55781;
    wire N__55780;
    wire N__55779;
    wire N__55778;
    wire N__55777;
    wire N__55776;
    wire N__55775;
    wire N__55774;
    wire N__55773;
    wire N__55644;
    wire N__55641;
    wire N__55638;
    wire N__55637;
    wire N__55634;
    wire N__55633;
    wire N__55630;
    wire N__55629;
    wire N__55626;
    wire N__55623;
    wire N__55620;
    wire N__55617;
    wire N__55612;
    wire N__55609;
    wire N__55606;
    wire N__55603;
    wire N__55596;
    wire N__55593;
    wire N__55592;
    wire N__55591;
    wire N__55590;
    wire N__55587;
    wire N__55584;
    wire N__55581;
    wire N__55578;
    wire N__55573;
    wire N__55568;
    wire N__55565;
    wire N__55560;
    wire N__55557;
    wire N__55554;
    wire N__55551;
    wire N__55548;
    wire N__55545;
    wire N__55542;
    wire N__55539;
    wire N__55536;
    wire N__55533;
    wire N__55530;
    wire N__55527;
    wire N__55524;
    wire N__55521;
    wire N__55518;
    wire N__55515;
    wire N__55512;
    wire N__55509;
    wire N__55506;
    wire N__55505;
    wire N__55504;
    wire N__55501;
    wire N__55496;
    wire N__55491;
    wire N__55488;
    wire N__55485;
    wire N__55482;
    wire N__55479;
    wire N__55476;
    wire N__55473;
    wire N__55470;
    wire N__55467;
    wire N__55466;
    wire N__55463;
    wire N__55460;
    wire N__55455;
    wire N__55452;
    wire N__55451;
    wire N__55448;
    wire N__55445;
    wire N__55440;
    wire N__55437;
    wire N__55436;
    wire N__55433;
    wire N__55430;
    wire N__55427;
    wire N__55422;
    wire N__55419;
    wire N__55416;
    wire N__55415;
    wire N__55412;
    wire N__55409;
    wire N__55404;
    wire N__55403;
    wire N__55402;
    wire N__55401;
    wire N__55400;
    wire N__55399;
    wire N__55396;
    wire N__55393;
    wire N__55390;
    wire N__55389;
    wire N__55386;
    wire N__55383;
    wire N__55380;
    wire N__55377;
    wire N__55374;
    wire N__55371;
    wire N__55368;
    wire N__55365;
    wire N__55362;
    wire N__55359;
    wire N__55354;
    wire N__55347;
    wire N__55344;
    wire N__55335;
    wire N__55334;
    wire N__55333;
    wire N__55332;
    wire N__55331;
    wire N__55330;
    wire N__55329;
    wire N__55328;
    wire N__55327;
    wire N__55326;
    wire N__55325;
    wire N__55324;
    wire N__55323;
    wire N__55322;
    wire N__55319;
    wire N__55316;
    wire N__55311;
    wire N__55310;
    wire N__55309;
    wire N__55308;
    wire N__55307;
    wire N__55306;
    wire N__55301;
    wire N__55298;
    wire N__55291;
    wire N__55284;
    wire N__55281;
    wire N__55278;
    wire N__55273;
    wire N__55272;
    wire N__55271;
    wire N__55264;
    wire N__55263;
    wire N__55262;
    wire N__55261;
    wire N__55260;
    wire N__55255;
    wire N__55252;
    wire N__55245;
    wire N__55242;
    wire N__55237;
    wire N__55232;
    wire N__55229;
    wire N__55224;
    wire N__55221;
    wire N__55218;
    wire N__55207;
    wire N__55202;
    wire N__55191;
    wire N__55188;
    wire N__55185;
    wire N__55182;
    wire N__55179;
    wire N__55176;
    wire N__55175;
    wire N__55172;
    wire N__55169;
    wire N__55164;
    wire N__55161;
    wire N__55160;
    wire N__55157;
    wire N__55154;
    wire N__55149;
    wire N__55146;
    wire N__55145;
    wire N__55142;
    wire N__55139;
    wire N__55134;
    wire N__55131;
    wire N__55130;
    wire N__55127;
    wire N__55124;
    wire N__55119;
    wire N__55116;
    wire N__55115;
    wire N__55112;
    wire N__55109;
    wire N__55104;
    wire N__55101;
    wire N__55100;
    wire N__55097;
    wire N__55094;
    wire N__55089;
    wire N__55086;
    wire N__55085;
    wire N__55082;
    wire N__55079;
    wire N__55076;
    wire N__55071;
    wire N__55068;
    wire N__55067;
    wire N__55064;
    wire N__55061;
    wire N__55056;
    wire N__55053;
    wire N__55052;
    wire N__55049;
    wire N__55046;
    wire N__55041;
    wire N__55038;
    wire N__55035;
    wire N__55034;
    wire N__55031;
    wire N__55030;
    wire N__55029;
    wire N__55028;
    wire N__55027;
    wire N__55022;
    wire N__55019;
    wire N__55016;
    wire N__55011;
    wire N__55008;
    wire N__54999;
    wire N__54996;
    wire N__54993;
    wire N__54990;
    wire N__54987;
    wire N__54986;
    wire N__54983;
    wire N__54980;
    wire N__54975;
    wire N__54974;
    wire N__54971;
    wire N__54968;
    wire N__54963;
    wire N__54960;
    wire N__54959;
    wire N__54956;
    wire N__54953;
    wire N__54948;
    wire N__54945;
    wire N__54944;
    wire N__54941;
    wire N__54938;
    wire N__54933;
    wire N__54930;
    wire N__54929;
    wire N__54926;
    wire N__54923;
    wire N__54920;
    wire N__54915;
    wire N__54912;
    wire N__54911;
    wire N__54908;
    wire N__54905;
    wire N__54900;
    wire N__54897;
    wire N__54894;
    wire N__54893;
    wire N__54888;
    wire N__54885;
    wire N__54882;
    wire N__54881;
    wire N__54878;
    wire N__54875;
    wire N__54874;
    wire N__54873;
    wire N__54870;
    wire N__54867;
    wire N__54864;
    wire N__54861;
    wire N__54852;
    wire N__54849;
    wire N__54848;
    wire N__54847;
    wire N__54844;
    wire N__54841;
    wire N__54838;
    wire N__54835;
    wire N__54834;
    wire N__54831;
    wire N__54828;
    wire N__54825;
    wire N__54822;
    wire N__54819;
    wire N__54810;
    wire N__54807;
    wire N__54806;
    wire N__54805;
    wire N__54802;
    wire N__54801;
    wire N__54798;
    wire N__54795;
    wire N__54792;
    wire N__54789;
    wire N__54786;
    wire N__54783;
    wire N__54780;
    wire N__54777;
    wire N__54774;
    wire N__54765;
    wire N__54764;
    wire N__54763;
    wire N__54762;
    wire N__54759;
    wire N__54756;
    wire N__54755;
    wire N__54752;
    wire N__54749;
    wire N__54748;
    wire N__54745;
    wire N__54742;
    wire N__54739;
    wire N__54736;
    wire N__54733;
    wire N__54730;
    wire N__54725;
    wire N__54714;
    wire N__54711;
    wire N__54708;
    wire N__54705;
    wire N__54702;
    wire N__54699;
    wire N__54698;
    wire N__54697;
    wire N__54694;
    wire N__54693;
    wire N__54690;
    wire N__54689;
    wire N__54688;
    wire N__54685;
    wire N__54684;
    wire N__54679;
    wire N__54672;
    wire N__54671;
    wire N__54670;
    wire N__54667;
    wire N__54664;
    wire N__54659;
    wire N__54656;
    wire N__54653;
    wire N__54642;
    wire N__54639;
    wire N__54638;
    wire N__54637;
    wire N__54636;
    wire N__54635;
    wire N__54634;
    wire N__54631;
    wire N__54628;
    wire N__54625;
    wire N__54624;
    wire N__54623;
    wire N__54620;
    wire N__54617;
    wire N__54610;
    wire N__54605;
    wire N__54602;
    wire N__54599;
    wire N__54596;
    wire N__54591;
    wire N__54582;
    wire N__54579;
    wire N__54576;
    wire N__54573;
    wire N__54570;
    wire N__54567;
    wire N__54566;
    wire N__54565;
    wire N__54564;
    wire N__54561;
    wire N__54558;
    wire N__54553;
    wire N__54546;
    wire N__54545;
    wire N__54544;
    wire N__54543;
    wire N__54540;
    wire N__54539;
    wire N__54536;
    wire N__54535;
    wire N__54534;
    wire N__54531;
    wire N__54530;
    wire N__54529;
    wire N__54528;
    wire N__54527;
    wire N__54526;
    wire N__54523;
    wire N__54522;
    wire N__54521;
    wire N__54520;
    wire N__54519;
    wire N__54518;
    wire N__54517;
    wire N__54516;
    wire N__54515;
    wire N__54514;
    wire N__54513;
    wire N__54512;
    wire N__54511;
    wire N__54510;
    wire N__54509;
    wire N__54508;
    wire N__54507;
    wire N__54506;
    wire N__54505;
    wire N__54504;
    wire N__54503;
    wire N__54502;
    wire N__54491;
    wire N__54484;
    wire N__54477;
    wire N__54466;
    wire N__54465;
    wire N__54462;
    wire N__54461;
    wire N__54460;
    wire N__54459;
    wire N__54458;
    wire N__54457;
    wire N__54456;
    wire N__54455;
    wire N__54452;
    wire N__54449;
    wire N__54446;
    wire N__54443;
    wire N__54440;
    wire N__54437;
    wire N__54434;
    wire N__54431;
    wire N__54428;
    wire N__54425;
    wire N__54424;
    wire N__54423;
    wire N__54422;
    wire N__54419;
    wire N__54418;
    wire N__54417;
    wire N__54416;
    wire N__54415;
    wire N__54414;
    wire N__54413;
    wire N__54410;
    wire N__54407;
    wire N__54406;
    wire N__54405;
    wire N__54404;
    wire N__54403;
    wire N__54402;
    wire N__54401;
    wire N__54400;
    wire N__54399;
    wire N__54396;
    wire N__54395;
    wire N__54392;
    wire N__54391;
    wire N__54390;
    wire N__54389;
    wire N__54386;
    wire N__54381;
    wire N__54376;
    wire N__54371;
    wire N__54366;
    wire N__54365;
    wire N__54362;
    wire N__54361;
    wire N__54360;
    wire N__54359;
    wire N__54358;
    wire N__54355;
    wire N__54354;
    wire N__54353;
    wire N__54352;
    wire N__54351;
    wire N__54350;
    wire N__54347;
    wire N__54346;
    wire N__54345;
    wire N__54342;
    wire N__54337;
    wire N__54334;
    wire N__54325;
    wire N__54316;
    wire N__54309;
    wire N__54298;
    wire N__54297;
    wire N__54296;
    wire N__54295;
    wire N__54294;
    wire N__54293;
    wire N__54292;
    wire N__54291;
    wire N__54290;
    wire N__54289;
    wire N__54288;
    wire N__54287;
    wire N__54286;
    wire N__54285;
    wire N__54284;
    wire N__54283;
    wire N__54282;
    wire N__54281;
    wire N__54280;
    wire N__54279;
    wire N__54278;
    wire N__54277;
    wire N__54276;
    wire N__54275;
    wire N__54274;
    wire N__54273;
    wire N__54272;
    wire N__54271;
    wire N__54270;
    wire N__54269;
    wire N__54268;
    wire N__54267;
    wire N__54266;
    wire N__54265;
    wire N__54264;
    wire N__54263;
    wire N__54262;
    wire N__54259;
    wire N__54252;
    wire N__54249;
    wire N__54242;
    wire N__54239;
    wire N__54232;
    wire N__54219;
    wire N__54216;
    wire N__54207;
    wire N__54202;
    wire N__54201;
    wire N__54198;
    wire N__54197;
    wire N__54194;
    wire N__54191;
    wire N__54190;
    wire N__54189;
    wire N__54188;
    wire N__54187;
    wire N__54186;
    wire N__54185;
    wire N__54184;
    wire N__54183;
    wire N__54182;
    wire N__54181;
    wire N__54180;
    wire N__54179;
    wire N__54178;
    wire N__54177;
    wire N__54176;
    wire N__54169;
    wire N__54164;
    wire N__54151;
    wire N__54138;
    wire N__54135;
    wire N__54134;
    wire N__54131;
    wire N__54128;
    wire N__54125;
    wire N__54122;
    wire N__54121;
    wire N__54118;
    wire N__54115;
    wire N__54112;
    wire N__54109;
    wire N__54106;
    wire N__54103;
    wire N__54102;
    wire N__54099;
    wire N__54098;
    wire N__54097;
    wire N__54096;
    wire N__54095;
    wire N__54094;
    wire N__54093;
    wire N__54092;
    wire N__54091;
    wire N__54088;
    wire N__54085;
    wire N__54082;
    wire N__54081;
    wire N__54080;
    wire N__54079;
    wire N__54078;
    wire N__54075;
    wire N__54072;
    wire N__54069;
    wire N__54066;
    wire N__54063;
    wire N__54062;
    wire N__54059;
    wire N__54056;
    wire N__54053;
    wire N__54052;
    wire N__54049;
    wire N__54046;
    wire N__54043;
    wire N__54040;
    wire N__54037;
    wire N__54034;
    wire N__54031;
    wire N__54028;
    wire N__54025;
    wire N__54022;
    wire N__54019;
    wire N__54018;
    wire N__54015;
    wire N__54012;
    wire N__54011;
    wire N__54010;
    wire N__54009;
    wire N__54008;
    wire N__54007;
    wire N__54006;
    wire N__54005;
    wire N__54004;
    wire N__54003;
    wire N__54002;
    wire N__54001;
    wire N__54000;
    wire N__53999;
    wire N__53998;
    wire N__53997;
    wire N__53996;
    wire N__53995;
    wire N__53994;
    wire N__53993;
    wire N__53992;
    wire N__53991;
    wire N__53990;
    wire N__53989;
    wire N__53988;
    wire N__53987;
    wire N__53986;
    wire N__53985;
    wire N__53984;
    wire N__53983;
    wire N__53982;
    wire N__53981;
    wire N__53968;
    wire N__53963;
    wire N__53958;
    wire N__53955;
    wire N__53948;
    wire N__53943;
    wire N__53938;
    wire N__53937;
    wire N__53936;
    wire N__53935;
    wire N__53934;
    wire N__53933;
    wire N__53930;
    wire N__53927;
    wire N__53926;
    wire N__53925;
    wire N__53922;
    wire N__53921;
    wire N__53918;
    wire N__53917;
    wire N__53916;
    wire N__53915;
    wire N__53912;
    wire N__53909;
    wire N__53906;
    wire N__53905;
    wire N__53904;
    wire N__53903;
    wire N__53902;
    wire N__53899;
    wire N__53898;
    wire N__53897;
    wire N__53896;
    wire N__53893;
    wire N__53892;
    wire N__53891;
    wire N__53890;
    wire N__53889;
    wire N__53888;
    wire N__53885;
    wire N__53882;
    wire N__53879;
    wire N__53872;
    wire N__53867;
    wire N__53860;
    wire N__53853;
    wire N__53846;
    wire N__53835;
    wire N__53828;
    wire N__53825;
    wire N__53822;
    wire N__53819;
    wire N__53818;
    wire N__53815;
    wire N__53814;
    wire N__53813;
    wire N__53812;
    wire N__53811;
    wire N__53810;
    wire N__53809;
    wire N__53808;
    wire N__53807;
    wire N__53802;
    wire N__53797;
    wire N__53794;
    wire N__53793;
    wire N__53792;
    wire N__53789;
    wire N__53786;
    wire N__53785;
    wire N__53784;
    wire N__53783;
    wire N__53776;
    wire N__53769;
    wire N__53766;
    wire N__53765;
    wire N__53764;
    wire N__53763;
    wire N__53758;
    wire N__53747;
    wire N__53738;
    wire N__53729;
    wire N__53718;
    wire N__53717;
    wire N__53716;
    wire N__53715;
    wire N__53714;
    wire N__53713;
    wire N__53710;
    wire N__53709;
    wire N__53708;
    wire N__53707;
    wire N__53704;
    wire N__53701;
    wire N__53698;
    wire N__53695;
    wire N__53694;
    wire N__53691;
    wire N__53688;
    wire N__53685;
    wire N__53682;
    wire N__53679;
    wire N__53676;
    wire N__53673;
    wire N__53670;
    wire N__53667;
    wire N__53664;
    wire N__53661;
    wire N__53658;
    wire N__53655;
    wire N__53652;
    wire N__53649;
    wire N__53646;
    wire N__53643;
    wire N__53640;
    wire N__53639;
    wire N__53638;
    wire N__53637;
    wire N__53636;
    wire N__53633;
    wire N__53630;
    wire N__53627;
    wire N__53624;
    wire N__53621;
    wire N__53620;
    wire N__53617;
    wire N__53616;
    wire N__53615;
    wire N__53614;
    wire N__53613;
    wire N__53612;
    wire N__53611;
    wire N__53610;
    wire N__53609;
    wire N__53608;
    wire N__53607;
    wire N__53596;
    wire N__53593;
    wire N__53590;
    wire N__53587;
    wire N__53586;
    wire N__53585;
    wire N__53584;
    wire N__53583;
    wire N__53580;
    wire N__53579;
    wire N__53578;
    wire N__53577;
    wire N__53576;
    wire N__53573;
    wire N__53572;
    wire N__53571;
    wire N__53568;
    wire N__53565;
    wire N__53564;
    wire N__53563;
    wire N__53562;
    wire N__53561;
    wire N__53560;
    wire N__53559;
    wire N__53558;
    wire N__53547;
    wire N__53546;
    wire N__53543;
    wire N__53536;
    wire N__53531;
    wire N__53526;
    wire N__53523;
    wire N__53516;
    wire N__53507;
    wire N__53498;
    wire N__53495;
    wire N__53492;
    wire N__53491;
    wire N__53484;
    wire N__53471;
    wire N__53468;
    wire N__53457;
    wire N__53454;
    wire N__53453;
    wire N__53452;
    wire N__53451;
    wire N__53450;
    wire N__53449;
    wire N__53446;
    wire N__53445;
    wire N__53442;
    wire N__53441;
    wire N__53440;
    wire N__53439;
    wire N__53438;
    wire N__53437;
    wire N__53436;
    wire N__53435;
    wire N__53434;
    wire N__53433;
    wire N__53432;
    wire N__53429;
    wire N__53426;
    wire N__53425;
    wire N__53422;
    wire N__53419;
    wire N__53418;
    wire N__53417;
    wire N__53414;
    wire N__53413;
    wire N__53412;
    wire N__53411;
    wire N__53406;
    wire N__53399;
    wire N__53388;
    wire N__53387;
    wire N__53386;
    wire N__53385;
    wire N__53380;
    wire N__53377;
    wire N__53370;
    wire N__53359;
    wire N__53356;
    wire N__53349;
    wire N__53340;
    wire N__53339;
    wire N__53330;
    wire N__53319;
    wire N__53310;
    wire N__53301;
    wire N__53292;
    wire N__53285;
    wire N__53282;
    wire N__53279;
    wire N__53276;
    wire N__53273;
    wire N__53268;
    wire N__53255;
    wire N__53254;
    wire N__53253;
    wire N__53252;
    wire N__53251;
    wire N__53248;
    wire N__53241;
    wire N__53234;
    wire N__53229;
    wire N__53220;
    wire N__53213;
    wire N__53202;
    wire N__53199;
    wire N__53198;
    wire N__53197;
    wire N__53196;
    wire N__53195;
    wire N__53194;
    wire N__53193;
    wire N__53192;
    wire N__53191;
    wire N__53190;
    wire N__53189;
    wire N__53188;
    wire N__53187;
    wire N__53180;
    wire N__53169;
    wire N__53164;
    wire N__53161;
    wire N__53160;
    wire N__53159;
    wire N__53158;
    wire N__53155;
    wire N__53154;
    wire N__53153;
    wire N__53152;
    wire N__53149;
    wire N__53144;
    wire N__53141;
    wire N__53128;
    wire N__53121;
    wire N__53116;
    wire N__53109;
    wire N__53104;
    wire N__53103;
    wire N__53102;
    wire N__53101;
    wire N__53100;
    wire N__53099;
    wire N__53096;
    wire N__53095;
    wire N__53092;
    wire N__53091;
    wire N__53090;
    wire N__53087;
    wire N__53086;
    wire N__53085;
    wire N__53082;
    wire N__53075;
    wire N__53066;
    wire N__53057;
    wire N__53048;
    wire N__53041;
    wire N__53032;
    wire N__53031;
    wire N__53030;
    wire N__53029;
    wire N__53028;
    wire N__53025;
    wire N__53022;
    wire N__53017;
    wire N__53016;
    wire N__53013;
    wire N__53012;
    wire N__53009;
    wire N__53008;
    wire N__53005;
    wire N__53004;
    wire N__53003;
    wire N__53002;
    wire N__53001;
    wire N__53000;
    wire N__52993;
    wire N__52986;
    wire N__52983;
    wire N__52982;
    wire N__52981;
    wire N__52980;
    wire N__52979;
    wire N__52976;
    wire N__52975;
    wire N__52974;
    wire N__52973;
    wire N__52972;
    wire N__52971;
    wire N__52966;
    wire N__52957;
    wire N__52954;
    wire N__52947;
    wire N__52942;
    wire N__52939;
    wire N__52932;
    wire N__52927;
    wire N__52922;
    wire N__52915;
    wire N__52910;
    wire N__52905;
    wire N__52904;
    wire N__52903;
    wire N__52902;
    wire N__52901;
    wire N__52900;
    wire N__52899;
    wire N__52898;
    wire N__52897;
    wire N__52896;
    wire N__52895;
    wire N__52894;
    wire N__52893;
    wire N__52892;
    wire N__52891;
    wire N__52890;
    wire N__52887;
    wire N__52886;
    wire N__52883;
    wire N__52880;
    wire N__52877;
    wire N__52874;
    wire N__52871;
    wire N__52868;
    wire N__52865;
    wire N__52862;
    wire N__52855;
    wire N__52846;
    wire N__52837;
    wire N__52832;
    wire N__52821;
    wire N__52818;
    wire N__52811;
    wire N__52810;
    wire N__52801;
    wire N__52794;
    wire N__52787;
    wire N__52786;
    wire N__52771;
    wire N__52768;
    wire N__52761;
    wire N__52758;
    wire N__52753;
    wire N__52742;
    wire N__52735;
    wire N__52734;
    wire N__52733;
    wire N__52732;
    wire N__52731;
    wire N__52730;
    wire N__52727;
    wire N__52726;
    wire N__52725;
    wire N__52724;
    wire N__52723;
    wire N__52722;
    wire N__52721;
    wire N__52718;
    wire N__52717;
    wire N__52714;
    wire N__52713;
    wire N__52712;
    wire N__52711;
    wire N__52704;
    wire N__52697;
    wire N__52694;
    wire N__52689;
    wire N__52684;
    wire N__52679;
    wire N__52672;
    wire N__52669;
    wire N__52662;
    wire N__52651;
    wire N__52646;
    wire N__52641;
    wire N__52634;
    wire N__52631;
    wire N__52624;
    wire N__52619;
    wire N__52616;
    wire N__52609;
    wire N__52600;
    wire N__52591;
    wire N__52590;
    wire N__52583;
    wire N__52576;
    wire N__52573;
    wire N__52570;
    wire N__52563;
    wire N__52560;
    wire N__52559;
    wire N__52558;
    wire N__52557;
    wire N__52542;
    wire N__52539;
    wire N__52532;
    wire N__52521;
    wire N__52514;
    wire N__52505;
    wire N__52500;
    wire N__52497;
    wire N__52494;
    wire N__52485;
    wire N__52478;
    wire N__52471;
    wire N__52460;
    wire N__52453;
    wire N__52450;
    wire N__52437;
    wire N__52430;
    wire N__52429;
    wire N__52428;
    wire N__52427;
    wire N__52412;
    wire N__52405;
    wire N__52398;
    wire N__52393;
    wire N__52388;
    wire N__52385;
    wire N__52380;
    wire N__52365;
    wire N__52362;
    wire N__52359;
    wire N__52356;
    wire N__52355;
    wire N__52352;
    wire N__52349;
    wire N__52344;
    wire N__52341;
    wire N__52338;
    wire N__52337;
    wire N__52334;
    wire N__52331;
    wire N__52326;
    wire N__52323;
    wire N__52322;
    wire N__52319;
    wire N__52316;
    wire N__52313;
    wire N__52310;
    wire N__52305;
    wire N__52304;
    wire N__52301;
    wire N__52296;
    wire N__52293;
    wire N__52290;
    wire N__52287;
    wire N__52284;
    wire N__52281;
    wire N__52278;
    wire N__52277;
    wire N__52276;
    wire N__52275;
    wire N__52274;
    wire N__52271;
    wire N__52268;
    wire N__52265;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52249;
    wire N__52246;
    wire N__52245;
    wire N__52242;
    wire N__52241;
    wire N__52240;
    wire N__52239;
    wire N__52236;
    wire N__52233;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52221;
    wire N__52218;
    wire N__52215;
    wire N__52200;
    wire N__52197;
    wire N__52196;
    wire N__52195;
    wire N__52192;
    wire N__52189;
    wire N__52186;
    wire N__52183;
    wire N__52180;
    wire N__52177;
    wire N__52170;
    wire N__52167;
    wire N__52164;
    wire N__52161;
    wire N__52158;
    wire N__52155;
    wire N__52152;
    wire N__52149;
    wire N__52146;
    wire N__52143;
    wire N__52140;
    wire N__52137;
    wire N__52136;
    wire N__52133;
    wire N__52130;
    wire N__52125;
    wire N__52122;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52109;
    wire N__52108;
    wire N__52107;
    wire N__52106;
    wire N__52103;
    wire N__52100;
    wire N__52099;
    wire N__52096;
    wire N__52095;
    wire N__52092;
    wire N__52091;
    wire N__52088;
    wire N__52087;
    wire N__52086;
    wire N__52085;
    wire N__52084;
    wire N__52083;
    wire N__52082;
    wire N__52081;
    wire N__52078;
    wire N__52061;
    wire N__52058;
    wire N__52057;
    wire N__52054;
    wire N__52053;
    wire N__52050;
    wire N__52049;
    wire N__52046;
    wire N__52045;
    wire N__52044;
    wire N__52043;
    wire N__52042;
    wire N__52039;
    wire N__52038;
    wire N__52037;
    wire N__52036;
    wire N__52035;
    wire N__52034;
    wire N__52033;
    wire N__52030;
    wire N__52025;
    wire N__52008;
    wire N__51999;
    wire N__51990;
    wire N__51985;
    wire N__51972;
    wire N__51969;
    wire N__51966;
    wire N__51963;
    wire N__51960;
    wire N__51957;
    wire N__51954;
    wire N__51953;
    wire N__51950;
    wire N__51947;
    wire N__51944;
    wire N__51939;
    wire N__51936;
    wire N__51933;
    wire N__51930;
    wire N__51927;
    wire N__51924;
    wire N__51921;
    wire N__51920;
    wire N__51917;
    wire N__51914;
    wire N__51913;
    wire N__51910;
    wire N__51907;
    wire N__51904;
    wire N__51901;
    wire N__51894;
    wire N__51891;
    wire N__51888;
    wire N__51885;
    wire N__51882;
    wire N__51881;
    wire N__51878;
    wire N__51875;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51865;
    wire N__51860;
    wire N__51857;
    wire N__51852;
    wire N__51849;
    wire N__51846;
    wire N__51843;
    wire N__51842;
    wire N__51839;
    wire N__51836;
    wire N__51833;
    wire N__51830;
    wire N__51825;
    wire N__51824;
    wire N__51821;
    wire N__51818;
    wire N__51813;
    wire N__51810;
    wire N__51807;
    wire N__51804;
    wire N__51803;
    wire N__51800;
    wire N__51797;
    wire N__51794;
    wire N__51791;
    wire N__51788;
    wire N__51787;
    wire N__51784;
    wire N__51781;
    wire N__51778;
    wire N__51771;
    wire N__51768;
    wire N__51765;
    wire N__51762;
    wire N__51761;
    wire N__51758;
    wire N__51755;
    wire N__51752;
    wire N__51749;
    wire N__51748;
    wire N__51745;
    wire N__51742;
    wire N__51739;
    wire N__51732;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51720;
    wire N__51719;
    wire N__51716;
    wire N__51713;
    wire N__51710;
    wire N__51707;
    wire N__51704;
    wire N__51699;
    wire N__51696;
    wire N__51693;
    wire N__51690;
    wire N__51687;
    wire N__51684;
    wire N__51683;
    wire N__51682;
    wire N__51679;
    wire N__51674;
    wire N__51669;
    wire N__51668;
    wire N__51665;
    wire N__51662;
    wire N__51659;
    wire N__51654;
    wire N__51651;
    wire N__51648;
    wire N__51645;
    wire N__51642;
    wire N__51639;
    wire N__51638;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51628;
    wire N__51625;
    wire N__51622;
    wire N__51619;
    wire N__51616;
    wire N__51609;
    wire N__51606;
    wire N__51603;
    wire N__51602;
    wire N__51601;
    wire N__51598;
    wire N__51597;
    wire N__51594;
    wire N__51591;
    wire N__51590;
    wire N__51589;
    wire N__51586;
    wire N__51583;
    wire N__51582;
    wire N__51581;
    wire N__51576;
    wire N__51573;
    wire N__51570;
    wire N__51569;
    wire N__51568;
    wire N__51567;
    wire N__51564;
    wire N__51557;
    wire N__51552;
    wire N__51547;
    wire N__51542;
    wire N__51531;
    wire N__51528;
    wire N__51525;
    wire N__51522;
    wire N__51521;
    wire N__51518;
    wire N__51515;
    wire N__51510;
    wire N__51507;
    wire N__51506;
    wire N__51505;
    wire N__51502;
    wire N__51497;
    wire N__51494;
    wire N__51489;
    wire N__51488;
    wire N__51487;
    wire N__51484;
    wire N__51481;
    wire N__51478;
    wire N__51475;
    wire N__51468;
    wire N__51465;
    wire N__51464;
    wire N__51463;
    wire N__51460;
    wire N__51455;
    wire N__51452;
    wire N__51449;
    wire N__51446;
    wire N__51441;
    wire N__51438;
    wire N__51435;
    wire N__51432;
    wire N__51429;
    wire N__51428;
    wire N__51425;
    wire N__51422;
    wire N__51419;
    wire N__51416;
    wire N__51413;
    wire N__51410;
    wire N__51405;
    wire N__51402;
    wire N__51401;
    wire N__51400;
    wire N__51399;
    wire N__51398;
    wire N__51397;
    wire N__51394;
    wire N__51393;
    wire N__51392;
    wire N__51391;
    wire N__51388;
    wire N__51387;
    wire N__51386;
    wire N__51383;
    wire N__51380;
    wire N__51379;
    wire N__51376;
    wire N__51375;
    wire N__51372;
    wire N__51369;
    wire N__51366;
    wire N__51363;
    wire N__51358;
    wire N__51351;
    wire N__51342;
    wire N__51339;
    wire N__51324;
    wire N__51321;
    wire N__51318;
    wire N__51317;
    wire N__51314;
    wire N__51311;
    wire N__51306;
    wire N__51303;
    wire N__51300;
    wire N__51297;
    wire N__51296;
    wire N__51295;
    wire N__51294;
    wire N__51291;
    wire N__51288;
    wire N__51287;
    wire N__51284;
    wire N__51283;
    wire N__51282;
    wire N__51281;
    wire N__51278;
    wire N__51277;
    wire N__51274;
    wire N__51271;
    wire N__51270;
    wire N__51267;
    wire N__51266;
    wire N__51261;
    wire N__51258;
    wire N__51255;
    wire N__51252;
    wire N__51249;
    wire N__51248;
    wire N__51243;
    wire N__51236;
    wire N__51227;
    wire N__51222;
    wire N__51213;
    wire N__51212;
    wire N__51211;
    wire N__51208;
    wire N__51205;
    wire N__51202;
    wire N__51199;
    wire N__51194;
    wire N__51189;
    wire N__51186;
    wire N__51183;
    wire N__51180;
    wire N__51177;
    wire N__51174;
    wire N__51171;
    wire N__51168;
    wire N__51167;
    wire N__51166;
    wire N__51161;
    wire N__51158;
    wire N__51153;
    wire N__51150;
    wire N__51147;
    wire N__51144;
    wire N__51141;
    wire N__51138;
    wire N__51137;
    wire N__51134;
    wire N__51131;
    wire N__51128;
    wire N__51125;
    wire N__51120;
    wire N__51119;
    wire N__51118;
    wire N__51115;
    wire N__51112;
    wire N__51109;
    wire N__51102;
    wire N__51099;
    wire N__51098;
    wire N__51095;
    wire N__51092;
    wire N__51091;
    wire N__51088;
    wire N__51085;
    wire N__51082;
    wire N__51075;
    wire N__51072;
    wire N__51069;
    wire N__51066;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51056;
    wire N__51055;
    wire N__51052;
    wire N__51049;
    wire N__51046;
    wire N__51043;
    wire N__51036;
    wire N__51033;
    wire N__51030;
    wire N__51027;
    wire N__51024;
    wire N__51021;
    wire N__51020;
    wire N__51017;
    wire N__51016;
    wire N__51013;
    wire N__51010;
    wire N__51007;
    wire N__51004;
    wire N__51001;
    wire N__50994;
    wire N__50991;
    wire N__50988;
    wire N__50985;
    wire N__50982;
    wire N__50979;
    wire N__50978;
    wire N__50975;
    wire N__50972;
    wire N__50969;
    wire N__50966;
    wire N__50961;
    wire N__50958;
    wire N__50955;
    wire N__50952;
    wire N__50949;
    wire N__50948;
    wire N__50947;
    wire N__50944;
    wire N__50939;
    wire N__50934;
    wire N__50931;
    wire N__50928;
    wire N__50925;
    wire N__50922;
    wire N__50921;
    wire N__50920;
    wire N__50917;
    wire N__50912;
    wire N__50907;
    wire N__50904;
    wire N__50901;
    wire N__50898;
    wire N__50895;
    wire N__50892;
    wire N__50889;
    wire N__50886;
    wire N__50883;
    wire N__50880;
    wire N__50879;
    wire N__50876;
    wire N__50875;
    wire N__50872;
    wire N__50869;
    wire N__50866;
    wire N__50859;
    wire N__50856;
    wire N__50853;
    wire N__50850;
    wire N__50847;
    wire N__50844;
    wire N__50841;
    wire N__50840;
    wire N__50837;
    wire N__50834;
    wire N__50831;
    wire N__50828;
    wire N__50823;
    wire N__50820;
    wire N__50817;
    wire N__50814;
    wire N__50813;
    wire N__50810;
    wire N__50807;
    wire N__50802;
    wire N__50799;
    wire N__50798;
    wire N__50795;
    wire N__50792;
    wire N__50789;
    wire N__50786;
    wire N__50781;
    wire N__50778;
    wire N__50775;
    wire N__50772;
    wire N__50769;
    wire N__50766;
    wire N__50765;
    wire N__50764;
    wire N__50761;
    wire N__50756;
    wire N__50751;
    wire N__50748;
    wire N__50747;
    wire N__50746;
    wire N__50743;
    wire N__50740;
    wire N__50737;
    wire N__50734;
    wire N__50727;
    wire N__50724;
    wire N__50721;
    wire N__50718;
    wire N__50715;
    wire N__50712;
    wire N__50711;
    wire N__50708;
    wire N__50705;
    wire N__50704;
    wire N__50701;
    wire N__50698;
    wire N__50695;
    wire N__50688;
    wire N__50685;
    wire N__50682;
    wire N__50679;
    wire N__50676;
    wire N__50673;
    wire N__50672;
    wire N__50669;
    wire N__50668;
    wire N__50667;
    wire N__50666;
    wire N__50663;
    wire N__50662;
    wire N__50661;
    wire N__50658;
    wire N__50655;
    wire N__50654;
    wire N__50653;
    wire N__50652;
    wire N__50649;
    wire N__50648;
    wire N__50647;
    wire N__50646;
    wire N__50643;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50633;
    wire N__50632;
    wire N__50629;
    wire N__50626;
    wire N__50623;
    wire N__50618;
    wire N__50607;
    wire N__50604;
    wire N__50595;
    wire N__50580;
    wire N__50577;
    wire N__50576;
    wire N__50575;
    wire N__50572;
    wire N__50569;
    wire N__50566;
    wire N__50563;
    wire N__50556;
    wire N__50555;
    wire N__50554;
    wire N__50551;
    wire N__50548;
    wire N__50545;
    wire N__50542;
    wire N__50539;
    wire N__50536;
    wire N__50529;
    wire N__50528;
    wire N__50525;
    wire N__50522;
    wire N__50521;
    wire N__50516;
    wire N__50513;
    wire N__50510;
    wire N__50507;
    wire N__50502;
    wire N__50499;
    wire N__50496;
    wire N__50493;
    wire N__50490;
    wire N__50489;
    wire N__50486;
    wire N__50483;
    wire N__50480;
    wire N__50477;
    wire N__50472;
    wire N__50469;
    wire N__50466;
    wire N__50463;
    wire N__50460;
    wire N__50457;
    wire N__50454;
    wire N__50453;
    wire N__50450;
    wire N__50447;
    wire N__50444;
    wire N__50443;
    wire N__50440;
    wire N__50437;
    wire N__50434;
    wire N__50427;
    wire N__50424;
    wire N__50421;
    wire N__50418;
    wire N__50415;
    wire N__50414;
    wire N__50411;
    wire N__50410;
    wire N__50407;
    wire N__50404;
    wire N__50401;
    wire N__50394;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50384;
    wire N__50381;
    wire N__50378;
    wire N__50375;
    wire N__50372;
    wire N__50371;
    wire N__50366;
    wire N__50363;
    wire N__50360;
    wire N__50355;
    wire N__50352;
    wire N__50349;
    wire N__50346;
    wire N__50343;
    wire N__50340;
    wire N__50339;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50313;
    wire N__50312;
    wire N__50309;
    wire N__50306;
    wire N__50303;
    wire N__50300;
    wire N__50299;
    wire N__50294;
    wire N__50291;
    wire N__50286;
    wire N__50285;
    wire N__50282;
    wire N__50279;
    wire N__50276;
    wire N__50273;
    wire N__50268;
    wire N__50267;
    wire N__50264;
    wire N__50261;
    wire N__50256;
    wire N__50253;
    wire N__50250;
    wire N__50249;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50223;
    wire N__50220;
    wire N__50217;
    wire N__50214;
    wire N__50211;
    wire N__50208;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50196;
    wire N__50195;
    wire N__50192;
    wire N__50189;
    wire N__50188;
    wire N__50187;
    wire N__50186;
    wire N__50183;
    wire N__50176;
    wire N__50175;
    wire N__50172;
    wire N__50171;
    wire N__50170;
    wire N__50169;
    wire N__50168;
    wire N__50167;
    wire N__50166;
    wire N__50165;
    wire N__50160;
    wire N__50153;
    wire N__50150;
    wire N__50147;
    wire N__50146;
    wire N__50145;
    wire N__50144;
    wire N__50137;
    wire N__50134;
    wire N__50129;
    wire N__50118;
    wire N__50109;
    wire N__50106;
    wire N__50105;
    wire N__50102;
    wire N__50099;
    wire N__50096;
    wire N__50093;
    wire N__50092;
    wire N__50087;
    wire N__50084;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50070;
    wire N__50067;
    wire N__50064;
    wire N__50061;
    wire N__50058;
    wire N__50055;
    wire N__50052;
    wire N__50051;
    wire N__50048;
    wire N__50045;
    wire N__50042;
    wire N__50039;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50022;
    wire N__50019;
    wire N__50016;
    wire N__50013;
    wire N__50012;
    wire N__50009;
    wire N__50006;
    wire N__50005;
    wire N__50000;
    wire N__49997;
    wire N__49992;
    wire N__49991;
    wire N__49988;
    wire N__49987;
    wire N__49984;
    wire N__49981;
    wire N__49978;
    wire N__49977;
    wire N__49974;
    wire N__49971;
    wire N__49968;
    wire N__49965;
    wire N__49956;
    wire N__49955;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49943;
    wire N__49940;
    wire N__49937;
    wire N__49934;
    wire N__49929;
    wire N__49928;
    wire N__49925;
    wire N__49922;
    wire N__49919;
    wire N__49914;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49908;
    wire N__49907;
    wire N__49904;
    wire N__49903;
    wire N__49900;
    wire N__49899;
    wire N__49896;
    wire N__49881;
    wire N__49878;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49866;
    wire N__49863;
    wire N__49862;
    wire N__49861;
    wire N__49858;
    wire N__49853;
    wire N__49848;
    wire N__49845;
    wire N__49842;
    wire N__49841;
    wire N__49840;
    wire N__49837;
    wire N__49834;
    wire N__49831;
    wire N__49824;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49800;
    wire N__49797;
    wire N__49794;
    wire N__49791;
    wire N__49790;
    wire N__49787;
    wire N__49784;
    wire N__49781;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49763;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49753;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49736;
    wire N__49735;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49713;
    wire N__49710;
    wire N__49707;
    wire N__49704;
    wire N__49703;
    wire N__49700;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49687;
    wire N__49682;
    wire N__49677;
    wire N__49674;
    wire N__49671;
    wire N__49668;
    wire N__49667;
    wire N__49666;
    wire N__49663;
    wire N__49658;
    wire N__49653;
    wire N__49650;
    wire N__49647;
    wire N__49644;
    wire N__49643;
    wire N__49640;
    wire N__49639;
    wire N__49636;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49620;
    wire N__49617;
    wire N__49614;
    wire N__49611;
    wire N__49610;
    wire N__49609;
    wire N__49606;
    wire N__49603;
    wire N__49600;
    wire N__49593;
    wire N__49590;
    wire N__49589;
    wire N__49586;
    wire N__49585;
    wire N__49582;
    wire N__49581;
    wire N__49578;
    wire N__49575;
    wire N__49572;
    wire N__49569;
    wire N__49566;
    wire N__49561;
    wire N__49554;
    wire N__49551;
    wire N__49548;
    wire N__49547;
    wire N__49544;
    wire N__49541;
    wire N__49538;
    wire N__49537;
    wire N__49534;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49521;
    wire N__49516;
    wire N__49513;
    wire N__49506;
    wire N__49503;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49485;
    wire N__49484;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49458;
    wire N__49455;
    wire N__49446;
    wire N__49443;
    wire N__49442;
    wire N__49439;
    wire N__49436;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49426;
    wire N__49425;
    wire N__49422;
    wire N__49419;
    wire N__49416;
    wire N__49413;
    wire N__49410;
    wire N__49407;
    wire N__49404;
    wire N__49395;
    wire N__49392;
    wire N__49389;
    wire N__49388;
    wire N__49387;
    wire N__49384;
    wire N__49381;
    wire N__49380;
    wire N__49377;
    wire N__49374;
    wire N__49371;
    wire N__49368;
    wire N__49365;
    wire N__49362;
    wire N__49359;
    wire N__49356;
    wire N__49347;
    wire N__49344;
    wire N__49341;
    wire N__49340;
    wire N__49337;
    wire N__49334;
    wire N__49333;
    wire N__49332;
    wire N__49329;
    wire N__49326;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49302;
    wire N__49299;
    wire N__49296;
    wire N__49293;
    wire N__49290;
    wire N__49289;
    wire N__49288;
    wire N__49285;
    wire N__49282;
    wire N__49281;
    wire N__49278;
    wire N__49275;
    wire N__49272;
    wire N__49269;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49253;
    wire N__49250;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49230;
    wire N__49227;
    wire N__49218;
    wire N__49215;
    wire N__49212;
    wire N__49211;
    wire N__49208;
    wire N__49207;
    wire N__49204;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49194;
    wire N__49191;
    wire N__49186;
    wire N__49183;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49166;
    wire N__49163;
    wire N__49160;
    wire N__49157;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49140;
    wire N__49137;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49114;
    wire N__49107;
    wire N__49104;
    wire N__49101;
    wire N__49100;
    wire N__49097;
    wire N__49094;
    wire N__49091;
    wire N__49090;
    wire N__49089;
    wire N__49086;
    wire N__49083;
    wire N__49078;
    wire N__49071;
    wire N__49068;
    wire N__49067;
    wire N__49064;
    wire N__49061;
    wire N__49058;
    wire N__49057;
    wire N__49056;
    wire N__49053;
    wire N__49050;
    wire N__49047;
    wire N__49044;
    wire N__49039;
    wire N__49036;
    wire N__49033;
    wire N__49030;
    wire N__49023;
    wire N__49020;
    wire N__49019;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49009;
    wire N__49008;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48987;
    wire N__48984;
    wire N__48981;
    wire N__48978;
    wire N__48977;
    wire N__48976;
    wire N__48973;
    wire N__48972;
    wire N__48969;
    wire N__48966;
    wire N__48963;
    wire N__48960;
    wire N__48957;
    wire N__48948;
    wire N__48945;
    wire N__48942;
    wire N__48941;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48931;
    wire N__48928;
    wire N__48927;
    wire N__48924;
    wire N__48921;
    wire N__48918;
    wire N__48915;
    wire N__48910;
    wire N__48903;
    wire N__48900;
    wire N__48897;
    wire N__48896;
    wire N__48893;
    wire N__48890;
    wire N__48889;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48879;
    wire N__48876;
    wire N__48871;
    wire N__48864;
    wire N__48861;
    wire N__48858;
    wire N__48855;
    wire N__48852;
    wire N__48849;
    wire N__48846;
    wire N__48843;
    wire N__48840;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48828;
    wire N__48825;
    wire N__48822;
    wire N__48819;
    wire N__48816;
    wire N__48815;
    wire N__48812;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48795;
    wire N__48792;
    wire N__48789;
    wire N__48788;
    wire N__48785;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48775;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48759;
    wire N__48756;
    wire N__48755;
    wire N__48752;
    wire N__48749;
    wire N__48746;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48729;
    wire N__48726;
    wire N__48725;
    wire N__48722;
    wire N__48721;
    wire N__48718;
    wire N__48715;
    wire N__48712;
    wire N__48705;
    wire N__48704;
    wire N__48703;
    wire N__48700;
    wire N__48695;
    wire N__48692;
    wire N__48687;
    wire N__48686;
    wire N__48685;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48669;
    wire N__48666;
    wire N__48663;
    wire N__48660;
    wire N__48659;
    wire N__48656;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48639;
    wire N__48636;
    wire N__48633;
    wire N__48630;
    wire N__48627;
    wire N__48624;
    wire N__48623;
    wire N__48620;
    wire N__48617;
    wire N__48614;
    wire N__48611;
    wire N__48606;
    wire N__48603;
    wire N__48600;
    wire N__48597;
    wire N__48594;
    wire N__48591;
    wire N__48588;
    wire N__48585;
    wire N__48582;
    wire N__48579;
    wire N__48576;
    wire N__48573;
    wire N__48570;
    wire N__48567;
    wire N__48564;
    wire N__48561;
    wire N__48558;
    wire N__48555;
    wire N__48552;
    wire N__48549;
    wire N__48546;
    wire N__48543;
    wire N__48540;
    wire N__48537;
    wire N__48534;
    wire N__48533;
    wire N__48530;
    wire N__48527;
    wire N__48522;
    wire N__48519;
    wire N__48516;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48506;
    wire N__48503;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48482;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48444;
    wire N__48441;
    wire N__48440;
    wire N__48437;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48420;
    wire N__48417;
    wire N__48416;
    wire N__48413;
    wire N__48410;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48393;
    wire N__48392;
    wire N__48391;
    wire N__48388;
    wire N__48383;
    wire N__48380;
    wire N__48375;
    wire N__48372;
    wire N__48369;
    wire N__48366;
    wire N__48363;
    wire N__48360;
    wire N__48357;
    wire N__48354;
    wire N__48351;
    wire N__48348;
    wire N__48345;
    wire N__48342;
    wire N__48341;
    wire N__48338;
    wire N__48335;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48315;
    wire N__48312;
    wire N__48309;
    wire N__48306;
    wire N__48305;
    wire N__48304;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48285;
    wire N__48282;
    wire N__48279;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48264;
    wire N__48263;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48253;
    wire N__48246;
    wire N__48243;
    wire N__48240;
    wire N__48237;
    wire N__48234;
    wire N__48231;
    wire N__48228;
    wire N__48225;
    wire N__48224;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48214;
    wire N__48211;
    wire N__48208;
    wire N__48205;
    wire N__48200;
    wire N__48197;
    wire N__48192;
    wire N__48189;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48181;
    wire N__48178;
    wire N__48173;
    wire N__48168;
    wire N__48167;
    wire N__48164;
    wire N__48161;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48132;
    wire N__48129;
    wire N__48126;
    wire N__48125;
    wire N__48122;
    wire N__48119;
    wire N__48116;
    wire N__48113;
    wire N__48112;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48097;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48072;
    wire N__48071;
    wire N__48070;
    wire N__48067;
    wire N__48064;
    wire N__48061;
    wire N__48058;
    wire N__48055;
    wire N__48052;
    wire N__48045;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48033;
    wire N__48030;
    wire N__48027;
    wire N__48026;
    wire N__48023;
    wire N__48022;
    wire N__48019;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48003;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47982;
    wire N__47981;
    wire N__47978;
    wire N__47975;
    wire N__47970;
    wire N__47967;
    wire N__47964;
    wire N__47963;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47946;
    wire N__47943;
    wire N__47942;
    wire N__47939;
    wire N__47936;
    wire N__47933;
    wire N__47930;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47910;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47900;
    wire N__47895;
    wire N__47892;
    wire N__47891;
    wire N__47888;
    wire N__47885;
    wire N__47884;
    wire N__47881;
    wire N__47876;
    wire N__47871;
    wire N__47868;
    wire N__47865;
    wire N__47862;
    wire N__47861;
    wire N__47858;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47841;
    wire N__47838;
    wire N__47835;
    wire N__47832;
    wire N__47829;
    wire N__47828;
    wire N__47825;
    wire N__47822;
    wire N__47817;
    wire N__47814;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47790;
    wire N__47787;
    wire N__47786;
    wire N__47785;
    wire N__47780;
    wire N__47777;
    wire N__47774;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47745;
    wire N__47744;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47734;
    wire N__47727;
    wire N__47724;
    wire N__47723;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47713;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47691;
    wire N__47690;
    wire N__47689;
    wire N__47686;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47676;
    wire N__47673;
    wire N__47672;
    wire N__47663;
    wire N__47662;
    wire N__47659;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47640;
    wire N__47637;
    wire N__47636;
    wire N__47635;
    wire N__47634;
    wire N__47633;
    wire N__47630;
    wire N__47627;
    wire N__47622;
    wire N__47621;
    wire N__47618;
    wire N__47611;
    wire N__47608;
    wire N__47603;
    wire N__47598;
    wire N__47597;
    wire N__47596;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47586;
    wire N__47585;
    wire N__47582;
    wire N__47581;
    wire N__47578;
    wire N__47575;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47559;
    wire N__47556;
    wire N__47553;
    wire N__47544;
    wire N__47543;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47519;
    wire N__47516;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47474;
    wire N__47469;
    wire N__47468;
    wire N__47465;
    wire N__47462;
    wire N__47459;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47435;
    wire N__47432;
    wire N__47429;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47417;
    wire N__47414;
    wire N__47411;
    wire N__47408;
    wire N__47403;
    wire N__47400;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47367;
    wire N__47364;
    wire N__47361;
    wire N__47358;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47346;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47325;
    wire N__47322;
    wire N__47319;
    wire N__47310;
    wire N__47307;
    wire N__47306;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47296;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47282;
    wire N__47277;
    wire N__47276;
    wire N__47273;
    wire N__47270;
    wire N__47269;
    wire N__47268;
    wire N__47263;
    wire N__47260;
    wire N__47257;
    wire N__47254;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47242;
    wire N__47239;
    wire N__47236;
    wire N__47229;
    wire N__47228;
    wire N__47225;
    wire N__47222;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47210;
    wire N__47207;
    wire N__47204;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47189;
    wire N__47188;
    wire N__47183;
    wire N__47180;
    wire N__47179;
    wire N__47178;
    wire N__47173;
    wire N__47170;
    wire N__47167;
    wire N__47164;
    wire N__47157;
    wire N__47156;
    wire N__47155;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47136;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47124;
    wire N__47121;
    wire N__47118;
    wire N__47115;
    wire N__47112;
    wire N__47111;
    wire N__47110;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47088;
    wire N__47087;
    wire N__47086;
    wire N__47083;
    wire N__47080;
    wire N__47077;
    wire N__47074;
    wire N__47067;
    wire N__47064;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47051;
    wire N__47048;
    wire N__47045;
    wire N__47040;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47028;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47013;
    wire N__47012;
    wire N__47009;
    wire N__47006;
    wire N__47001;
    wire N__47000;
    wire N__46997;
    wire N__46994;
    wire N__46989;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46977;
    wire N__46974;
    wire N__46973;
    wire N__46970;
    wire N__46967;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46953;
    wire N__46952;
    wire N__46951;
    wire N__46948;
    wire N__46945;
    wire N__46942;
    wire N__46935;
    wire N__46932;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46914;
    wire N__46911;
    wire N__46908;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46889;
    wire N__46886;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46869;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46841;
    wire N__46838;
    wire N__46835;
    wire N__46832;
    wire N__46827;
    wire N__46826;
    wire N__46823;
    wire N__46820;
    wire N__46817;
    wire N__46812;
    wire N__46811;
    wire N__46808;
    wire N__46805;
    wire N__46802;
    wire N__46797;
    wire N__46794;
    wire N__46793;
    wire N__46790;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46780;
    wire N__46773;
    wire N__46772;
    wire N__46771;
    wire N__46768;
    wire N__46765;
    wire N__46762;
    wire N__46759;
    wire N__46752;
    wire N__46749;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46741;
    wire N__46740;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46722;
    wire N__46713;
    wire N__46710;
    wire N__46709;
    wire N__46708;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46698;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46680;
    wire N__46679;
    wire N__46678;
    wire N__46675;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46659;
    wire N__46658;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46645;
    wire N__46638;
    wire N__46637;
    wire N__46634;
    wire N__46633;
    wire N__46630;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46614;
    wire N__46613;
    wire N__46612;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46593;
    wire N__46592;
    wire N__46591;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46581;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46569;
    wire N__46560;
    wire N__46559;
    wire N__46558;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46542;
    wire N__46541;
    wire N__46538;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46518;
    wire N__46515;
    wire N__46514;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46497;
    wire N__46496;
    wire N__46495;
    wire N__46492;
    wire N__46489;
    wire N__46486;
    wire N__46483;
    wire N__46476;
    wire N__46475;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46462;
    wire N__46455;
    wire N__46454;
    wire N__46451;
    wire N__46448;
    wire N__46445;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46425;
    wire N__46424;
    wire N__46421;
    wire N__46420;
    wire N__46419;
    wire N__46418;
    wire N__46415;
    wire N__46414;
    wire N__46411;
    wire N__46410;
    wire N__46409;
    wire N__46408;
    wire N__46405;
    wire N__46404;
    wire N__46399;
    wire N__46394;
    wire N__46391;
    wire N__46388;
    wire N__46385;
    wire N__46382;
    wire N__46377;
    wire N__46374;
    wire N__46371;
    wire N__46356;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46331;
    wire N__46328;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46310;
    wire N__46305;
    wire N__46302;
    wire N__46299;
    wire N__46296;
    wire N__46293;
    wire N__46290;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46266;
    wire N__46265;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46247;
    wire N__46244;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46199;
    wire N__46198;
    wire N__46197;
    wire N__46196;
    wire N__46195;
    wire N__46194;
    wire N__46193;
    wire N__46192;
    wire N__46191;
    wire N__46190;
    wire N__46189;
    wire N__46188;
    wire N__46187;
    wire N__46186;
    wire N__46185;
    wire N__46184;
    wire N__46183;
    wire N__46182;
    wire N__46181;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46173;
    wire N__46166;
    wire N__46165;
    wire N__46164;
    wire N__46161;
    wire N__46160;
    wire N__46159;
    wire N__46158;
    wire N__46155;
    wire N__46154;
    wire N__46153;
    wire N__46152;
    wire N__46151;
    wire N__46150;
    wire N__46145;
    wire N__46142;
    wire N__46133;
    wire N__46124;
    wire N__46121;
    wire N__46118;
    wire N__46115;
    wire N__46112;
    wire N__46107;
    wire N__46104;
    wire N__46103;
    wire N__46102;
    wire N__46099;
    wire N__46098;
    wire N__46091;
    wire N__46086;
    wire N__46083;
    wire N__46076;
    wire N__46071;
    wire N__46062;
    wire N__46061;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46032;
    wire N__46031;
    wire N__46030;
    wire N__46029;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46004;
    wire N__46001;
    wire N__45998;
    wire N__45987;
    wire N__45980;
    wire N__45971;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45941;
    wire N__45938;
    wire N__45935;
    wire N__45934;
    wire N__45931;
    wire N__45928;
    wire N__45925;
    wire N__45918;
    wire N__45915;
    wire N__45914;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45876;
    wire N__45875;
    wire N__45874;
    wire N__45871;
    wire N__45868;
    wire N__45865;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45815;
    wire N__45810;
    wire N__45809;
    wire N__45806;
    wire N__45803;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45789;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45761;
    wire N__45758;
    wire N__45755;
    wire N__45752;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45735;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45725;
    wire N__45722;
    wire N__45719;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45690;
    wire N__45687;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45669;
    wire N__45666;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45658;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45642;
    wire N__45641;
    wire N__45638;
    wire N__45635;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45586;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45545;
    wire N__45540;
    wire N__45537;
    wire N__45536;
    wire N__45535;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45515;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45494;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45471;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45459;
    wire N__45458;
    wire N__45455;
    wire N__45452;
    wire N__45449;
    wire N__45444;
    wire N__45443;
    wire N__45440;
    wire N__45437;
    wire N__45432;
    wire N__45429;
    wire N__45426;
    wire N__45423;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45381;
    wire N__45380;
    wire N__45379;
    wire N__45374;
    wire N__45371;
    wire N__45366;
    wire N__45365;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45348;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45285;
    wire N__45284;
    wire N__45281;
    wire N__45278;
    wire N__45275;
    wire N__45270;
    wire N__45269;
    wire N__45266;
    wire N__45263;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45188;
    wire N__45183;
    wire N__45180;
    wire N__45179;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45140;
    wire N__45137;
    wire N__45134;
    wire N__45133;
    wire N__45130;
    wire N__45125;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45083;
    wire N__45082;
    wire N__45079;
    wire N__45074;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45056;
    wire N__45053;
    wire N__45048;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45029;
    wire N__45026;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45009;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44987;
    wire N__44984;
    wire N__44981;
    wire N__44980;
    wire N__44977;
    wire N__44974;
    wire N__44971;
    wire N__44964;
    wire N__44963;
    wire N__44960;
    wire N__44957;
    wire N__44956;
    wire N__44955;
    wire N__44954;
    wire N__44953;
    wire N__44952;
    wire N__44949;
    wire N__44944;
    wire N__44941;
    wire N__44934;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44891;
    wire N__44888;
    wire N__44887;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44871;
    wire N__44870;
    wire N__44867;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44817;
    wire N__44814;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44804;
    wire N__44799;
    wire N__44798;
    wire N__44795;
    wire N__44792;
    wire N__44789;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44756;
    wire N__44753;
    wire N__44750;
    wire N__44745;
    wire N__44744;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44730;
    wire N__44729;
    wire N__44728;
    wire N__44723;
    wire N__44720;
    wire N__44717;
    wire N__44714;
    wire N__44711;
    wire N__44706;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44687;
    wire N__44684;
    wire N__44681;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44640;
    wire N__44637;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44606;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44583;
    wire N__44580;
    wire N__44579;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44569;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44544;
    wire N__44543;
    wire N__44540;
    wire N__44537;
    wire N__44534;
    wire N__44531;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44519;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44504;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44484;
    wire N__44481;
    wire N__44478;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44372;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44312;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44186;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44165;
    wire N__44164;
    wire N__44163;
    wire N__44160;
    wire N__44153;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44138;
    wire N__44135;
    wire N__44132;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44093;
    wire N__44090;
    wire N__44087;
    wire N__44084;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44063;
    wire N__44058;
    wire N__44055;
    wire N__44054;
    wire N__44051;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43958;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43934;
    wire N__43931;
    wire N__43928;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43908;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43898;
    wire N__43895;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43857;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43847;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43827;
    wire N__43824;
    wire N__43821;
    wire N__43820;
    wire N__43819;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43782;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43767;
    wire N__43764;
    wire N__43763;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43674;
    wire N__43673;
    wire N__43670;
    wire N__43667;
    wire N__43662;
    wire N__43659;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43611;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43598;
    wire N__43595;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43535;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43514;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43500;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43479;
    wire N__43478;
    wire N__43475;
    wire N__43472;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43448;
    wire N__43443;
    wire N__43440;
    wire N__43437;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43422;
    wire N__43421;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43352;
    wire N__43349;
    wire N__43346;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43325;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43311;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43226;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43208;
    wire N__43205;
    wire N__43202;
    wire N__43197;
    wire N__43194;
    wire N__43191;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43178;
    wire N__43175;
    wire N__43174;
    wire N__43173;
    wire N__43172;
    wire N__43171;
    wire N__43170;
    wire N__43169;
    wire N__43168;
    wire N__43167;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43156;
    wire N__43153;
    wire N__43152;
    wire N__43151;
    wire N__43150;
    wire N__43149;
    wire N__43148;
    wire N__43147;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43135;
    wire N__43134;
    wire N__43133;
    wire N__43130;
    wire N__43129;
    wire N__43126;
    wire N__43125;
    wire N__43124;
    wire N__43121;
    wire N__43118;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43106;
    wire N__43097;
    wire N__43094;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43086;
    wire N__43085;
    wire N__43082;
    wire N__43073;
    wire N__43066;
    wire N__43057;
    wire N__43048;
    wire N__43039;
    wire N__43026;
    wire N__43011;
    wire N__43010;
    wire N__43007;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42995;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42983;
    wire N__42978;
    wire N__42975;
    wire N__42972;
    wire N__42969;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42948;
    wire N__42945;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42932;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42912;
    wire N__42909;
    wire N__42906;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42873;
    wire N__42870;
    wire N__42867;
    wire N__42866;
    wire N__42865;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42849;
    wire N__42848;
    wire N__42847;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42829;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42815;
    wire N__42814;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42798;
    wire N__42793;
    wire N__42786;
    wire N__42783;
    wire N__42782;
    wire N__42779;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42729;
    wire N__42728;
    wire N__42725;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42715;
    wire N__42710;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42683;
    wire N__42682;
    wire N__42679;
    wire N__42676;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42539;
    wire N__42538;
    wire N__42535;
    wire N__42530;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42515;
    wire N__42512;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42500;
    wire N__42495;
    wire N__42492;
    wire N__42489;
    wire N__42486;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42443;
    wire N__42438;
    wire N__42437;
    wire N__42434;
    wire N__42431;
    wire N__42428;
    wire N__42423;
    wire N__42420;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42410;
    wire N__42407;
    wire N__42406;
    wire N__42403;
    wire N__42400;
    wire N__42397;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42374;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42316;
    wire N__42311;
    wire N__42308;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42290;
    wire N__42289;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42267;
    wire N__42264;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42251;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42225;
    wire N__42224;
    wire N__42221;
    wire N__42220;
    wire N__42217;
    wire N__42214;
    wire N__42211;
    wire N__42204;
    wire N__42201;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42191;
    wire N__42190;
    wire N__42189;
    wire N__42188;
    wire N__42187;
    wire N__42186;
    wire N__42185;
    wire N__42184;
    wire N__42183;
    wire N__42182;
    wire N__42181;
    wire N__42180;
    wire N__42179;
    wire N__42178;
    wire N__42177;
    wire N__42176;
    wire N__42175;
    wire N__42174;
    wire N__42173;
    wire N__42172;
    wire N__42171;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42102;
    wire N__42093;
    wire N__42084;
    wire N__42075;
    wire N__42066;
    wire N__42057;
    wire N__42048;
    wire N__42045;
    wire N__42040;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42022;
    wire N__42017;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41993;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41977;
    wire N__41974;
    wire N__41971;
    wire N__41968;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41918;
    wire N__41915;
    wire N__41912;
    wire N__41909;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41855;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41845;
    wire N__41838;
    wire N__41835;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41827;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41810;
    wire N__41805;
    wire N__41804;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41796;
    wire N__41793;
    wire N__41792;
    wire N__41791;
    wire N__41790;
    wire N__41789;
    wire N__41786;
    wire N__41785;
    wire N__41780;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41770;
    wire N__41769;
    wire N__41768;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41760;
    wire N__41759;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41747;
    wire N__41738;
    wire N__41727;
    wire N__41722;
    wire N__41709;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41693;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41681;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41660;
    wire N__41657;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41628;
    wire N__41627;
    wire N__41626;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41591;
    wire N__41588;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41530;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41499;
    wire N__41496;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41486;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41471;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41432;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41321;
    wire N__41320;
    wire N__41317;
    wire N__41312;
    wire N__41309;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41291;
    wire N__41290;
    wire N__41287;
    wire N__41282;
    wire N__41279;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41261;
    wire N__41258;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41197;
    wire N__41192;
    wire N__41189;
    wire N__41184;
    wire N__41181;
    wire N__41180;
    wire N__41179;
    wire N__41174;
    wire N__41171;
    wire N__41166;
    wire N__41163;
    wire N__41162;
    wire N__41161;
    wire N__41156;
    wire N__41153;
    wire N__41148;
    wire N__41145;
    wire N__41144;
    wire N__41143;
    wire N__41138;
    wire N__41135;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40910;
    wire N__40909;
    wire N__40906;
    wire N__40901;
    wire N__40896;
    wire N__40895;
    wire N__40894;
    wire N__40891;
    wire N__40886;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40866;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40752;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40736;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40707;
    wire N__40706;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40694;
    wire N__40689;
    wire N__40688;
    wire N__40685;
    wire N__40684;
    wire N__40681;
    wire N__40680;
    wire N__40675;
    wire N__40670;
    wire N__40665;
    wire N__40664;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40632;
    wire N__40629;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40589;
    wire N__40586;
    wire N__40583;
    wire N__40580;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40563;
    wire N__40560;
    wire N__40559;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40524;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40493;
    wire N__40490;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40473;
    wire N__40472;
    wire N__40467;
    wire N__40464;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40452;
    wire N__40449;
    wire N__40446;
    wire N__40443;
    wire N__40442;
    wire N__40441;
    wire N__40438;
    wire N__40433;
    wire N__40428;
    wire N__40427;
    wire N__40426;
    wire N__40423;
    wire N__40420;
    wire N__40417;
    wire N__40416;
    wire N__40413;
    wire N__40408;
    wire N__40405;
    wire N__40398;
    wire N__40397;
    wire N__40394;
    wire N__40393;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40355;
    wire N__40352;
    wire N__40351;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40328;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40305;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40274;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40263;
    wire N__40262;
    wire N__40261;
    wire N__40258;
    wire N__40247;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40125;
    wire N__40122;
    wire N__40121;
    wire N__40118;
    wire N__40117;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40105;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40076;
    wire N__40073;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40056;
    wire N__40055;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40008;
    wire N__40007;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39950;
    wire N__39947;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39932;
    wire N__39927;
    wire N__39926;
    wire N__39923;
    wire N__39920;
    wire N__39915;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39884;
    wire N__39883;
    wire N__39882;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39874;
    wire N__39873;
    wire N__39872;
    wire N__39869;
    wire N__39868;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39860;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39845;
    wire N__39842;
    wire N__39841;
    wire N__39840;
    wire N__39839;
    wire N__39838;
    wire N__39835;
    wire N__39830;
    wire N__39821;
    wire N__39816;
    wire N__39807;
    wire N__39802;
    wire N__39795;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39737;
    wire N__39734;
    wire N__39731;
    wire N__39730;
    wire N__39725;
    wire N__39722;
    wire N__39717;
    wire N__39716;
    wire N__39713;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39703;
    wire N__39698;
    wire N__39695;
    wire N__39690;
    wire N__39687;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39666;
    wire N__39663;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39635;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39543;
    wire N__39540;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39516;
    wire N__39513;
    wire N__39508;
    wire N__39505;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39399;
    wire N__39396;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39384;
    wire N__39383;
    wire N__39382;
    wire N__39379;
    wire N__39374;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39212;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39161;
    wire N__39160;
    wire N__39159;
    wire N__39152;
    wire N__39149;
    wire N__39144;
    wire N__39143;
    wire N__39138;
    wire N__39135;
    wire N__39134;
    wire N__39133;
    wire N__39130;
    wire N__39125;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39113;
    wire N__39112;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39081;
    wire N__39080;
    wire N__39077;
    wire N__39076;
    wire N__39075;
    wire N__39074;
    wire N__39071;
    wire N__39070;
    wire N__39067;
    wire N__39060;
    wire N__39055;
    wire N__39048;
    wire N__39045;
    wire N__39044;
    wire N__39043;
    wire N__39042;
    wire N__39039;
    wire N__39034;
    wire N__39031;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38961;
    wire N__38958;
    wire N__38957;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38942;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38927;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38456;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38423;
    wire N__38420;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38403;
    wire N__38402;
    wire N__38399;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38378;
    wire N__38375;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38360;
    wire N__38359;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38302;
    wire N__38297;
    wire N__38294;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38269;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38255;
    wire N__38250;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38234;
    wire N__38233;
    wire N__38228;
    wire N__38225;
    wire N__38222;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38210;
    wire N__38209;
    wire N__38208;
    wire N__38207;
    wire N__38206;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38198;
    wire N__38197;
    wire N__38196;
    wire N__38195;
    wire N__38192;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38184;
    wire N__38181;
    wire N__38180;
    wire N__38179;
    wire N__38178;
    wire N__38175;
    wire N__38174;
    wire N__38173;
    wire N__38168;
    wire N__38161;
    wire N__38148;
    wire N__38143;
    wire N__38134;
    wire N__38131;
    wire N__38118;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38100;
    wire N__38099;
    wire N__38096;
    wire N__38093;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38011;
    wire N__38006;
    wire N__38003;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37952;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37926;
    wire N__37923;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37887;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37874;
    wire N__37871;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37825;
    wire N__37818;
    wire N__37817;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37787;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37770;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37752;
    wire N__37749;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37725;
    wire N__37722;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37646;
    wire N__37641;
    wire N__37640;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37578;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37467;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37424;
    wire N__37423;
    wire N__37422;
    wire N__37421;
    wire N__37420;
    wire N__37419;
    wire N__37418;
    wire N__37417;
    wire N__37416;
    wire N__37415;
    wire N__37414;
    wire N__37413;
    wire N__37412;
    wire N__37411;
    wire N__37408;
    wire N__37407;
    wire N__37404;
    wire N__37403;
    wire N__37400;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37392;
    wire N__37389;
    wire N__37388;
    wire N__37385;
    wire N__37384;
    wire N__37381;
    wire N__37380;
    wire N__37379;
    wire N__37376;
    wire N__37375;
    wire N__37372;
    wire N__37371;
    wire N__37368;
    wire N__37367;
    wire N__37366;
    wire N__37365;
    wire N__37362;
    wire N__37361;
    wire N__37358;
    wire N__37357;
    wire N__37354;
    wire N__37353;
    wire N__37336;
    wire N__37319;
    wire N__37304;
    wire N__37287;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37269;
    wire N__37266;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37223;
    wire N__37220;
    wire N__37219;
    wire N__37218;
    wire N__37217;
    wire N__37216;
    wire N__37215;
    wire N__37212;
    wire N__37211;
    wire N__37210;
    wire N__37207;
    wire N__37206;
    wire N__37205;
    wire N__37204;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37196;
    wire N__37195;
    wire N__37194;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37171;
    wire N__37170;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37162;
    wire N__37159;
    wire N__37158;
    wire N__37157;
    wire N__37156;
    wire N__37155;
    wire N__37154;
    wire N__37153;
    wire N__37150;
    wire N__37149;
    wire N__37146;
    wire N__37141;
    wire N__37132;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37113;
    wire N__37110;
    wire N__37101;
    wire N__37096;
    wire N__37093;
    wire N__37088;
    wire N__37079;
    wire N__37070;
    wire N__37065;
    wire N__37044;
    wire N__37043;
    wire N__37040;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36992;
    wire N__36991;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36909;
    wire N__36906;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36876;
    wire N__36875;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36845;
    wire N__36842;
    wire N__36837;
    wire N__36836;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36773;
    wire N__36768;
    wire N__36765;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36719;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36665;
    wire N__36664;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36632;
    wire N__36627;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36612;
    wire N__36609;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36578;
    wire N__36573;
    wire N__36570;
    wire N__36569;
    wire N__36566;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36551;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36536;
    wire N__36533;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36503;
    wire N__36500;
    wire N__36499;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36414;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36381;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36336;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36317;
    wire N__36316;
    wire N__36313;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36243;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36207;
    wire N__36204;
    wire N__36203;
    wire N__36200;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36182;
    wire N__36177;
    wire N__36174;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36036;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36014;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35987;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35969;
    wire N__35968;
    wire N__35965;
    wire N__35960;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35918;
    wire N__35917;
    wire N__35914;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35879;
    wire N__35876;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35834;
    wire N__35833;
    wire N__35830;
    wire N__35825;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35802;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35705;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35670;
    wire N__35667;
    wire N__35666;
    wire N__35663;
    wire N__35660;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35619;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35577;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35560;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35546;
    wire N__35543;
    wire N__35538;
    wire N__35535;
    wire N__35532;
    wire N__35529;
    wire N__35526;
    wire N__35525;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35481;
    wire N__35478;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35470;
    wire N__35465;
    wire N__35462;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35358;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35350;
    wire N__35345;
    wire N__35342;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35260;
    wire N__35257;
    wire N__35252;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35232;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35205;
    wire N__35202;
    wire N__35199;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35126;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35099;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35042;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34952;
    wire N__34949;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34824;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34781;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34730;
    wire N__34729;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34725;
    wire N__34722;
    wire N__34721;
    wire N__34720;
    wire N__34717;
    wire N__34716;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34708;
    wire N__34707;
    wire N__34704;
    wire N__34703;
    wire N__34702;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34696;
    wire N__34687;
    wire N__34678;
    wire N__34665;
    wire N__34664;
    wire N__34663;
    wire N__34660;
    wire N__34657;
    wire N__34656;
    wire N__34655;
    wire N__34652;
    wire N__34651;
    wire N__34648;
    wire N__34641;
    wire N__34636;
    wire N__34635;
    wire N__34634;
    wire N__34633;
    wire N__34632;
    wire N__34631;
    wire N__34630;
    wire N__34629;
    wire N__34626;
    wire N__34615;
    wire N__34608;
    wire N__34599;
    wire N__34594;
    wire N__34591;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34556;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34517;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34457;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34331;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34248;
    wire N__34245;
    wire N__34244;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34173;
    wire N__34170;
    wire N__34169;
    wire N__34168;
    wire N__34167;
    wire N__34164;
    wire N__34163;
    wire N__34162;
    wire N__34161;
    wire N__34160;
    wire N__34159;
    wire N__34156;
    wire N__34155;
    wire N__34154;
    wire N__34153;
    wire N__34152;
    wire N__34149;
    wire N__34148;
    wire N__34145;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34137;
    wire N__34134;
    wire N__34133;
    wire N__34130;
    wire N__34129;
    wire N__34128;
    wire N__34127;
    wire N__34122;
    wire N__34119;
    wire N__34114;
    wire N__34109;
    wire N__34104;
    wire N__34099;
    wire N__34094;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34070;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34029;
    wire N__34028;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34024;
    wire N__34021;
    wire N__34020;
    wire N__34019;
    wire N__34018;
    wire N__34017;
    wire N__34016;
    wire N__34015;
    wire N__34012;
    wire N__34011;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34003;
    wire N__34002;
    wire N__33997;
    wire N__33994;
    wire N__33989;
    wire N__33986;
    wire N__33985;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33977;
    wire N__33974;
    wire N__33967;
    wire N__33958;
    wire N__33955;
    wire N__33948;
    wire N__33943;
    wire N__33936;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33900;
    wire N__33897;
    wire N__33896;
    wire N__33895;
    wire N__33894;
    wire N__33893;
    wire N__33892;
    wire N__33891;
    wire N__33888;
    wire N__33887;
    wire N__33886;
    wire N__33881;
    wire N__33874;
    wire N__33873;
    wire N__33872;
    wire N__33871;
    wire N__33868;
    wire N__33867;
    wire N__33866;
    wire N__33865;
    wire N__33864;
    wire N__33863;
    wire N__33862;
    wire N__33859;
    wire N__33858;
    wire N__33855;
    wire N__33854;
    wire N__33851;
    wire N__33850;
    wire N__33849;
    wire N__33846;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33830;
    wire N__33825;
    wire N__33818;
    wire N__33815;
    wire N__33808;
    wire N__33805;
    wire N__33804;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33796;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33777;
    wire N__33770;
    wire N__33759;
    wire N__33756;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33714;
    wire N__33713;
    wire N__33710;
    wire N__33709;
    wire N__33708;
    wire N__33707;
    wire N__33706;
    wire N__33705;
    wire N__33702;
    wire N__33701;
    wire N__33700;
    wire N__33699;
    wire N__33698;
    wire N__33697;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33669;
    wire N__33668;
    wire N__33667;
    wire N__33664;
    wire N__33663;
    wire N__33662;
    wire N__33661;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33655;
    wire N__33652;
    wire N__33651;
    wire N__33648;
    wire N__33647;
    wire N__33646;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33616;
    wire N__33607;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33583;
    wire N__33574;
    wire N__33555;
    wire N__33552;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33528;
    wire N__33525;
    wire N__33524;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33518;
    wire N__33517;
    wire N__33516;
    wire N__33515;
    wire N__33514;
    wire N__33513;
    wire N__33512;
    wire N__33511;
    wire N__33510;
    wire N__33507;
    wire N__33506;
    wire N__33505;
    wire N__33504;
    wire N__33503;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33492;
    wire N__33491;
    wire N__33488;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33470;
    wire N__33465;
    wire N__33464;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33456;
    wire N__33453;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33445;
    wire N__33432;
    wire N__33427;
    wire N__33416;
    wire N__33413;
    wire N__33408;
    wire N__33405;
    wire N__33400;
    wire N__33389;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33351;
    wire N__33350;
    wire N__33349;
    wire N__33346;
    wire N__33345;
    wire N__33344;
    wire N__33343;
    wire N__33342;
    wire N__33341;
    wire N__33340;
    wire N__33339;
    wire N__33336;
    wire N__33335;
    wire N__33334;
    wire N__33331;
    wire N__33330;
    wire N__33329;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33314;
    wire N__33311;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33303;
    wire N__33302;
    wire N__33301;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33293;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33278;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33270;
    wire N__33265;
    wire N__33260;
    wire N__33253;
    wire N__33244;
    wire N__33235;
    wire N__33226;
    wire N__33215;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33171;
    wire N__33170;
    wire N__33167;
    wire N__33166;
    wire N__33165;
    wire N__33164;
    wire N__33163;
    wire N__33160;
    wire N__33159;
    wire N__33158;
    wire N__33157;
    wire N__33156;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33148;
    wire N__33145;
    wire N__33140;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33128;
    wire N__33127;
    wire N__33126;
    wire N__33125;
    wire N__33122;
    wire N__33121;
    wire N__33120;
    wire N__33119;
    wire N__33118;
    wire N__33115;
    wire N__33114;
    wire N__33111;
    wire N__33110;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33095;
    wire N__33092;
    wire N__33083;
    wire N__33070;
    wire N__33065;
    wire N__33054;
    wire N__33045;
    wire N__33042;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33000;
    wire N__32999;
    wire N__32998;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32977;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32966;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32958;
    wire N__32955;
    wire N__32954;
    wire N__32953;
    wire N__32952;
    wire N__32947;
    wire N__32946;
    wire N__32945;
    wire N__32942;
    wire N__32941;
    wire N__32940;
    wire N__32937;
    wire N__32930;
    wire N__32927;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32907;
    wire N__32906;
    wire N__32905;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32887;
    wire N__32882;
    wire N__32879;
    wire N__32866;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32846;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32829;
    wire N__32828;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32820;
    wire N__32819;
    wire N__32818;
    wire N__32817;
    wire N__32814;
    wire N__32813;
    wire N__32812;
    wire N__32809;
    wire N__32808;
    wire N__32807;
    wire N__32806;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32798;
    wire N__32795;
    wire N__32794;
    wire N__32793;
    wire N__32792;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32782;
    wire N__32779;
    wire N__32772;
    wire N__32769;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32753;
    wire N__32742;
    wire N__32731;
    wire N__32726;
    wire N__32721;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32685;
    wire N__32684;
    wire N__32683;
    wire N__32682;
    wire N__32681;
    wire N__32680;
    wire N__32677;
    wire N__32676;
    wire N__32673;
    wire N__32672;
    wire N__32671;
    wire N__32668;
    wire N__32665;
    wire N__32664;
    wire N__32661;
    wire N__32660;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32632;
    wire N__32627;
    wire N__32618;
    wire N__32615;
    wire N__32614;
    wire N__32613;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32597;
    wire N__32594;
    wire N__32589;
    wire N__32586;
    wire N__32581;
    wire N__32578;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32562;
    wire N__32555;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32511;
    wire N__32508;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32474;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32453;
    wire N__32450;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32433;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32425;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32336;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32289;
    wire N__32286;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32236;
    wire N__32231;
    wire N__32228;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32193;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32183;
    wire N__32182;
    wire N__32179;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32124;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32107;
    wire N__32100;
    wire N__32097;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32057;
    wire N__32054;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32037;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31977;
    wire N__31974;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31944;
    wire N__31941;
    wire N__31940;
    wire N__31937;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31908;
    wire N__31905;
    wire N__31904;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31848;
    wire N__31847;
    wire N__31844;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31827;
    wire N__31824;
    wire N__31823;
    wire N__31822;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31797;
    wire N__31794;
    wire N__31793;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31751;
    wire N__31748;
    wire N__31745;
    wire N__31742;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31629;
    wire N__31628;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31585;
    wire N__31580;
    wire N__31577;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31496;
    wire N__31493;
    wire N__31490;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31441;
    wire N__31436;
    wire N__31433;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31385;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31370;
    wire N__31367;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31202;
    wire N__31201;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31139;
    wire N__31138;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31126;
    wire N__31121;
    wire N__31118;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31076;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31055;
    wire N__31050;
    wire N__31047;
    wire N__31046;
    wire N__31043;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30988;
    wire N__30985;
    wire N__30982;
    wire N__30979;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30920;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30897;
    wire N__30894;
    wire N__30893;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30876;
    wire N__30873;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30848;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30819;
    wire N__30816;
    wire N__30815;
    wire N__30814;
    wire N__30811;
    wire N__30806;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30672;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30548;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30456;
    wire N__30453;
    wire N__30452;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30405;
    wire N__30404;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30381;
    wire N__30380;
    wire N__30377;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30353;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30320;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30251;
    wire N__30248;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30173;
    wire N__30172;
    wire N__30169;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30146;
    wire N__30145;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30078;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30046;
    wire N__30041;
    wire N__30038;
    wire N__30033;
    wire N__30030;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30002;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29940;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29925;
    wire N__29924;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29906;
    wire N__29901;
    wire N__29898;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29848;
    wire N__29843;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29816;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29753;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29702;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29666;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29649;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29637;
    wire N__29634;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29570;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29558;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29504;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29400;
    wire N__29397;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29360;
    wire N__29357;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29234;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29216;
    wire N__29211;
    wire N__29208;
    wire N__29207;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29171;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29093;
    wire N__29092;
    wire N__29089;
    wire N__29084;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29037;
    wire N__29034;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28718;
    wire N__28713;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28691;
    wire N__28688;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28670;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28638;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28618;
    wire N__28613;
    wire N__28610;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28536;
    wire N__28535;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28506;
    wire N__28503;
    wire N__28502;
    wire N__28499;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28166;
    wire N__28163;
    wire N__28162;
    wire N__28159;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28143;
    wire N__28140;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28075;
    wire N__28070;
    wire N__28067;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27912;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27833;
    wire N__27830;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27809;
    wire N__27804;
    wire N__27801;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27751;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27709;
    wire N__27704;
    wire N__27701;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27641;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27575;
    wire N__27572;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27555;
    wire N__27552;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27453;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27404;
    wire N__27401;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27371;
    wire N__27368;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27315;
    wire N__27312;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27284;
    wire N__27283;
    wire N__27280;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27197;
    wire N__27194;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27095;
    wire N__27092;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27028;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26998;
    wire N__26993;
    wire N__26990;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26822;
    wire N__26819;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26783;
    wire N__26780;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26718;
    wire N__26717;
    wire N__26714;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26697;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26673;
    wire N__26670;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26609;
    wire N__26606;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26514;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26478;
    wire N__26475;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26424;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26351;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26297;
    wire N__26292;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26265;
    wire N__26262;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26242;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26177;
    wire N__26174;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26100;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26075;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26060;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26032;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25997;
    wire N__25996;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25829;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25763;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25730;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25655;
    wire N__25654;
    wire N__25651;
    wire N__25646;
    wire N__25641;
    wire N__25638;
    wire N__25637;
    wire N__25636;
    wire N__25633;
    wire N__25628;
    wire N__25623;
    wire N__25620;
    wire N__25619;
    wire N__25616;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25503;
    wire N__25502;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25485;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25460;
    wire N__25457;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24985;
    wire N__24980;
    wire N__24977;
    wire N__24972;
    wire N__24971;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24911;
    wire N__24910;
    wire N__24907;
    wire N__24902;
    wire N__24897;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24873;
    wire N__24872;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24862;
    wire N__24857;
    wire N__24854;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24788;
    wire N__24785;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24704;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24650;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24536;
    wire N__24535;
    wire N__24532;
    wire N__24527;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24515;
    wire N__24514;
    wire N__24511;
    wire N__24506;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24494;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24477;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24410;
    wire N__24405;
    wire N__24402;
    wire N__24401;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24329;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24312;
    wire N__24311;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24291;
    wire N__24288;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24233;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24218;
    wire N__24213;
    wire N__24210;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24192;
    wire N__24189;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24178;
    wire N__24175;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24114;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24062;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23964;
    wire N__23963;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23945;
    wire N__23942;
    wire N__23937;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23929;
    wire N__23924;
    wire N__23921;
    wire N__23916;
    wire N__23913;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23892;
    wire N__23889;
    wire N__23888;
    wire N__23887;
    wire N__23884;
    wire N__23879;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23658;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23645;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23627;
    wire N__23624;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23565;
    wire N__23564;
    wire N__23561;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23446;
    wire N__23441;
    wire N__23438;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23372;
    wire N__23369;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23352;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23341;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23325;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23298;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23286;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23253;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23196;
    wire N__23193;
    wire N__23192;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23175;
    wire N__23174;
    wire N__23171;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23144;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23124;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23103;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23079;
    wire N__23076;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23022;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23010;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22865;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22848;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22793;
    wire N__22792;
    wire N__22789;
    wire N__22784;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22757;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22727;
    wire N__22724;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22706;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22492;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22348;
    wire N__22343;
    wire N__22340;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22312;
    wire N__22307;
    wire N__22304;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22196;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_17_0_;
    wire n12703;
    wire n12704;
    wire n12705;
    wire n12706;
    wire n12707;
    wire n12708;
    wire n12709;
    wire n12710;
    wire bfn_1_18_0_;
    wire n12711;
    wire n12712;
    wire n12713;
    wire n12714;
    wire n12715;
    wire n12716;
    wire n12717;
    wire n12718;
    wire bfn_1_19_0_;
    wire n12719;
    wire n12720;
    wire n12721;
    wire n12722;
    wire n12723;
    wire n12724;
    wire bfn_1_20_0_;
    wire n12725;
    wire n12726;
    wire n12727;
    wire n12728;
    wire n12729;
    wire n12730;
    wire n12731;
    wire n12732;
    wire bfn_1_21_0_;
    wire n12733;
    wire n12734;
    wire n12735;
    wire n12736;
    wire n12737;
    wire n12738;
    wire n12739;
    wire n12740;
    wire bfn_1_22_0_;
    wire n12741;
    wire n12742;
    wire n12743;
    wire n12744;
    wire n12745;
    wire n12746;
    wire n12747;
    wire n2719_cascade_;
    wire n2486;
    wire n2816_cascade_;
    wire n2829_cascade_;
    wire n13845_cascade_;
    wire n14702;
    wire bfn_1_26_0_;
    wire n12797;
    wire n12798;
    wire n12799;
    wire n12800;
    wire n12801;
    wire n12802;
    wire n12803;
    wire n12804;
    wire bfn_1_27_0_;
    wire n12805;
    wire n12806;
    wire n12807;
    wire n12808;
    wire n12809;
    wire n12810;
    wire n12811;
    wire n12812;
    wire bfn_1_28_0_;
    wire n12813;
    wire n12814;
    wire n12815;
    wire n12816;
    wire n12817;
    wire n12818;
    wire n12819;
    wire n12820;
    wire bfn_1_29_0_;
    wire n2876;
    wire n12821;
    wire n12822;
    wire n11956;
    wire n2899;
    wire n2833;
    wire n2900;
    wire n2833_cascade_;
    wire n2932_cascade_;
    wire n2901;
    wire n2933_cascade_;
    wire bfn_1_31_0_;
    wire \debounce.n13016 ;
    wire \debounce.n13017 ;
    wire \debounce.n13018 ;
    wire \debounce.n13019 ;
    wire \debounce.n13020 ;
    wire \debounce.n13021 ;
    wire \debounce.n13022 ;
    wire \debounce.n13023 ;
    wire bfn_1_32_0_;
    wire \debounce.n13024 ;
    wire n2501;
    wire n2500;
    wire n2433_cascade_;
    wire n2532_cascade_;
    wire n2498;
    wire n2487;
    wire n2497;
    wire n2499;
    wire n2496;
    wire n2418_cascade_;
    wire n2495;
    wire n2428_cascade_;
    wire n2527_cascade_;
    wire n2488;
    wire n2493;
    wire n2490;
    wire n2418;
    wire n2485;
    wire n2491;
    wire n2481;
    wire n14310;
    wire n2494;
    wire n2483;
    wire n2416;
    wire n2480;
    wire n2482;
    wire n14650_cascade_;
    wire n2595;
    wire n2528;
    wire n2627_cascade_;
    wire n14646;
    wire n2520;
    wire n2587;
    wire n2589;
    wire n2522;
    wire n2596;
    wire n2628_cascade_;
    wire n14644;
    wire n2527;
    wire n2594;
    wire n2579;
    wire n2586;
    wire n2519;
    wire n2484;
    wire n2583;
    wire n2516_cascade_;
    wire n2588;
    wire n2580;
    wire n2612_cascade_;
    wire n2801;
    wire bfn_2_23_0_;
    wire n12772;
    wire n2799;
    wire n12773;
    wire n2798;
    wire n12774;
    wire n2797;
    wire n12775;
    wire n12776;
    wire n12777;
    wire n12778;
    wire n12779;
    wire bfn_2_24_0_;
    wire n12780;
    wire n12781;
    wire n12782;
    wire n12783;
    wire n12784;
    wire n12785;
    wire n2719;
    wire n2786;
    wire n12786;
    wire n12787;
    wire n2785;
    wire bfn_2_25_0_;
    wire n2784;
    wire n12788;
    wire n2783;
    wire n12789;
    wire n2782;
    wire n12790;
    wire n12791;
    wire n12792;
    wire n12793;
    wire n12794;
    wire n12795;
    wire bfn_2_26_0_;
    wire n12796;
    wire n14158_cascade_;
    wire n2790;
    wire n2742_cascade_;
    wire n2789;
    wire n2711;
    wire n2778;
    wire n2781;
    wire n2714;
    wire n2800;
    wire n2832;
    wire n2794;
    wire n2887;
    wire n2779;
    wire n2811_cascade_;
    wire n14708;
    wire n2780;
    wire n2817;
    wire n2884;
    wire n2877;
    wire n2897;
    wire n2830;
    wire n2811;
    wire n2878;
    wire bfn_2_29_0_;
    wire n2933;
    wire n3000;
    wire n12823;
    wire n12824;
    wire n12825;
    wire n12826;
    wire n12827;
    wire n12828;
    wire n12829;
    wire n12830;
    wire bfn_2_30_0_;
    wire n12831;
    wire n12832;
    wire n12833;
    wire n12834;
    wire n12835;
    wire n12836;
    wire n12837;
    wire n12838;
    wire bfn_2_31_0_;
    wire n12839;
    wire n12840;
    wire n12841;
    wire n12842;
    wire n12843;
    wire n12844;
    wire n12845;
    wire n12846;
    wire bfn_2_32_0_;
    wire n12847;
    wire n12848;
    wire n12849;
    wire \debounce.cnt_reg_0 ;
    wire \debounce.cnt_reg_7 ;
    wire \debounce.cnt_reg_1 ;
    wire \debounce.cnt_reg_2 ;
    wire \debounce.cnt_reg_9 ;
    wire \debounce.cnt_reg_8 ;
    wire \debounce.cnt_reg_4 ;
    wire \debounce.cnt_reg_5 ;
    wire n2976;
    wire n2432;
    wire n2432_cascade_;
    wire n2433;
    wire n2431;
    wire n2430;
    wire n11946_cascade_;
    wire n2429;
    wire n2427;
    wire n2424;
    wire n2427_cascade_;
    wire n2428;
    wire n2529;
    wire n11942;
    wire n13816;
    wire n14622_cascade_;
    wire n14638;
    wire n2420;
    wire n2420_cascade_;
    wire n14612;
    wire n14616;
    wire n2426;
    wire n2421;
    wire n2413;
    wire n2423;
    wire n2425_cascade_;
    wire n14632;
    wire n2419;
    wire n2415;
    wire n14456_cascade_;
    wire n2346_cascade_;
    wire n2417;
    wire n2414;
    wire n13790;
    wire n14318;
    wire n2328_cascade_;
    wire n14442_cascade_;
    wire n14448_cascade_;
    wire n14450;
    wire n2593;
    wire n2422;
    wire n2489;
    wire n2521;
    wire n2526;
    wire n2521_cascade_;
    wire n14312;
    wire n14324;
    wire n2516;
    wire n2512;
    wire n2513;
    wire n14330_cascade_;
    wire n2511;
    wire n2523;
    wire n2544_cascade_;
    wire n2590;
    wire n2591;
    wire n2530;
    wire n2597;
    wire n2629_cascade_;
    wire n14656;
    wire n2601;
    wire n2584;
    wire n2517;
    wire n2582;
    wire n2515;
    wire n2531;
    wire n2598;
    wire n2727;
    wire n2585;
    wire n2518;
    wire n14658;
    wire n2617_cascade_;
    wire n2514;
    wire n2581;
    wire n2613_cascade_;
    wire n14664;
    wire n14670_cascade_;
    wire n2643_cascade_;
    wire n2713;
    wire n2592;
    wire n14889_cascade_;
    wire n2525;
    wire n2721_cascade_;
    wire n2717;
    wire n2718;
    wire n14140_cascade_;
    wire n14138;
    wire n2716;
    wire n2715;
    wire n14146_cascade_;
    wire n14152;
    wire n2722;
    wire n2787;
    wire n2795;
    wire n2728;
    wire n2712;
    wire n2725;
    wire n2792;
    wire n2721;
    wire n2788;
    wire n2793;
    wire n2889;
    wire n2921_cascade_;
    wire n2888;
    wire n2791;
    wire n2822;
    wire n2823_cascade_;
    wire n2821;
    wire n2777;
    wire n2710;
    wire n2809;
    wire n2810;
    wire n2808;
    wire n2809_cascade_;
    wire n14714;
    wire n2823;
    wire n2841_cascade_;
    wire n2890;
    wire n2920;
    wire n2987;
    wire n2898;
    wire n2831;
    wire n2879;
    wire n2812;
    wire n2911_cascade_;
    wire n2829;
    wire n2896;
    wire n2893;
    wire n2826;
    wire n2882;
    wire n2815;
    wire n2813;
    wire n2880;
    wire bfn_3_29_0_;
    wire n12850;
    wire n12851;
    wire n12852;
    wire n12853;
    wire n12854;
    wire n12855;
    wire n12856;
    wire n12857;
    wire bfn_3_30_0_;
    wire n12858;
    wire n12859;
    wire n12860;
    wire n12861;
    wire n12862;
    wire n12863;
    wire n3086;
    wire n12864;
    wire n12865;
    wire bfn_3_31_0_;
    wire n12866;
    wire n12867;
    wire n12868;
    wire n12869;
    wire n12870;
    wire n12871;
    wire n12872;
    wire n12873;
    wire bfn_3_32_0_;
    wire n12874;
    wire n12875;
    wire n12876;
    wire n12877;
    wire \debounce.cnt_reg_6 ;
    wire \debounce.n16 ;
    wire \debounce.cnt_reg_3 ;
    wire \debounce.n17 ;
    wire n2401;
    wire bfn_4_17_0_;
    wire n2400;
    wire n12682;
    wire n2399;
    wire n12683;
    wire n2398;
    wire n12684;
    wire n2397;
    wire n12685;
    wire n2329;
    wire n2396;
    wire n12686;
    wire n2328;
    wire n2395;
    wire n12687;
    wire n2394;
    wire n12688;
    wire n12689;
    wire n2393;
    wire bfn_4_18_0_;
    wire n2392;
    wire n12690;
    wire n2391;
    wire n12691;
    wire n2390;
    wire n12692;
    wire n2389;
    wire n12693;
    wire n2388;
    wire n12694;
    wire n2387;
    wire n12695;
    wire n2386;
    wire n12696;
    wire n12697;
    wire n2385;
    wire bfn_4_19_0_;
    wire n2384;
    wire n12698;
    wire n2383;
    wire n12699;
    wire n2382;
    wire n12700;
    wire n2381;
    wire n12701;
    wire n12702;
    wire n2412;
    wire n2314_adj_622;
    wire n2327;
    wire n2327_cascade_;
    wire n2326;
    wire n14440;
    wire n2492;
    wire n2425;
    wire n2524;
    wire n2318;
    wire n2320;
    wire n2319;
    wire bfn_4_21_0_;
    wire n2700;
    wire n12748;
    wire n12749;
    wire n12750;
    wire n12751;
    wire n2629;
    wire n2696;
    wire n12752;
    wire n2628;
    wire n2695;
    wire n12753;
    wire n2627;
    wire n2694;
    wire n12754;
    wire n12755;
    wire n2626;
    wire n2693;
    wire bfn_4_22_0_;
    wire n2625;
    wire n2692;
    wire n12756;
    wire n2624;
    wire n2691;
    wire n12757;
    wire n2623;
    wire n2690;
    wire n12758;
    wire n2622;
    wire n2689;
    wire n12759;
    wire n12760;
    wire n2620;
    wire n2687;
    wire n12761;
    wire n2619;
    wire n2686;
    wire n12762;
    wire n12763;
    wire n2618;
    wire n2685;
    wire bfn_4_23_0_;
    wire n2617;
    wire n2684;
    wire n12764;
    wire n2616;
    wire n2683;
    wire n12765;
    wire n2615;
    wire n2682;
    wire n12766;
    wire n2614;
    wire n2681;
    wire n12767;
    wire n2613;
    wire n2680;
    wire n12768;
    wire n2612;
    wire n2679;
    wire n12769;
    wire n2611;
    wire n2678;
    wire n12770;
    wire n12771;
    wire n2610;
    wire bfn_4_24_0_;
    wire n2709;
    wire n2816;
    wire n2883;
    wire n2621;
    wire n2688;
    wire n2720;
    wire n2726;
    wire n2724;
    wire n2720_cascade_;
    wire n2723;
    wire n14136;
    wire n2699;
    wire n2698;
    wire n2820;
    wire n14688_cascade_;
    wire n14690;
    wire n14696;
    wire ENCODER0_B_N;
    wire n2697;
    wire n2630;
    wire n2731;
    wire n2730;
    wire n2729_cascade_;
    wire n13796;
    wire n3094;
    wire n2701;
    wire n2733;
    wire n2733_cascade_;
    wire n2732;
    wire n11936;
    wire n2729;
    wire n2796;
    wire n2819;
    wire n2886;
    wire n2918_cascade_;
    wire n2827;
    wire n2894;
    wire n2926_cascade_;
    wire n14346;
    wire n14336_cascade_;
    wire n14352_cascade_;
    wire n14350;
    wire n2828;
    wire n2895;
    wire n2885;
    wire n2818;
    wire n2881;
    wire n2814;
    wire n12038;
    wire n14358;
    wire n14360_cascade_;
    wire n14366;
    wire n2927;
    wire n2994;
    wire n2909;
    wire n2907;
    wire n14372;
    wire n2929;
    wire n2940_cascade_;
    wire n2996;
    wire n2921;
    wire n2988;
    wire n3083;
    wire n2995;
    wire n2928;
    wire n2997;
    wire n2930;
    wire n3096;
    wire n3029_cascade_;
    wire n2991;
    wire n3019;
    wire n3023_cascade_;
    wire n2922;
    wire n2989;
    wire n3078;
    wire n3075;
    wire n2984;
    wire n2917;
    wire n2931;
    wire n2998;
    wire n3097;
    wire n3030_cascade_;
    wire n3020;
    wire n3087;
    wire n2985;
    wire n2918;
    wire n2911;
    wire n2978;
    wire n2825;
    wire n2892;
    wire n2924;
    wire n2913;
    wire n2980;
    wire n2915;
    wire n2982;
    wire n2912;
    wire n2979;
    wire n2919;
    wire n2986;
    wire n3016;
    wire n3018_cascade_;
    wire n2914;
    wire n2981;
    wire n2908;
    wire n2975;
    wire n3074;
    wire n3007_cascade_;
    wire n2910;
    wire n2977;
    wire \debounce.reg_A_2 ;
    wire \debounce.cnt_next_9__N_424 ;
    wire bfn_5_17_0_;
    wire n12643;
    wire n12644;
    wire n12645;
    wire n12646;
    wire n12647;
    wire n12648;
    wire n12649;
    wire n12650;
    wire bfn_5_18_0_;
    wire n12651;
    wire n12652;
    wire n12653;
    wire n12654;
    wire n12655;
    wire n12656;
    wire n12657;
    wire n12658;
    wire bfn_5_19_0_;
    wire n12659;
    wire n12660;
    wire n12661;
    wire n2315;
    wire n2325;
    wire n2195;
    wire bfn_5_20_0_;
    wire n12662;
    wire n12663;
    wire n12664;
    wire n2297;
    wire n12665;
    wire n2296;
    wire n12666;
    wire n2295;
    wire n12667;
    wire n2294;
    wire n12668;
    wire n12669;
    wire n2293;
    wire bfn_5_21_0_;
    wire n12670;
    wire n12671;
    wire n12672;
    wire n12673;
    wire n2288;
    wire n12674;
    wire n2287;
    wire n12675;
    wire n2286;
    wire n12676;
    wire n12677;
    wire bfn_5_22_0_;
    wire n12678;
    wire n2283;
    wire n12679;
    wire n2282;
    wire n12680;
    wire n12681;
    wire n2313;
    wire n2299;
    wire n2196;
    wire n2198;
    wire n2230;
    wire n2230_cascade_;
    wire n2289;
    wire n2321;
    wire n2331;
    wire n11954;
    wire n311;
    wire n2533;
    wire n2600;
    wire n2532;
    wire n2599;
    wire n2631;
    wire n2633;
    wire n2631_cascade_;
    wire n2632;
    wire n12044;
    wire n2301;
    wire n2333;
    wire bfn_5_25_0_;
    wire n12878;
    wire n12879;
    wire n12880;
    wire n12881;
    wire n12882;
    wire n12883;
    wire n12884;
    wire n12885;
    wire bfn_5_26_0_;
    wire n12886;
    wire n12887;
    wire n12888;
    wire n12889;
    wire n12890;
    wire n12891;
    wire n12892;
    wire n12893;
    wire bfn_5_27_0_;
    wire n12894;
    wire n12895;
    wire n12896;
    wire n12897;
    wire n12898;
    wire n12899;
    wire n12900;
    wire n12901;
    wire bfn_5_28_0_;
    wire n12902;
    wire n12903;
    wire n12904;
    wire n12905;
    wire n12906;
    wire n3180;
    wire n2925;
    wire n2992;
    wire n3099;
    wire n3076;
    wire n2926;
    wire n2993;
    wire n3027;
    wire n3025_cascade_;
    wire n14736;
    wire n3014;
    wire n3081;
    wire n3100;
    wire n3001;
    wire n3033;
    wire n3033_cascade_;
    wire n3032;
    wire n2990;
    wire n3022_cascade_;
    wire n14732;
    wire n3030;
    wire n3029;
    wire n11932;
    wire n13859_cascade_;
    wire n14738;
    wire n2999;
    wire n2932;
    wire n3031;
    wire n3098;
    wire n3031_cascade_;
    wire n2916;
    wire n2983;
    wire n3015;
    wire n3082;
    wire n3015_cascade_;
    wire n3089;
    wire n3022;
    wire n3095;
    wire n3028;
    wire n3127_cascade_;
    wire n3011;
    wire n14744;
    wire n14816;
    wire n14750_cascade_;
    wire n3009;
    wire n3007;
    wire n3008;
    wire n14754_cascade_;
    wire n3006;
    wire n3079;
    wire n3039_cascade_;
    wire n3012;
    wire n14194_cascade_;
    wire n14196;
    wire n3018;
    wire n3085;
    wire n3117_cascade_;
    wire n14198;
    wire n3017;
    wire n3084;
    wire n3025;
    wire n3092;
    wire n3010;
    wire n3077;
    wire n2192;
    wire n2291;
    wire n2224_cascade_;
    wire n2323;
    wire n2193;
    wire n2126_cascade_;
    wire n2292;
    wire n2225_cascade_;
    wire n2324;
    wire n2116_cascade_;
    wire n2183;
    wire n2049_cascade_;
    wire n2186;
    wire n2290;
    wire n2322;
    wire n2116;
    wire n2117_cascade_;
    wire n2148_cascade_;
    wire n2197;
    wire n2229;
    wire n2189;
    wire n2184;
    wire n2117;
    wire n2216;
    wire n2215;
    wire n2214;
    wire n2216_cascade_;
    wire n2298;
    wire n2247_cascade_;
    wire n2330;
    wire n2187;
    wire n2199;
    wire n2285;
    wire n2317;
    wire n2200;
    wire n2191;
    wire n2185;
    wire n2218;
    wire n2219;
    wire n2217_cascade_;
    wire n14598;
    wire n2188;
    wire n2300;
    wire n2332;
    wire n2190;
    wire n2228;
    wire n2224;
    wire n2227;
    wire n14578_cascade_;
    wire n2225;
    wire n2223;
    wire n2222;
    wire n14582_cascade_;
    wire n2221;
    wire n2220;
    wire n14588_cascade_;
    wire n14812;
    wire n14592;
    wire n309;
    wire n17_adj_710_cascade_;
    wire n19_adj_711_cascade_;
    wire n14236;
    wire n14230_cascade_;
    wire n61;
    wire n14268_cascade_;
    wire n14806_cascade_;
    wire n3237_cascade_;
    wire n14228;
    wire n14270;
    wire n14272;
    wire n3173;
    wire n3182;
    wire n3214_cascade_;
    wire n3190;
    wire n3222_cascade_;
    wire n27_adj_713;
    wire n3183;
    wire n3116;
    wire n14794;
    wire n14800;
    wire n2891;
    wire n2824;
    wire n2923;
    wire n3187;
    wire n3189;
    wire n3221_cascade_;
    wire n3175;
    wire n3121;
    wire n3188;
    wire n3191;
    wire n3124;
    wire n3179;
    wire n3113;
    wire n3108;
    wire n14216_cascade_;
    wire n3105;
    wire n14222_cascade_;
    wire n3106;
    wire n3138_cascade_;
    wire n3107;
    wire n3174;
    wire n3201;
    wire n11861;
    wire n3233_cascade_;
    wire n3111;
    wire n3178;
    wire n3023;
    wire n3090;
    wire n3122;
    wire n3181;
    wire n3199;
    wire n3198;
    wire n3115;
    wire n3114;
    wire n14204;
    wire n14210;
    wire n3101;
    wire n3200;
    wire n3133_cascade_;
    wire n3232_cascade_;
    wire n25_adj_712_cascade_;
    wire n37_adj_715;
    wire n14234;
    wire n14238_cascade_;
    wire n14248;
    wire n14250_cascade_;
    wire n3026;
    wire n3093;
    wire n59;
    wire n14252;
    wire n5_adj_703;
    wire n14254_cascade_;
    wire n11926;
    wire n14256_cascade_;
    wire n7_adj_708;
    wire n14264_cascade_;
    wire n14266;
    wire n14258;
    wire n14260_cascade_;
    wire n14262;
    wire n3021;
    wire n3088;
    wire n3120;
    wire bfn_7_17_0_;
    wire n12625;
    wire n2099;
    wire n12626;
    wire n12627;
    wire n2097;
    wire n12628;
    wire n2096;
    wire n12629;
    wire n12630;
    wire n2094;
    wire n12631;
    wire n12632;
    wire n2093;
    wire bfn_7_18_0_;
    wire n12633;
    wire n2091;
    wire n12634;
    wire n12635;
    wire n12636;
    wire n2088;
    wire n12637;
    wire n2087;
    wire n12638;
    wire n12639;
    wire n12640;
    wire n2085;
    wire bfn_7_19_0_;
    wire n2084;
    wire n12641;
    wire n12642;
    wire n2115;
    wire n2095;
    wire n2123;
    wire n2127_cascade_;
    wire n2126;
    wire n2018;
    wire n2092;
    wire n2124;
    wire n2098;
    wire n2130;
    wire n2131;
    wire n2129;
    wire n2130_cascade_;
    wire n2119;
    wire n13775_cascade_;
    wire n14398;
    wire n2090;
    wire n2122;
    wire n2125;
    wire n2122_cascade_;
    wire n2128;
    wire n2120;
    wire n14386_cascade_;
    wire n14384;
    wire n14392;
    wire n2089;
    wire n2121;
    wire n2127;
    wire n2194;
    wire n2226;
    wire n2101;
    wire n2133;
    wire n2133_cascade_;
    wire n11892;
    wire n307;
    wire n2201;
    wire n2233;
    wire n2231;
    wire n2233_cascade_;
    wire n2232;
    wire n11950;
    wire n2086;
    wire n2118;
    wire n308;
    wire n2284;
    wire n2217;
    wire n2316;
    wire n2100;
    wire n2132;
    wire n315;
    wire n15484;
    wire n12034;
    wire bfn_7_23_0_;
    wire n12938;
    wire n15445;
    wire n12939;
    wire n15412;
    wire n12940;
    wire n15378;
    wire n2940;
    wire n12941;
    wire n15346;
    wire n2841;
    wire n12942;
    wire n15310;
    wire n2742;
    wire n12943;
    wire n15852;
    wire n2643;
    wire n12944;
    wire n12945;
    wire n15821;
    wire n2544;
    wire bfn_7_24_0_;
    wire n15791;
    wire n2445;
    wire n12946;
    wire n15765;
    wire n2346;
    wire n12947;
    wire n15739;
    wire n2247;
    wire n12948;
    wire n15714;
    wire n2148;
    wire n12949;
    wire n15689;
    wire n2049;
    wire n12950;
    wire n12951;
    wire n12952;
    wire n12953;
    wire bfn_7_25_0_;
    wire n12954;
    wire n12955;
    wire n12956;
    wire n12957;
    wire n12958;
    wire n12959;
    wire n12960;
    wire n3177;
    wire n3110;
    wire n31_adj_714_cascade_;
    wire n14232;
    wire n3126;
    wire n3193;
    wire n3225_cascade_;
    wire n14776_cascade_;
    wire n14764;
    wire n14780_cascade_;
    wire n3128;
    wire n3195;
    wire n3117;
    wire n3184;
    wire n3119;
    wire n3186;
    wire n3218_cascade_;
    wire n14778;
    wire n12030;
    wire n14786;
    wire n14788;
    wire encoder0_position_scaled_12;
    wire n3194;
    wire n3127;
    wire n3013;
    wire n3080;
    wire n3112;
    wire n3192;
    wire n3125;
    wire n3196;
    wire \debounce.reg_A_0 ;
    wire reg_B_0;
    wire \debounce.reg_A_1 ;
    wire \debounce.n6 ;
    wire n3185;
    wire n3118;
    wire n3197;
    wire n3229_cascade_;
    wire n3237;
    wire n13_adj_709;
    wire n319;
    wire bfn_7_29_0_;
    wire n3301;
    wire n12907;
    wire n3233;
    wire n3300;
    wire n12908;
    wire n3232;
    wire n3299;
    wire n12909;
    wire n3231;
    wire n12910;
    wire n3298;
    wire n3230;
    wire n15097;
    wire n12911;
    wire n3229;
    wire n3296;
    wire n12912;
    wire n3228;
    wire n3295;
    wire n12913;
    wire n12914;
    wire n3227;
    wire n3294;
    wire bfn_7_30_0_;
    wire n3226;
    wire n3293;
    wire n12915;
    wire n3225;
    wire n3292;
    wire n12916;
    wire n3224;
    wire n3291;
    wire n12917;
    wire n3223;
    wire n3290;
    wire n12918;
    wire n3222;
    wire n3289;
    wire n12919;
    wire n3221;
    wire n3288;
    wire n12920;
    wire n3220;
    wire n3287;
    wire n12921;
    wire n12922;
    wire n3219;
    wire n3286;
    wire bfn_7_31_0_;
    wire n3218;
    wire n3285;
    wire n12923;
    wire n3217;
    wire n3284;
    wire n12924;
    wire n3216;
    wire n3283;
    wire n12925;
    wire n3215;
    wire n3282;
    wire n12926;
    wire n3214;
    wire n3281;
    wire n12927;
    wire n3213;
    wire n3280;
    wire n12928;
    wire n3212;
    wire n3279;
    wire n12929;
    wire n12930;
    wire n3211;
    wire n3278;
    wire bfn_7_32_0_;
    wire n3210;
    wire n3277;
    wire n12931;
    wire n3209;
    wire n3276;
    wire n12932;
    wire n3275;
    wire n12933;
    wire n3207;
    wire n3274;
    wire n12934;
    wire n3206;
    wire n3273;
    wire n12935;
    wire n3205;
    wire n3272;
    wire n12936;
    wire n15450;
    wire n3204;
    wire n12937;
    wire n14873;
    wire bfn_9_17_0_;
    wire n12608;
    wire n12609;
    wire n12610;
    wire n12611;
    wire n12612;
    wire n12613;
    wire n12614;
    wire n12615;
    wire bfn_9_18_0_;
    wire n12616;
    wire n12617;
    wire n12618;
    wire n12619;
    wire n12620;
    wire n12621;
    wire n1986;
    wire n12622;
    wire n12623;
    wire bfn_9_19_0_;
    wire n12624;
    wire n2016;
    wire n1993;
    wire n1990;
    wire n1985;
    wire n2017;
    wire n1992;
    wire n1997;
    wire n1987;
    wire n2025;
    wire n2022;
    wire n2024;
    wire n14550_cascade_;
    wire n2029;
    wire n14556_cascade_;
    wire n14558_cascade_;
    wire n2019;
    wire n14564;
    wire n1991;
    wire n2023;
    wire n1994;
    wire n2026;
    wire encoder0_position_0;
    wire bfn_9_22_0_;
    wire \quad_counter0.n13025 ;
    wire \quad_counter0.n13026 ;
    wire \quad_counter0.n13027 ;
    wire encoder0_position_4;
    wire \quad_counter0.n13028 ;
    wire \quad_counter0.n13029 ;
    wire \quad_counter0.n13030 ;
    wire \quad_counter0.n13031 ;
    wire \quad_counter0.n13032 ;
    wire encoder0_position_8;
    wire bfn_9_23_0_;
    wire \quad_counter0.n13033 ;
    wire \quad_counter0.n13034 ;
    wire encoder0_position_11;
    wire \quad_counter0.n13035 ;
    wire encoder0_position_12;
    wire \quad_counter0.n13036 ;
    wire encoder0_position_13;
    wire \quad_counter0.n13037 ;
    wire \quad_counter0.n13038 ;
    wire \quad_counter0.n13039 ;
    wire \quad_counter0.n13040 ;
    wire bfn_9_24_0_;
    wire \quad_counter0.n13041 ;
    wire \quad_counter0.n13042 ;
    wire \quad_counter0.n13043 ;
    wire \quad_counter0.n13044 ;
    wire \quad_counter0.n13045 ;
    wire \quad_counter0.n13046 ;
    wire \quad_counter0.n13047 ;
    wire \quad_counter0.n13048 ;
    wire bfn_9_25_0_;
    wire \quad_counter0.n13049 ;
    wire \quad_counter0.n13050 ;
    wire \quad_counter0.n13051 ;
    wire \quad_counter0.n13052 ;
    wire \quad_counter0.n13053 ;
    wire \quad_counter0.n13054 ;
    wire \quad_counter0.n13055 ;
    wire encoder0_position_scaled_17;
    wire encoder0_position_14;
    wire encoder0_position_scaled_4;
    wire encoder0_position_scaled_5;
    wire encoder0_position_scaled_22;
    wire n3133;
    wire n3132;
    wire n3129;
    wire n3130;
    wire n11930_cascade_;
    wire n3131;
    wire n13819;
    wire \quad_counter0.a_prev_N_543_cascade_ ;
    wire \quad_counter0.direction_N_536 ;
    wire n3024;
    wire n3091;
    wire n3039;
    wire n3123;
    wire ENCODER0_A_N;
    wire \quad_counter0.a_new_0 ;
    wire encoder0_position_scaled_21;
    wire encoder0_position_scaled_19;
    wire n25_adj_605;
    wire pwm_setpoint_23_N_171_0;
    wire bfn_9_30_0_;
    wire n24_adj_604;
    wire pwm_setpoint_23_N_171_1;
    wire n12412;
    wire n23_adj_603;
    wire n12413;
    wire n22_adj_602;
    wire n12414;
    wire n12415;
    wire n12416;
    wire n12417;
    wire n18_adj_598;
    wire n12418;
    wire n12419;
    wire n17_adj_597;
    wire bfn_9_31_0_;
    wire n12420;
    wire n12421;
    wire n14_adj_594;
    wire n12422;
    wire n13_adj_593;
    wire n12423;
    wire n12424;
    wire n12425;
    wire n10_adj_590;
    wire n12426;
    wire n12427;
    wire bfn_9_32_0_;
    wire n12428;
    wire n12429;
    wire n6_adj_586;
    wire n12430;
    wire n12431;
    wire n12432;
    wire n12433;
    wire n12434;
    wire encoder0_position_9;
    wire n310;
    wire n1927;
    wire n1923;
    wire n1926;
    wire n1923_cascade_;
    wire n1924;
    wire n14408;
    wire n1921_cascade_;
    wire n14410;
    wire n1995;
    wire n2027;
    wire n1925;
    wire n1922;
    wire n1989;
    wire n1922_cascade_;
    wire n2021;
    wire n14416;
    wire n14420_cascade_;
    wire n1950_cascade_;
    wire n1998;
    wire n2030;
    wire n15666;
    wire n1917;
    wire n1988;
    wire n1921;
    wire n2020;
    wire n11966;
    wire n1932;
    wire n1932_cascade_;
    wire n1999;
    wire n2031;
    wire n306;
    wire n2031_cascade_;
    wire n11964;
    wire n305;
    wire n2001;
    wire n2033;
    wire n1996;
    wire n2028;
    wire n2000;
    wire n1933;
    wire n1950;
    wire n2032;
    wire n33_adj_654;
    wire n33;
    wire bfn_10_21_0_;
    wire n32_adj_653;
    wire n12968;
    wire n31_adj_652;
    wire n12969;
    wire n12970;
    wire n29_adj_650;
    wire n29;
    wire n12971;
    wire n28_adj_649;
    wire n12972;
    wire n27_adj_648;
    wire n12973;
    wire n26_adj_647;
    wire n12974;
    wire n12975;
    wire n25_adj_646;
    wire n25_adj_551;
    wire bfn_10_22_0_;
    wire n24_adj_645;
    wire n24;
    wire n12976;
    wire n23;
    wire n12977;
    wire n22_adj_643;
    wire n22;
    wire n12978;
    wire n21_adj_642;
    wire n21;
    wire n12979;
    wire n20_adj_641;
    wire n20;
    wire n12980;
    wire n19_adj_640;
    wire n19;
    wire n12981;
    wire n12982;
    wire n12983;
    wire n17_adj_638;
    wire bfn_10_23_0_;
    wire n12984;
    wire n15_adj_636;
    wire n12985;
    wire n12986;
    wire n13_adj_634;
    wire n12987;
    wire n12988;
    wire n12989;
    wire n12990;
    wire n12991;
    wire bfn_10_24_0_;
    wire n12992;
    wire n12993;
    wire n12994;
    wire n12995;
    wire n12996;
    wire n12997;
    wire n12998;
    wire n5_adj_626;
    wire n6_adj_627;
    wire n8_adj_629;
    wire n7_adj_628;
    wire n4_adj_625;
    wire pwm_setpoint_1;
    wire pwm_setpoint_0;
    wire n28;
    wire encoder0_position_5;
    wire n314;
    wire \quad_counter0.b_new_0 ;
    wire encoder0_position_scaled_0;
    wire encoder0_position_scaled_15;
    wire encoder0_position_scaled_13;
    wire n3_adj_624;
    wire encoder0_position_scaled_2;
    wire n4_adj_655;
    wire \quad_counter0.a_prev_N_543 ;
    wire \quad_counter0.b_new_1 ;
    wire \quad_counter0.a_prev ;
    wire \quad_counter0.debounce_cnt ;
    wire \quad_counter0.direction_N_540_cascade_ ;
    wire direction_N_537;
    wire a_new_1;
    wire direction_N_537_cascade_;
    wire b_prev;
    wire n1302;
    wire n29_adj_672_cascade_;
    wire n15233;
    wire n15234;
    wire encoder0_position_scaled_16;
    wire n33_adj_675_cascade_;
    wire n12_adj_592;
    wire pwm_setpoint_23_N_171_16;
    wire pwm_setpoint_23_N_171_2;
    wire pwm_setpoint_23_N_171_14;
    wire pwm_setpoint_14;
    wire n15121;
    wire n15182;
    wire n29_adj_672;
    wire n30_adj_673_cascade_;
    wire n10_adj_659;
    wire n15267;
    wire n20_adj_600;
    wire n16_adj_596;
    wire n15_adj_595;
    wire n21_adj_601;
    wire pwm_setpoint_23_N_171_5;
    wire n19_adj_599;
    wire pwm_setpoint_23_N_171_6;
    wire pwm_setpoint_23_N_171_10;
    wire pwm_setpoint_23_N_171_9;
    wire pwm_setpoint_23_N_171_4;
    wire n7_adj_587;
    wire pwm_setpoint_23_N_171_15;
    wire reg_B_1;
    wire pwm_setpoint_15;
    wire n31_adj_674;
    wire n11_adj_591;
    wire pwm_setpoint_23_N_171_18;
    wire n3_adj_583;
    wire n9_adj_589;
    wire reg_B_2;
    wire n14125;
    wire n14937;
    wire n14936_cascade_;
    wire LED_c;
    wire pwm_setpoint_23_N_171_22;
    wire n1826_cascade_;
    wire n1928;
    wire n14526;
    wire n14530_cascade_;
    wire n1819_cascade_;
    wire n14532;
    wire n1851_cascade_;
    wire n1920;
    wire n1919;
    wire n1930;
    wire n1930_cascade_;
    wire n1929;
    wire n14540;
    wire n1931;
    wire n1918;
    wire n14520;
    wire n14176_cascade_;
    wire n1752_cascade_;
    wire n1851;
    wire n15644;
    wire n1832_cascade_;
    wire n11968;
    wire n1820_cascade_;
    wire n14538;
    wire n30_adj_651;
    wire n26;
    wire encoder0_position_7;
    wire n312;
    wire n31;
    wire encoder0_position_2;
    wire n317;
    wire encoder0_position_10;
    wire n23_adj_644;
    wire encoder0_position_scaled_1;
    wire bfn_11_22_0_;
    wire n12487;
    wire n12488;
    wire n12489;
    wire n12490;
    wire n12491;
    wire n12492;
    wire n901;
    wire n896;
    wire n900;
    wire n899;
    wire n931_cascade_;
    wire n10;
    wire n897;
    wire encoder0_position_25;
    wire n8;
    wire n294;
    wire n14574;
    wire n828;
    wire n828_cascade_;
    wire n12012;
    wire n861;
    wire n861_cascade_;
    wire n898;
    wire n13644_cascade_;
    wire n830;
    wire n7;
    wire n5_adj_676;
    wire n5_adj_676_cascade_;
    wire n13641_cascade_;
    wire n13646_cascade_;
    wire n831;
    wire encoder0_position_28;
    wire n5;
    wire encoder0_position_29;
    wire n4;
    wire n3;
    wire encoder0_position_30;
    wire n13642_cascade_;
    wire n829;
    wire n32;
    wire encoder0_position_1;
    wire n318;
    wire encoder0_position_scaled_14;
    wire n10_adj_606_cascade_;
    wire n15_adj_565_cascade_;
    wire n16_adj_564;
    wire encoder0_position_scaled_10;
    wire pwm_setpoint_23_N_171_3;
    wire encoder0_position_scaled_11;
    wire pwm_setpoint_23_N_171_13;
    wire n15_adj_663_cascade_;
    wire n15125;
    wire encoder0_position_scaled_18;
    wire encoder0_position_scaled_20;
    wire encoder0_position_scaled_23;
    wire n12_adj_661;
    wire pwm_setpoint_23_N_171_7;
    wire pwm_setpoint_16;
    wire pwm_setpoint_7;
    wire n15119;
    wire encoder0_position_scaled_9;
    wire n26_adj_697;
    wire bfn_11_29_0_;
    wire n25_adj_696;
    wire n13087;
    wire n24_adj_695;
    wire n13088;
    wire n23_adj_694;
    wire n13089;
    wire n22_adj_693;
    wire n13090;
    wire n21_adj_692;
    wire n13091;
    wire n20_adj_691;
    wire n13092;
    wire n19_adj_690;
    wire n13093;
    wire n13094;
    wire n18_adj_689;
    wire bfn_11_30_0_;
    wire n17_adj_688;
    wire n13095;
    wire n16_adj_687;
    wire n13096;
    wire n15_adj_686;
    wire n13097;
    wire n14_adj_685;
    wire n13098;
    wire n13_adj_684;
    wire n13099;
    wire n12_adj_683;
    wire n13100;
    wire n11_adj_682;
    wire n13101;
    wire n13102;
    wire n10_adj_681;
    wire bfn_11_31_0_;
    wire n9_adj_680;
    wire n13103;
    wire n8_adj_679;
    wire n13104;
    wire n7_adj_678;
    wire n13105;
    wire n6_adj_677;
    wire n13106;
    wire blink_counter_21;
    wire n13107;
    wire blink_counter_22;
    wire n13108;
    wire blink_counter_23;
    wire n13109;
    wire n13110;
    wire blink_counter_24;
    wire bfn_11_32_0_;
    wire n13111;
    wire blink_counter_25;
    wire pwm_setpoint_23_N_171_19;
    wire n8_adj_588;
    wire n5_adj_585;
    wire n1901;
    wire bfn_12_17_0_;
    wire n1833;
    wire n1900;
    wire n12592;
    wire n1832;
    wire n1899;
    wire n12593;
    wire n1831;
    wire n1898;
    wire n12594;
    wire n1830;
    wire n1897;
    wire n12595;
    wire n1829;
    wire n1896;
    wire n12596;
    wire n1828;
    wire n1895;
    wire n12597;
    wire n1894;
    wire n12598;
    wire n12599;
    wire n1826;
    wire n1893;
    wire bfn_12_18_0_;
    wire n1825;
    wire n1892;
    wire n12600;
    wire n1824;
    wire n1891;
    wire n12601;
    wire n1823;
    wire n1890;
    wire n12602;
    wire n1822;
    wire n1889;
    wire n12603;
    wire n1888;
    wire n12604;
    wire n1820;
    wire n1887;
    wire n12605;
    wire n1819;
    wire n1886;
    wire n12606;
    wire n12607;
    wire bfn_12_19_0_;
    wire n1885;
    wire n1722_cascade_;
    wire n1821;
    wire n1827;
    wire n1752;
    wire n16_adj_637;
    wire n2;
    wire n16;
    wire encoder0_position_17;
    wire n30;
    wire encoder0_position_3;
    wire n316;
    wire n2_adj_623;
    wire encoder0_position_scaled_7;
    wire encoder0_position_23;
    wire n10_adj_631;
    wire n18_adj_639;
    wire n17;
    wire encoder0_position_16;
    wire n18;
    wire encoder0_position_15;
    wire n304;
    wire n15;
    wire encoder0_position_18;
    wire bfn_12_22_0_;
    wire n12493;
    wire n12494;
    wire n12495;
    wire n12496;
    wire n12497;
    wire n12498;
    wire n12499;
    wire n1001;
    wire n927;
    wire n14466_cascade_;
    wire n11940;
    wire n930;
    wire n960_cascade_;
    wire n997;
    wire n929;
    wire n996;
    wire n1028_cascade_;
    wire n998;
    wire n931;
    wire encoder0_position_scaled_8;
    wire n6;
    wire n13641;
    wire n13648_cascade_;
    wire encoder0_position_27;
    wire n832;
    wire n999;
    wire n932;
    wire encoder0_position_26;
    wire n13650;
    wire n833;
    wire encoder0_position_scaled_3;
    wire n293;
    wire n2542;
    wire bfn_12_25_0_;
    wire n292;
    wire n2541;
    wire n12482;
    wire n174;
    wire n2540;
    wire n12483;
    wire n404;
    wire n2539;
    wire n12484;
    wire n403;
    wire n2538;
    wire n12485;
    wire n402;
    wire n12486;
    wire n2537;
    wire encoder0_position_scaled_6;
    wire n3109;
    wire n3176;
    wire n3138;
    wire n3208;
    wire n25_adj_552;
    wire duty_0;
    wire bfn_12_26_0_;
    wire n24_adj_553;
    wire duty_1;
    wire n12459;
    wire n23_adj_554;
    wire duty_2;
    wire n12460;
    wire n22_adj_555;
    wire duty_3;
    wire n12461;
    wire n21_adj_556;
    wire duty_4;
    wire n12462;
    wire n20_adj_557;
    wire duty_5;
    wire n12463;
    wire n19_adj_558;
    wire duty_6;
    wire n12464;
    wire n18_adj_559;
    wire duty_7;
    wire n12465;
    wire n12466;
    wire n17_adj_560;
    wire bfn_12_27_0_;
    wire n16_adj_563;
    wire duty_9;
    wire n12467;
    wire n15_adj_568;
    wire duty_10;
    wire n12468;
    wire n14_adj_569;
    wire n12469;
    wire n13_adj_570;
    wire n12470;
    wire n12_adj_571;
    wire duty_13;
    wire n12471;
    wire n11_adj_572;
    wire duty_14;
    wire n12472;
    wire n10_adj_573;
    wire duty_15;
    wire n12473;
    wire n12474;
    wire n9_adj_574;
    wire duty_16;
    wire bfn_12_28_0_;
    wire n8_adj_575;
    wire n12475;
    wire n7_adj_576;
    wire duty_18;
    wire n12476;
    wire n6_adj_577;
    wire duty_19;
    wire n12477;
    wire n5_adj_578;
    wire n12478;
    wire n4_adj_579;
    wire n12479;
    wire n3_adj_580;
    wire duty_22;
    wire n12480;
    wire n2_adj_581;
    wire n12481;
    wire n35;
    wire n33_adj_675;
    wire n35_cascade_;
    wire n15225;
    wire pwm_setpoint_13;
    wire n27_adj_671;
    wire duty_12;
    wire pwm_setpoint_23_N_171_12;
    wire n37;
    wire pwm_setpoint_18;
    wire n15277;
    wire n6_adj_656;
    wire n15235_cascade_;
    wire n15236_cascade_;
    wire duty_11;
    wire pwm_setpoint_23_N_171_11;
    wire duty_17;
    wire pwm_setpoint_23_N_171_17;
    wire pwm_setpoint_17;
    wire n15278;
    wire n8_adj_657_cascade_;
    wire n15180;
    wire n15219_cascade_;
    wire n24_adj_669;
    wire pwm_setpoint_22;
    wire n15274;
    wire n45;
    wire n15255;
    wire n40_cascade_;
    wire duty_20;
    wire pwm_setpoint_23_N_171_20;
    wire n4_adj_584;
    wire n16_adj_664;
    wire pwm_setpoint_23__N_195;
    wire pwm_setpoint_23_N_171_21;
    wire duty_21;
    wire n1801;
    wire bfn_13_17_0_;
    wire n1800;
    wire n12577;
    wire n1799;
    wire n12578;
    wire n1798;
    wire n12579;
    wire n1797;
    wire n12580;
    wire n1796;
    wire n12581;
    wire n1795;
    wire n12582;
    wire n1794;
    wire n12583;
    wire n12584;
    wire n1793;
    wire bfn_13_18_0_;
    wire n1792;
    wire n12585;
    wire n1791;
    wire n12586;
    wire n1790;
    wire n12587;
    wire n1722;
    wire n1789;
    wire n12588;
    wire n1721;
    wire n1788;
    wire n12589;
    wire n1720;
    wire n1787;
    wire n12590;
    wire n15622;
    wire n12591;
    wire n1818;
    wire bfn_13_19_0_;
    wire n12550;
    wire n12551;
    wire n12552;
    wire n12553;
    wire n12554;
    wire n12555;
    wire n12556;
    wire n12557;
    wire bfn_13_20_0_;
    wire n12558;
    wire n1591;
    wire n12559;
    wire n12560;
    wire n12561;
    wire n12562;
    wire n13;
    wire encoder0_position_20;
    wire n27;
    wire encoder0_position_6;
    wire n313;
    wire n11;
    wire encoder0_position_22;
    wire n11_adj_632;
    wire n9;
    wire n295;
    wire encoder0_position_24;
    wire n9_adj_630;
    wire n933;
    wire n1000;
    wire n1032_cascade_;
    wire n11914_cascade_;
    wire n13716_cascade_;
    wire n1059_cascade_;
    wire n1126_cascade_;
    wire n928;
    wire n960;
    wire n995;
    wire bfn_13_23_0_;
    wire n12500;
    wire n12501;
    wire n12502;
    wire n12503;
    wire n1029;
    wire n1096;
    wire n12504;
    wire n1028;
    wire n1095;
    wire n12505;
    wire n1027;
    wire n1094;
    wire n12506;
    wire n12507;
    wire bfn_13_24_0_;
    wire n1026;
    wire n1093;
    wire n1030;
    wire n1097;
    wire pwm_counter_0;
    wire bfn_13_26_0_;
    wire pwm_counter_1;
    wire \PWM.n13056 ;
    wire \PWM.n13057 ;
    wire \PWM.n13058 ;
    wire \PWM.n13059 ;
    wire \PWM.n13060 ;
    wire \PWM.n13061 ;
    wire \PWM.n13062 ;
    wire \PWM.n13063 ;
    wire bfn_13_27_0_;
    wire \PWM.n13064 ;
    wire \PWM.n13065 ;
    wire \PWM.n13066 ;
    wire \PWM.n13067 ;
    wire \PWM.n13068 ;
    wire \PWM.n13069 ;
    wire \PWM.n13070 ;
    wire \PWM.n13071 ;
    wire bfn_13_28_0_;
    wire \PWM.n13072 ;
    wire \PWM.n13073 ;
    wire \PWM.n13074 ;
    wire \PWM.n13075 ;
    wire \PWM.n13076 ;
    wire \PWM.n13077 ;
    wire \PWM.n13078 ;
    wire \PWM.n13079 ;
    wire bfn_13_29_0_;
    wire \PWM.n13080 ;
    wire \PWM.n13081 ;
    wire \PWM.n13082 ;
    wire \PWM.n13083 ;
    wire \PWM.n13084 ;
    wire \PWM.n13085 ;
    wire \PWM.n13086 ;
    wire n6_adj_717;
    wire pwm_setpoint_5;
    wire pwm_setpoint_6;
    wire pwm_setpoint_10;
    wire pwm_setpoint_11;
    wire pwm_setpoint_12;
    wire pwm_setpoint_20;
    wire n41;
    wire n41_cascade_;
    wire n15265;
    wire n15112;
    wire pwm_setpoint_23;
    wire n15257;
    wire n15108;
    wire pwm_setpoint_21;
    wire pwm_setpoint_19;
    wire n39;
    wire n14910_cascade_;
    wire n1730;
    wire n14514_cascade_;
    wire n1653_cascade_;
    wire n1598;
    wire n1630_adj_617_cascade_;
    wire n1729;
    wire n11902_cascade_;
    wire n13736;
    wire n1599;
    wire n1731;
    wire n1733;
    wire n303;
    wire n1731_cascade_;
    wire n11970;
    wire n1732;
    wire n1590;
    wire n1589;
    wire n1531;
    wire n1531_cascade_;
    wire n1592;
    wire n1533;
    wire n1600;
    wire n1533_cascade_;
    wire n15582;
    wire n14294_cascade_;
    wire n11974;
    wire n1527_cascade_;
    wire n14288;
    wire n14;
    wire n1324_cascade_;
    wire encoder0_position_19;
    wire n14_adj_635;
    wire n1032;
    wire n1099;
    wire n11908_cascade_;
    wire n13708_cascade_;
    wire n1356_cascade_;
    wire n1433_cascade_;
    wire n1031;
    wire n1098;
    wire n296;
    wire n1101;
    wire n1133_cascade_;
    wire n14428;
    wire n12000_cascade_;
    wire n1158_cascade_;
    wire n1232_cascade_;
    wire n12;
    wire encoder0_position_31;
    wire n1100;
    wire n1033;
    wire n1132_cascade_;
    wire n1059;
    wire n15499;
    wire n14470;
    wire encoder0_position_21;
    wire n12_adj_633;
    wire n16_adj_701_cascade_;
    wire n24_adj_561;
    wire n25;
    wire n13932_cascade_;
    wire n14110_cascade_;
    wire n10_adj_567;
    wire n15_adj_702;
    wire n11853;
    wire n23_adj_562;
    wire pwm_setpoint_2;
    wire pwm_setpoint_3;
    wire pwm_counter_2;
    wire pwm_counter_3;
    wire pwm_counter_5;
    wire pwm_counter_7;
    wire pwm_counter_6;
    wire pwm_counter_11;
    wire pwm_counter_10;
    wire pwm_counter_14;
    wire pwm_counter_20;
    wire pwm_counter_16;
    wire pwm_counter_17;
    wire pwm_counter_13;
    wire pwm_counter_23;
    wire pwm_counter_22;
    wire pwm_counter_18;
    wire pwm_counter_15;
    wire pwm_counter_21;
    wire pwm_counter_12;
    wire \PWM.n26_cascade_ ;
    wire \PWM.n28 ;
    wire \PWM.n29_cascade_ ;
    wire \PWM.n27 ;
    wire \PWM.pwm_counter_31__N_407 ;
    wire pwm_counter_19;
    wire \PWM.n13995 ;
    wire \PWM.n17 ;
    wire pwm_counter_24;
    wire pwm_counter_29;
    wire pwm_counter_27;
    wire pwm_counter_26;
    wire pwm_counter_30;
    wire pwm_counter_25;
    wire n12_adj_566_cascade_;
    wire pwm_counter_28;
    wire n5162;
    wire n5162_cascade_;
    wire pwm_counter_31;
    wire n5164;
    wire pwm_setpoint_23_N_171_8;
    wire duty_8;
    wire pwm_setpoint_4;
    wire pwm_counter_4;
    wire n15150;
    wire n11_adj_660;
    wire n9_adj_658_cascade_;
    wire n13_adj_662;
    wire n15_adj_663;
    wire n15205;
    wire n15201_cascade_;
    wire n15261;
    wire pwm_setpoint_8;
    wire pwm_counter_8;
    wire pwm_setpoint_9;
    wire pwm_counter_9;
    wire n21_adj_667;
    wire n19_adj_666;
    wire n17_adj_665;
    wire n9_adj_658;
    wire n43;
    wire n23_adj_668;
    wire n15132_cascade_;
    wire n25_adj_670;
    wire n15110;
    wire commutation_state_7__N_261;
    wire h3;
    wire h1;
    wire h2;
    wire n302;
    wire n1701;
    wire bfn_15_17_0_;
    wire n1700;
    wire n12563;
    wire n1632_adj_619;
    wire n1699;
    wire n12564;
    wire n1631_adj_618;
    wire n1698;
    wire n12565;
    wire n1630_adj_617;
    wire n1697;
    wire n12566;
    wire n12567;
    wire n12568;
    wire n1694;
    wire n12569;
    wire n12570;
    wire bfn_15_18_0_;
    wire n12571;
    wire n1624_adj_611;
    wire n1691;
    wire n12572;
    wire n1623_adj_610;
    wire n1690;
    wire n12573;
    wire n1622_adj_609;
    wire n1689;
    wire n12574;
    wire n1621_adj_608;
    wire n1688;
    wire n12575;
    wire n15603;
    wire n1620_adj_607;
    wire n12576;
    wire n1719;
    wire n1692;
    wire n1523;
    wire n1522;
    wire n1523_cascade_;
    wire n14296;
    wire n1601;
    wire n1554_cascade_;
    wire n301;
    wire n1633_adj_620;
    wire n1532;
    wire n11906;
    wire n14490_cascade_;
    wire n13727;
    wire n14496_cascade_;
    wire n1455_cascade_;
    wire n1525;
    wire n1524;
    wire n299;
    wire n1401;
    wire bfn_15_21_0_;
    wire n1400;
    wire n12527;
    wire n1399;
    wire n12528;
    wire n1331;
    wire n1398;
    wire n12529;
    wire n1330;
    wire n1397;
    wire n12530;
    wire n1396;
    wire n12531;
    wire n12532;
    wire n1394;
    wire n12533;
    wire n12534;
    wire n1393;
    wire bfn_15_22_0_;
    wire n12535;
    wire n1324;
    wire n1391;
    wire n12536;
    wire n15544;
    wire n12537;
    wire n1332;
    wire n1329;
    wire n1333;
    wire n298;
    wire n1301;
    wire bfn_15_23_0_;
    wire n1233;
    wire n1300;
    wire n12517;
    wire n1232;
    wire n1299;
    wire n12518;
    wire n1298;
    wire n12519;
    wire n1297;
    wire n12520;
    wire n12521;
    wire n12522;
    wire n12523;
    wire n12524;
    wire bfn_15_24_0_;
    wire n1292;
    wire n12525;
    wire n12526;
    wire n1323;
    wire bfn_15_25_0_;
    wire encoder0_position_target_0;
    wire n12435;
    wire encoder0_position_target_1;
    wire n12436;
    wire encoder0_position_target_2;
    wire n12437;
    wire encoder0_position_target_3;
    wire n12438;
    wire encoder0_position_target_4;
    wire n12439;
    wire encoder0_position_target_5;
    wire n12440;
    wire encoder0_position_target_6;
    wire n12441;
    wire n12442;
    wire encoder0_position_target_7;
    wire bfn_15_26_0_;
    wire encoder0_position_target_8;
    wire n12443;
    wire encoder0_position_target_9;
    wire n12444;
    wire encoder0_position_target_10;
    wire n12445;
    wire encoder0_position_target_11;
    wire n12446;
    wire encoder0_position_target_12;
    wire n12447;
    wire encoder0_position_target_13;
    wire n12448;
    wire encoder0_position_target_14;
    wire n12449;
    wire n12450;
    wire bfn_15_27_0_;
    wire encoder0_position_target_16;
    wire n12451;
    wire encoder0_position_target_17;
    wire n12452;
    wire encoder0_position_target_18;
    wire n12453;
    wire n12454;
    wire encoder0_position_target_20;
    wire n12455;
    wire n12456;
    wire encoder0_position_target_22;
    wire n12457;
    wire n12458;
    wire bfn_15_28_0_;
    wire n14_adj_718_cascade_;
    wire n10_adj_719;
    wire n5119_cascade_;
    wire n15088;
    wire dti_counter_0;
    wire bfn_15_31_0_;
    wire n15095;
    wire dti_counter_1;
    wire n12961;
    wire n15094;
    wire dti_counter_2;
    wire n12962;
    wire n15093;
    wire dti_counter_3;
    wire n12963;
    wire n15092;
    wire dti_counter_4;
    wire n12964;
    wire n15091;
    wire dti_counter_5;
    wire n12965;
    wire n12966;
    wire n11514;
    wire n15089;
    wire n12967;
    wire dti_counter_7;
    wire n4_adj_716_cascade_;
    wire dti_counter_6;
    wire n15090;
    wire commutation_state_prev_1;
    wire commutation_state_prev_2;
    wire n1693_adj_621;
    wire n1695;
    wire n1727;
    wire n1727_cascade_;
    wire n1726;
    wire n1724;
    wire n1725;
    wire n14166_cascade_;
    wire n1723;
    wire n14172;
    wire n1696;
    wire n1653;
    wire n1728;
    wire n14508;
    wire n1395;
    wire n1427_cascade_;
    wire n1526;
    wire n1526_cascade_;
    wire n1593;
    wire n1625_adj_612;
    wire n1528;
    wire n1595;
    wire n1627_adj_614;
    wire n1527;
    wire n1594;
    wire n1626_adj_613;
    wire n1529;
    wire n1596;
    wire n1628_adj_615;
    wire n1597;
    wire n1554;
    wire n1530;
    wire n1629_adj_616;
    wire n300;
    wire n1501;
    wire bfn_16_19_0_;
    wire n1433;
    wire n1500;
    wire n12538;
    wire n1432;
    wire n1499;
    wire n12539;
    wire n1431;
    wire n1498;
    wire n12540;
    wire n1430;
    wire n1497;
    wire n12541;
    wire n1429;
    wire n1496;
    wire n12542;
    wire n1428;
    wire n1495;
    wire n12543;
    wire n1427;
    wire n1494;
    wire n12544;
    wire n12545;
    wire n1426;
    wire n1493;
    wire bfn_16_20_0_;
    wire n1425;
    wire n1492;
    wire n12546;
    wire n1491;
    wire n12547;
    wire n1423;
    wire n1490;
    wire n12548;
    wire n1422;
    wire n12549;
    wire n1521;
    wire n1455;
    wire n15562;
    wire n1392;
    wire n1356;
    wire n1424;
    wire n1294;
    wire n1295;
    wire n1227;
    wire n14482_cascade_;
    wire n1296;
    wire n1257_cascade_;
    wire n1328;
    wire n1327;
    wire n1328_cascade_;
    wire n1326;
    wire n14282;
    wire n1226;
    wire n1226_cascade_;
    wire n1293;
    wire n1325;
    wire n1229;
    wire n11910;
    wire n1229_cascade_;
    wire n1231;
    wire n13711;
    wire n1257;
    wire n15528;
    wire n1228;
    wire n1230;
    wire n297;
    wire n1201;
    wire bfn_16_23_0_;
    wire n1133;
    wire n1200;
    wire n12508;
    wire n1132;
    wire n1199;
    wire n12509;
    wire n1131;
    wire n1198;
    wire n12510;
    wire n1130;
    wire n1197;
    wire n12511;
    wire n1129;
    wire n1196;
    wire n12512;
    wire n1128;
    wire n1195;
    wire n12513;
    wire n1127;
    wire n1194;
    wire n12514;
    wire n12515;
    wire bfn_16_24_0_;
    wire CONSTANT_ONE_NET;
    wire n15513;
    wire n1125;
    wire n12516;
    wire n1224;
    wire n1126;
    wire n1193;
    wire n1158;
    wire n1225;
    wire n23_adj_700;
    wire n25_adj_698;
    wire direction_N_342_cascade_;
    wire n1693;
    wire direction_N_340;
    wire direction_N_342;
    wire n13661_cascade_;
    wire direction_c;
    wire n22_adj_705_cascade_;
    wire n6_adj_582_cascade_;
    wire n14108;
    wire encoder0_position_target_15;
    wire encoder0_position_target_21;
    wire encoder0_position_target_19;
    wire encoder0_position_target_23;
    wire n24_adj_699;
    wire n16_adj_707;
    wire commutation_state_prev_0;
    wire dti_N_333_cascade_;
    wire n4_adj_716;
    wire n5169;
    wire n1377;
    wire n5119;
    wire n5183_cascade_;
    wire dti;
    wire n20_adj_706_cascade_;
    wire n24_adj_704;
    wire n13187;
    wire sweep_counter_0;
    wire bfn_17_26_0_;
    wire sweep_counter_1;
    wire n12999;
    wire sweep_counter_2;
    wire n13000;
    wire sweep_counter_3;
    wire n13001;
    wire sweep_counter_4;
    wire n13002;
    wire sweep_counter_5;
    wire n13003;
    wire sweep_counter_6;
    wire n13004;
    wire sweep_counter_7;
    wire n13005;
    wire n13006;
    wire sweep_counter_8;
    wire bfn_17_27_0_;
    wire sweep_counter_9;
    wire n13007;
    wire sweep_counter_10;
    wire n13008;
    wire sweep_counter_11;
    wire n13009;
    wire sweep_counter_12;
    wire n13010;
    wire sweep_counter_13;
    wire n13011;
    wire sweep_counter_14;
    wire n13012;
    wire sweep_counter_15;
    wire n13013;
    wire n13014;
    wire sweep_counter_16;
    wire bfn_17_28_0_;
    wire n13015;
    wire sweep_counter_17;
    wire n5197;
    wire duty_23;
    wire INLB_c_0;
    wire INLA_c_0;
    wire commutation_state_0;
    wire commutation_state_1;
    wire commutation_state_2;
    wire dir;
    wire INLC_c_0;
    wire CLK_N;
    wire n5183;
    wire n5235;
    wire GHB;
    wire INHB_c_0;
    wire GHC;
    wire INHC_c_0;
    wire pwm_out;
    wire GHA;
    wire INHA_c_0;
    wire _gnd_net_;

    defparam CS_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_CLK_pad_iopad (
            .OE(N__56344),
            .DIN(N__56343),
            .DOUT(N__56342),
            .PACKAGEPIN(CS_CLK));
    defparam CS_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_CLK_pad_preio (
            .PADOEN(N__56344),
            .PADOUT(N__56343),
            .PADIN(N__56342),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_pad_iopad (
            .OE(N__56335),
            .DIN(N__56334),
            .DOUT(N__56333),
            .PACKAGEPIN(CS));
    defparam CS_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_pad_preio (
            .PADOEN(N__56335),
            .PADOUT(N__56334),
            .PADIN(N__56333),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam DE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DE_pad_iopad.PULLUP=1'b0;
    IO_PAD DE_pad_iopad (
            .OE(N__56326),
            .DIN(N__56325),
            .DOUT(N__56324),
            .PACKAGEPIN(DE));
    defparam DE_pad_preio.PIN_TYPE=6'b011001;
    defparam DE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DE_pad_preio (
            .PADOEN(N__56326),
            .PADOUT(N__56325),
            .PADIN(N__56324),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ENCODER0_A_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ENCODER0_A_pad_iopad.PULLUP=1'b0;
    IO_PAD ENCODER0_A_pad_iopad (
            .OE(N__56317),
            .DIN(N__56316),
            .DOUT(N__56315),
            .PACKAGEPIN(ENCODER0_A));
    defparam ENCODER0_A_pad_preio.PIN_TYPE=6'b000001;
    defparam ENCODER0_A_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ENCODER0_A_pad_preio (
            .PADOEN(N__56317),
            .PADOUT(N__56316),
            .PADIN(N__56315),
            .CLOCKENABLE(),
            .DIN0(ENCODER0_A_N),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ENCODER0_B_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ENCODER0_B_pad_iopad.PULLUP=1'b0;
    IO_PAD ENCODER0_B_pad_iopad (
            .OE(N__56308),
            .DIN(N__56307),
            .DOUT(N__56306),
            .PACKAGEPIN(ENCODER0_B));
    defparam ENCODER0_B_pad_preio.PIN_TYPE=6'b000001;
    defparam ENCODER0_B_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ENCODER0_B_pad_preio (
            .PADOEN(N__56308),
            .PADOUT(N__56307),
            .PADIN(N__56306),
            .CLOCKENABLE(),
            .DIN0(ENCODER0_B_N),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHA_pad_iopad.PULLUP=1'b0;
    IO_PAD INHA_pad_iopad (
            .OE(N__56299),
            .DIN(N__56298),
            .DOUT(N__56297),
            .PACKAGEPIN(INHA));
    defparam INHA_pad_preio.PIN_TYPE=6'b011001;
    defparam INHA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHA_pad_preio (
            .PADOEN(N__56299),
            .PADOUT(N__56298),
            .PADIN(N__56297),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55479),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHB_pad_iopad.PULLUP=1'b0;
    IO_PAD INHB_pad_iopad (
            .OE(N__56290),
            .DIN(N__56289),
            .DOUT(N__56288),
            .PACKAGEPIN(INHB));
    defparam INHB_pad_preio.PIN_TYPE=6'b011001;
    defparam INHB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHB_pad_preio (
            .PADOEN(N__56290),
            .PADOUT(N__56289),
            .PADIN(N__56288),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55548),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHC_pad_iopad.PULLUP=1'b0;
    IO_PAD INHC_pad_iopad (
            .OE(N__56281),
            .DIN(N__56280),
            .DOUT(N__56279),
            .PACKAGEPIN(INHC));
    defparam INHC_pad_preio.PIN_TYPE=6'b011001;
    defparam INHC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHC_pad_preio (
            .PADOEN(N__56281),
            .PADOUT(N__56280),
            .PADIN(N__56279),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55527),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLA_pad_iopad.PULLUP=1'b0;
    IO_PAD INLA_pad_iopad (
            .OE(N__56272),
            .DIN(N__56271),
            .DOUT(N__56270),
            .PACKAGEPIN(INLA));
    defparam INLA_pad_preio.PIN_TYPE=6'b011001;
    defparam INLA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLA_pad_preio (
            .PADOEN(N__56272),
            .PADOUT(N__56271),
            .PADIN(N__56270),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56163),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLB_pad_iopad.PULLUP=1'b0;
    IO_PAD INLB_pad_iopad (
            .OE(N__56263),
            .DIN(N__56262),
            .DOUT(N__56261),
            .PACKAGEPIN(INLB));
    defparam INLB_pad_preio.PIN_TYPE=6'b011001;
    defparam INLB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLB_pad_preio (
            .PADOEN(N__56263),
            .PADOUT(N__56262),
            .PADIN(N__56261),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55191),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLC_pad_iopad.PULLUP=1'b0;
    IO_PAD INLC_pad_iopad (
            .OE(N__56254),
            .DIN(N__56253),
            .DOUT(N__56252),
            .PACKAGEPIN(INLC));
    defparam INLC_pad_preio.PIN_TYPE=6'b011001;
    defparam INLC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLC_pad_preio (
            .PADOEN(N__56254),
            .PADOUT(N__56253),
            .PADIN(N__56252),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55854),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__56245),
            .DIN(N__56244),
            .DOUT(N__56243),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__56245),
            .PADOUT(N__56244),
            .PADIN(N__56243),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__39489),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__56236),
            .DIN(N__56235),
            .DOUT(N__56234),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__56236),
            .PADOUT(N__56235),
            .PADIN(N__56234),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TX_pad_iopad.PULLUP=1'b0;
    IO_PAD TX_pad_iopad (
            .OE(N__56227),
            .DIN(N__56226),
            .DOUT(N__56225),
            .PACKAGEPIN(TX));
    defparam TX_pad_preio.PIN_TYPE=6'b011001;
    defparam TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TX_pad_preio (
            .PADOEN(N__56227),
            .PADOUT(N__56226),
            .PADIN(N__56225),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__56218),
            .DIN(N__56217),
            .DOUT(N__56216),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__56218),
            .PADOUT(N__56217),
            .PADIN(N__56216),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__56209),
            .DIN(N__56208),
            .DOUT(N__56207),
            .PACKAGEPIN(HALL1));
    defparam hall1_input_preio.PIN_TYPE=6'b000000;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__56209),
            .PADOUT(N__56208),
            .PADIN(N__56207),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_2 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__55776),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__56200),
            .DIN(N__56199),
            .DOUT(N__56198),
            .PACKAGEPIN(HALL2));
    defparam hall2_input_preio.PIN_TYPE=6'b000000;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__56200),
            .PADOUT(N__56199),
            .PADIN(N__56198),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_1 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__55774),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__56191),
            .DIN(N__56190),
            .DOUT(N__56189),
            .PACKAGEPIN(HALL3));
    defparam hall3_input_preio.PIN_TYPE=6'b000000;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__56191),
            .PADOUT(N__56190),
            .PADIN(N__56189),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_0 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__55774),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__56182),
            .DIN(N__56181),
            .DOUT(N__56180),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__56182),
            .PADOUT(N__56181),
            .PADIN(N__56180),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__13316 (
            .O(N__56163),
            .I(N__56160));
    LocalMux I__13315 (
            .O(N__56160),
            .I(N__56157));
    IoSpan4Mux I__13314 (
            .O(N__56157),
            .I(N__56154));
    Span4Mux_s0_v I__13313 (
            .O(N__56154),
            .I(N__56151));
    Odrv4 I__13312 (
            .O(N__56151),
            .I(INLA_c_0));
    InMux I__13311 (
            .O(N__56148),
            .I(N__56140));
    InMux I__13310 (
            .O(N__56147),
            .I(N__56137));
    InMux I__13309 (
            .O(N__56146),
            .I(N__56132));
    InMux I__13308 (
            .O(N__56145),
            .I(N__56132));
    InMux I__13307 (
            .O(N__56144),
            .I(N__56127));
    InMux I__13306 (
            .O(N__56143),
            .I(N__56127));
    LocalMux I__13305 (
            .O(N__56140),
            .I(N__56119));
    LocalMux I__13304 (
            .O(N__56137),
            .I(N__56119));
    LocalMux I__13303 (
            .O(N__56132),
            .I(N__56113));
    LocalMux I__13302 (
            .O(N__56127),
            .I(N__56113));
    InMux I__13301 (
            .O(N__56126),
            .I(N__56107));
    InMux I__13300 (
            .O(N__56125),
            .I(N__56102));
    InMux I__13299 (
            .O(N__56124),
            .I(N__56102));
    Span4Mux_v I__13298 (
            .O(N__56119),
            .I(N__56096));
    InMux I__13297 (
            .O(N__56118),
            .I(N__56093));
    Span4Mux_s2_v I__13296 (
            .O(N__56113),
            .I(N__56090));
    InMux I__13295 (
            .O(N__56112),
            .I(N__56083));
    InMux I__13294 (
            .O(N__56111),
            .I(N__56083));
    InMux I__13293 (
            .O(N__56110),
            .I(N__56083));
    LocalMux I__13292 (
            .O(N__56107),
            .I(N__56080));
    LocalMux I__13291 (
            .O(N__56102),
            .I(N__56077));
    InMux I__13290 (
            .O(N__56101),
            .I(N__56074));
    InMux I__13289 (
            .O(N__56100),
            .I(N__56069));
    InMux I__13288 (
            .O(N__56099),
            .I(N__56069));
    Span4Mux_h I__13287 (
            .O(N__56096),
            .I(N__56064));
    LocalMux I__13286 (
            .O(N__56093),
            .I(N__56064));
    Span4Mux_h I__13285 (
            .O(N__56090),
            .I(N__56055));
    LocalMux I__13284 (
            .O(N__56083),
            .I(N__56055));
    Span4Mux_h I__13283 (
            .O(N__56080),
            .I(N__56055));
    Span4Mux_s2_v I__13282 (
            .O(N__56077),
            .I(N__56055));
    LocalMux I__13281 (
            .O(N__56074),
            .I(commutation_state_0));
    LocalMux I__13280 (
            .O(N__56069),
            .I(commutation_state_0));
    Odrv4 I__13279 (
            .O(N__56064),
            .I(commutation_state_0));
    Odrv4 I__13278 (
            .O(N__56055),
            .I(commutation_state_0));
    CascadeMux I__13277 (
            .O(N__56046),
            .I(N__56040));
    CascadeMux I__13276 (
            .O(N__56045),
            .I(N__56037));
    InMux I__13275 (
            .O(N__56044),
            .I(N__56031));
    InMux I__13274 (
            .O(N__56043),
            .I(N__56031));
    InMux I__13273 (
            .O(N__56040),
            .I(N__56024));
    InMux I__13272 (
            .O(N__56037),
            .I(N__56024));
    InMux I__13271 (
            .O(N__56036),
            .I(N__56021));
    LocalMux I__13270 (
            .O(N__56031),
            .I(N__56018));
    InMux I__13269 (
            .O(N__56030),
            .I(N__56014));
    CascadeMux I__13268 (
            .O(N__56029),
            .I(N__56010));
    LocalMux I__13267 (
            .O(N__56024),
            .I(N__56003));
    LocalMux I__13266 (
            .O(N__56021),
            .I(N__56003));
    Span4Mux_s1_v I__13265 (
            .O(N__56018),
            .I(N__56003));
    CascadeMux I__13264 (
            .O(N__56017),
            .I(N__55999));
    LocalMux I__13263 (
            .O(N__56014),
            .I(N__55996));
    InMux I__13262 (
            .O(N__56013),
            .I(N__55993));
    InMux I__13261 (
            .O(N__56010),
            .I(N__55990));
    Span4Mux_h I__13260 (
            .O(N__56003),
            .I(N__55987));
    InMux I__13259 (
            .O(N__56002),
            .I(N__55982));
    InMux I__13258 (
            .O(N__55999),
            .I(N__55982));
    Span4Mux_s1_v I__13257 (
            .O(N__55996),
            .I(N__55977));
    LocalMux I__13256 (
            .O(N__55993),
            .I(N__55977));
    LocalMux I__13255 (
            .O(N__55990),
            .I(commutation_state_1));
    Odrv4 I__13254 (
            .O(N__55987),
            .I(commutation_state_1));
    LocalMux I__13253 (
            .O(N__55982),
            .I(commutation_state_1));
    Odrv4 I__13252 (
            .O(N__55977),
            .I(commutation_state_1));
    CascadeMux I__13251 (
            .O(N__55968),
            .I(N__55965));
    InMux I__13250 (
            .O(N__55965),
            .I(N__55957));
    InMux I__13249 (
            .O(N__55964),
            .I(N__55952));
    InMux I__13248 (
            .O(N__55963),
            .I(N__55952));
    CascadeMux I__13247 (
            .O(N__55962),
            .I(N__55947));
    CascadeMux I__13246 (
            .O(N__55961),
            .I(N__55944));
    CascadeMux I__13245 (
            .O(N__55960),
            .I(N__55941));
    LocalMux I__13244 (
            .O(N__55957),
            .I(N__55936));
    LocalMux I__13243 (
            .O(N__55952),
            .I(N__55936));
    InMux I__13242 (
            .O(N__55951),
            .I(N__55933));
    CascadeMux I__13241 (
            .O(N__55950),
            .I(N__55930));
    InMux I__13240 (
            .O(N__55947),
            .I(N__55927));
    InMux I__13239 (
            .O(N__55944),
            .I(N__55922));
    InMux I__13238 (
            .O(N__55941),
            .I(N__55922));
    Span4Mux_h I__13237 (
            .O(N__55936),
            .I(N__55915));
    LocalMux I__13236 (
            .O(N__55933),
            .I(N__55915));
    InMux I__13235 (
            .O(N__55930),
            .I(N__55912));
    LocalMux I__13234 (
            .O(N__55927),
            .I(N__55907));
    LocalMux I__13233 (
            .O(N__55922),
            .I(N__55907));
    InMux I__13232 (
            .O(N__55921),
            .I(N__55902));
    InMux I__13231 (
            .O(N__55920),
            .I(N__55902));
    Span4Mux_h I__13230 (
            .O(N__55915),
            .I(N__55899));
    LocalMux I__13229 (
            .O(N__55912),
            .I(commutation_state_2));
    Odrv12 I__13228 (
            .O(N__55907),
            .I(commutation_state_2));
    LocalMux I__13227 (
            .O(N__55902),
            .I(commutation_state_2));
    Odrv4 I__13226 (
            .O(N__55899),
            .I(commutation_state_2));
    InMux I__13225 (
            .O(N__55890),
            .I(N__55884));
    InMux I__13224 (
            .O(N__55889),
            .I(N__55884));
    LocalMux I__13223 (
            .O(N__55884),
            .I(N__55878));
    InMux I__13222 (
            .O(N__55883),
            .I(N__55873));
    InMux I__13221 (
            .O(N__55882),
            .I(N__55873));
    InMux I__13220 (
            .O(N__55881),
            .I(N__55869));
    Span4Mux_v I__13219 (
            .O(N__55878),
            .I(N__55864));
    LocalMux I__13218 (
            .O(N__55873),
            .I(N__55864));
    InMux I__13217 (
            .O(N__55872),
            .I(N__55861));
    LocalMux I__13216 (
            .O(N__55869),
            .I(dir));
    Odrv4 I__13215 (
            .O(N__55864),
            .I(dir));
    LocalMux I__13214 (
            .O(N__55861),
            .I(dir));
    IoInMux I__13213 (
            .O(N__55854),
            .I(N__55851));
    LocalMux I__13212 (
            .O(N__55851),
            .I(N__55848));
    Span4Mux_s0_v I__13211 (
            .O(N__55848),
            .I(N__55845));
    Span4Mux_h I__13210 (
            .O(N__55845),
            .I(N__55842));
    Span4Mux_h I__13209 (
            .O(N__55842),
            .I(N__55839));
    Odrv4 I__13208 (
            .O(N__55839),
            .I(INLC_c_0));
    ClkMux I__13207 (
            .O(N__55836),
            .I(N__55644));
    ClkMux I__13206 (
            .O(N__55835),
            .I(N__55644));
    ClkMux I__13205 (
            .O(N__55834),
            .I(N__55644));
    ClkMux I__13204 (
            .O(N__55833),
            .I(N__55644));
    ClkMux I__13203 (
            .O(N__55832),
            .I(N__55644));
    ClkMux I__13202 (
            .O(N__55831),
            .I(N__55644));
    ClkMux I__13201 (
            .O(N__55830),
            .I(N__55644));
    ClkMux I__13200 (
            .O(N__55829),
            .I(N__55644));
    ClkMux I__13199 (
            .O(N__55828),
            .I(N__55644));
    ClkMux I__13198 (
            .O(N__55827),
            .I(N__55644));
    ClkMux I__13197 (
            .O(N__55826),
            .I(N__55644));
    ClkMux I__13196 (
            .O(N__55825),
            .I(N__55644));
    ClkMux I__13195 (
            .O(N__55824),
            .I(N__55644));
    ClkMux I__13194 (
            .O(N__55823),
            .I(N__55644));
    ClkMux I__13193 (
            .O(N__55822),
            .I(N__55644));
    ClkMux I__13192 (
            .O(N__55821),
            .I(N__55644));
    ClkMux I__13191 (
            .O(N__55820),
            .I(N__55644));
    ClkMux I__13190 (
            .O(N__55819),
            .I(N__55644));
    ClkMux I__13189 (
            .O(N__55818),
            .I(N__55644));
    ClkMux I__13188 (
            .O(N__55817),
            .I(N__55644));
    ClkMux I__13187 (
            .O(N__55816),
            .I(N__55644));
    ClkMux I__13186 (
            .O(N__55815),
            .I(N__55644));
    ClkMux I__13185 (
            .O(N__55814),
            .I(N__55644));
    ClkMux I__13184 (
            .O(N__55813),
            .I(N__55644));
    ClkMux I__13183 (
            .O(N__55812),
            .I(N__55644));
    ClkMux I__13182 (
            .O(N__55811),
            .I(N__55644));
    ClkMux I__13181 (
            .O(N__55810),
            .I(N__55644));
    ClkMux I__13180 (
            .O(N__55809),
            .I(N__55644));
    ClkMux I__13179 (
            .O(N__55808),
            .I(N__55644));
    ClkMux I__13178 (
            .O(N__55807),
            .I(N__55644));
    ClkMux I__13177 (
            .O(N__55806),
            .I(N__55644));
    ClkMux I__13176 (
            .O(N__55805),
            .I(N__55644));
    ClkMux I__13175 (
            .O(N__55804),
            .I(N__55644));
    ClkMux I__13174 (
            .O(N__55803),
            .I(N__55644));
    ClkMux I__13173 (
            .O(N__55802),
            .I(N__55644));
    ClkMux I__13172 (
            .O(N__55801),
            .I(N__55644));
    ClkMux I__13171 (
            .O(N__55800),
            .I(N__55644));
    ClkMux I__13170 (
            .O(N__55799),
            .I(N__55644));
    ClkMux I__13169 (
            .O(N__55798),
            .I(N__55644));
    ClkMux I__13168 (
            .O(N__55797),
            .I(N__55644));
    ClkMux I__13167 (
            .O(N__55796),
            .I(N__55644));
    ClkMux I__13166 (
            .O(N__55795),
            .I(N__55644));
    ClkMux I__13165 (
            .O(N__55794),
            .I(N__55644));
    ClkMux I__13164 (
            .O(N__55793),
            .I(N__55644));
    ClkMux I__13163 (
            .O(N__55792),
            .I(N__55644));
    ClkMux I__13162 (
            .O(N__55791),
            .I(N__55644));
    ClkMux I__13161 (
            .O(N__55790),
            .I(N__55644));
    ClkMux I__13160 (
            .O(N__55789),
            .I(N__55644));
    ClkMux I__13159 (
            .O(N__55788),
            .I(N__55644));
    ClkMux I__13158 (
            .O(N__55787),
            .I(N__55644));
    ClkMux I__13157 (
            .O(N__55786),
            .I(N__55644));
    ClkMux I__13156 (
            .O(N__55785),
            .I(N__55644));
    ClkMux I__13155 (
            .O(N__55784),
            .I(N__55644));
    ClkMux I__13154 (
            .O(N__55783),
            .I(N__55644));
    ClkMux I__13153 (
            .O(N__55782),
            .I(N__55644));
    ClkMux I__13152 (
            .O(N__55781),
            .I(N__55644));
    ClkMux I__13151 (
            .O(N__55780),
            .I(N__55644));
    ClkMux I__13150 (
            .O(N__55779),
            .I(N__55644));
    ClkMux I__13149 (
            .O(N__55778),
            .I(N__55644));
    ClkMux I__13148 (
            .O(N__55777),
            .I(N__55644));
    ClkMux I__13147 (
            .O(N__55776),
            .I(N__55644));
    ClkMux I__13146 (
            .O(N__55775),
            .I(N__55644));
    ClkMux I__13145 (
            .O(N__55774),
            .I(N__55644));
    ClkMux I__13144 (
            .O(N__55773),
            .I(N__55644));
    GlobalMux I__13143 (
            .O(N__55644),
            .I(N__55641));
    gio2CtrlBuf I__13142 (
            .O(N__55641),
            .I(CLK_N));
    CEMux I__13141 (
            .O(N__55638),
            .I(N__55634));
    CEMux I__13140 (
            .O(N__55637),
            .I(N__55630));
    LocalMux I__13139 (
            .O(N__55634),
            .I(N__55626));
    CEMux I__13138 (
            .O(N__55633),
            .I(N__55623));
    LocalMux I__13137 (
            .O(N__55630),
            .I(N__55620));
    CEMux I__13136 (
            .O(N__55629),
            .I(N__55617));
    Span4Mux_s1_v I__13135 (
            .O(N__55626),
            .I(N__55612));
    LocalMux I__13134 (
            .O(N__55623),
            .I(N__55612));
    Span4Mux_s1_v I__13133 (
            .O(N__55620),
            .I(N__55609));
    LocalMux I__13132 (
            .O(N__55617),
            .I(N__55606));
    Span4Mux_v I__13131 (
            .O(N__55612),
            .I(N__55603));
    Odrv4 I__13130 (
            .O(N__55609),
            .I(n5183));
    Odrv12 I__13129 (
            .O(N__55606),
            .I(n5183));
    Odrv4 I__13128 (
            .O(N__55603),
            .I(n5183));
    SRMux I__13127 (
            .O(N__55596),
            .I(N__55593));
    LocalMux I__13126 (
            .O(N__55593),
            .I(N__55587));
    SRMux I__13125 (
            .O(N__55592),
            .I(N__55584));
    SRMux I__13124 (
            .O(N__55591),
            .I(N__55581));
    SRMux I__13123 (
            .O(N__55590),
            .I(N__55578));
    Span4Mux_h I__13122 (
            .O(N__55587),
            .I(N__55573));
    LocalMux I__13121 (
            .O(N__55584),
            .I(N__55573));
    LocalMux I__13120 (
            .O(N__55581),
            .I(N__55568));
    LocalMux I__13119 (
            .O(N__55578),
            .I(N__55568));
    Span4Mux_h I__13118 (
            .O(N__55573),
            .I(N__55565));
    Span4Mux_s1_v I__13117 (
            .O(N__55568),
            .I(N__55560));
    Span4Mux_s1_v I__13116 (
            .O(N__55565),
            .I(N__55560));
    Odrv4 I__13115 (
            .O(N__55560),
            .I(n5235));
    InMux I__13114 (
            .O(N__55557),
            .I(N__55554));
    LocalMux I__13113 (
            .O(N__55554),
            .I(N__55551));
    Odrv12 I__13112 (
            .O(N__55551),
            .I(GHB));
    IoInMux I__13111 (
            .O(N__55548),
            .I(N__55545));
    LocalMux I__13110 (
            .O(N__55545),
            .I(N__55542));
    Span4Mux_s1_v I__13109 (
            .O(N__55542),
            .I(N__55539));
    Span4Mux_h I__13108 (
            .O(N__55539),
            .I(N__55536));
    Odrv4 I__13107 (
            .O(N__55536),
            .I(INHB_c_0));
    InMux I__13106 (
            .O(N__55533),
            .I(N__55530));
    LocalMux I__13105 (
            .O(N__55530),
            .I(GHC));
    IoInMux I__13104 (
            .O(N__55527),
            .I(N__55524));
    LocalMux I__13103 (
            .O(N__55524),
            .I(N__55521));
    Span4Mux_s1_v I__13102 (
            .O(N__55521),
            .I(N__55518));
    Span4Mux_h I__13101 (
            .O(N__55518),
            .I(N__55515));
    Odrv4 I__13100 (
            .O(N__55515),
            .I(INHC_c_0));
    InMux I__13099 (
            .O(N__55512),
            .I(N__55509));
    LocalMux I__13098 (
            .O(N__55509),
            .I(N__55506));
    Span4Mux_s1_v I__13097 (
            .O(N__55506),
            .I(N__55501));
    InMux I__13096 (
            .O(N__55505),
            .I(N__55496));
    InMux I__13095 (
            .O(N__55504),
            .I(N__55496));
    Sp12to4 I__13094 (
            .O(N__55501),
            .I(N__55491));
    LocalMux I__13093 (
            .O(N__55496),
            .I(N__55491));
    Odrv12 I__13092 (
            .O(N__55491),
            .I(pwm_out));
    InMux I__13091 (
            .O(N__55488),
            .I(N__55485));
    LocalMux I__13090 (
            .O(N__55485),
            .I(N__55482));
    Odrv12 I__13089 (
            .O(N__55482),
            .I(GHA));
    IoInMux I__13088 (
            .O(N__55479),
            .I(N__55476));
    LocalMux I__13087 (
            .O(N__55476),
            .I(N__55473));
    Span4Mux_s0_v I__13086 (
            .O(N__55473),
            .I(N__55470));
    Odrv4 I__13085 (
            .O(N__55470),
            .I(INHA_c_0));
    InMux I__13084 (
            .O(N__55467),
            .I(N__55463));
    InMux I__13083 (
            .O(N__55466),
            .I(N__55460));
    LocalMux I__13082 (
            .O(N__55463),
            .I(sweep_counter_14));
    LocalMux I__13081 (
            .O(N__55460),
            .I(sweep_counter_14));
    InMux I__13080 (
            .O(N__55455),
            .I(n13012));
    InMux I__13079 (
            .O(N__55452),
            .I(N__55448));
    InMux I__13078 (
            .O(N__55451),
            .I(N__55445));
    LocalMux I__13077 (
            .O(N__55448),
            .I(sweep_counter_15));
    LocalMux I__13076 (
            .O(N__55445),
            .I(sweep_counter_15));
    InMux I__13075 (
            .O(N__55440),
            .I(n13013));
    InMux I__13074 (
            .O(N__55437),
            .I(N__55433));
    InMux I__13073 (
            .O(N__55436),
            .I(N__55430));
    LocalMux I__13072 (
            .O(N__55433),
            .I(N__55427));
    LocalMux I__13071 (
            .O(N__55430),
            .I(sweep_counter_16));
    Odrv4 I__13070 (
            .O(N__55427),
            .I(sweep_counter_16));
    InMux I__13069 (
            .O(N__55422),
            .I(bfn_17_28_0_));
    InMux I__13068 (
            .O(N__55419),
            .I(n13015));
    InMux I__13067 (
            .O(N__55416),
            .I(N__55412));
    InMux I__13066 (
            .O(N__55415),
            .I(N__55409));
    LocalMux I__13065 (
            .O(N__55412),
            .I(sweep_counter_17));
    LocalMux I__13064 (
            .O(N__55409),
            .I(sweep_counter_17));
    CEMux I__13063 (
            .O(N__55404),
            .I(N__55396));
    SRMux I__13062 (
            .O(N__55403),
            .I(N__55393));
    CEMux I__13061 (
            .O(N__55402),
            .I(N__55390));
    SRMux I__13060 (
            .O(N__55401),
            .I(N__55386));
    SRMux I__13059 (
            .O(N__55400),
            .I(N__55383));
    CEMux I__13058 (
            .O(N__55399),
            .I(N__55380));
    LocalMux I__13057 (
            .O(N__55396),
            .I(N__55377));
    LocalMux I__13056 (
            .O(N__55393),
            .I(N__55374));
    LocalMux I__13055 (
            .O(N__55390),
            .I(N__55371));
    CEMux I__13054 (
            .O(N__55389),
            .I(N__55368));
    LocalMux I__13053 (
            .O(N__55386),
            .I(N__55365));
    LocalMux I__13052 (
            .O(N__55383),
            .I(N__55362));
    LocalMux I__13051 (
            .O(N__55380),
            .I(N__55359));
    Span4Mux_h I__13050 (
            .O(N__55377),
            .I(N__55354));
    Span4Mux_h I__13049 (
            .O(N__55374),
            .I(N__55354));
    Span4Mux_h I__13048 (
            .O(N__55371),
            .I(N__55347));
    LocalMux I__13047 (
            .O(N__55368),
            .I(N__55347));
    Span4Mux_h I__13046 (
            .O(N__55365),
            .I(N__55347));
    Span4Mux_h I__13045 (
            .O(N__55362),
            .I(N__55344));
    Odrv4 I__13044 (
            .O(N__55359),
            .I(n5197));
    Odrv4 I__13043 (
            .O(N__55354),
            .I(n5197));
    Odrv4 I__13042 (
            .O(N__55347),
            .I(n5197));
    Odrv4 I__13041 (
            .O(N__55344),
            .I(n5197));
    InMux I__13040 (
            .O(N__55335),
            .I(N__55319));
    InMux I__13039 (
            .O(N__55334),
            .I(N__55316));
    InMux I__13038 (
            .O(N__55333),
            .I(N__55311));
    InMux I__13037 (
            .O(N__55332),
            .I(N__55311));
    InMux I__13036 (
            .O(N__55331),
            .I(N__55301));
    InMux I__13035 (
            .O(N__55330),
            .I(N__55301));
    InMux I__13034 (
            .O(N__55329),
            .I(N__55298));
    InMux I__13033 (
            .O(N__55328),
            .I(N__55291));
    InMux I__13032 (
            .O(N__55327),
            .I(N__55291));
    InMux I__13031 (
            .O(N__55326),
            .I(N__55291));
    InMux I__13030 (
            .O(N__55325),
            .I(N__55284));
    InMux I__13029 (
            .O(N__55324),
            .I(N__55284));
    InMux I__13028 (
            .O(N__55323),
            .I(N__55284));
    InMux I__13027 (
            .O(N__55322),
            .I(N__55281));
    LocalMux I__13026 (
            .O(N__55319),
            .I(N__55278));
    LocalMux I__13025 (
            .O(N__55316),
            .I(N__55273));
    LocalMux I__13024 (
            .O(N__55311),
            .I(N__55273));
    InMux I__13023 (
            .O(N__55310),
            .I(N__55264));
    InMux I__13022 (
            .O(N__55309),
            .I(N__55264));
    InMux I__13021 (
            .O(N__55308),
            .I(N__55264));
    InMux I__13020 (
            .O(N__55307),
            .I(N__55255));
    InMux I__13019 (
            .O(N__55306),
            .I(N__55255));
    LocalMux I__13018 (
            .O(N__55301),
            .I(N__55252));
    LocalMux I__13017 (
            .O(N__55298),
            .I(N__55245));
    LocalMux I__13016 (
            .O(N__55291),
            .I(N__55245));
    LocalMux I__13015 (
            .O(N__55284),
            .I(N__55245));
    LocalMux I__13014 (
            .O(N__55281),
            .I(N__55242));
    Span4Mux_h I__13013 (
            .O(N__55278),
            .I(N__55237));
    Span4Mux_h I__13012 (
            .O(N__55273),
            .I(N__55237));
    InMux I__13011 (
            .O(N__55272),
            .I(N__55232));
    InMux I__13010 (
            .O(N__55271),
            .I(N__55232));
    LocalMux I__13009 (
            .O(N__55264),
            .I(N__55229));
    InMux I__13008 (
            .O(N__55263),
            .I(N__55224));
    InMux I__13007 (
            .O(N__55262),
            .I(N__55224));
    InMux I__13006 (
            .O(N__55261),
            .I(N__55221));
    InMux I__13005 (
            .O(N__55260),
            .I(N__55218));
    LocalMux I__13004 (
            .O(N__55255),
            .I(N__55207));
    Span4Mux_v I__13003 (
            .O(N__55252),
            .I(N__55207));
    Span4Mux_v I__13002 (
            .O(N__55245),
            .I(N__55207));
    Span4Mux_v I__13001 (
            .O(N__55242),
            .I(N__55207));
    Span4Mux_v I__13000 (
            .O(N__55237),
            .I(N__55207));
    LocalMux I__12999 (
            .O(N__55232),
            .I(N__55202));
    Span4Mux_s1_v I__12998 (
            .O(N__55229),
            .I(N__55202));
    LocalMux I__12997 (
            .O(N__55224),
            .I(duty_23));
    LocalMux I__12996 (
            .O(N__55221),
            .I(duty_23));
    LocalMux I__12995 (
            .O(N__55218),
            .I(duty_23));
    Odrv4 I__12994 (
            .O(N__55207),
            .I(duty_23));
    Odrv4 I__12993 (
            .O(N__55202),
            .I(duty_23));
    IoInMux I__12992 (
            .O(N__55191),
            .I(N__55188));
    LocalMux I__12991 (
            .O(N__55188),
            .I(N__55185));
    IoSpan4Mux I__12990 (
            .O(N__55185),
            .I(N__55182));
    Span4Mux_s1_v I__12989 (
            .O(N__55182),
            .I(N__55179));
    Odrv4 I__12988 (
            .O(N__55179),
            .I(INLB_c_0));
    InMux I__12987 (
            .O(N__55176),
            .I(N__55172));
    InMux I__12986 (
            .O(N__55175),
            .I(N__55169));
    LocalMux I__12985 (
            .O(N__55172),
            .I(sweep_counter_5));
    LocalMux I__12984 (
            .O(N__55169),
            .I(sweep_counter_5));
    InMux I__12983 (
            .O(N__55164),
            .I(n13003));
    InMux I__12982 (
            .O(N__55161),
            .I(N__55157));
    InMux I__12981 (
            .O(N__55160),
            .I(N__55154));
    LocalMux I__12980 (
            .O(N__55157),
            .I(sweep_counter_6));
    LocalMux I__12979 (
            .O(N__55154),
            .I(sweep_counter_6));
    InMux I__12978 (
            .O(N__55149),
            .I(n13004));
    InMux I__12977 (
            .O(N__55146),
            .I(N__55142));
    InMux I__12976 (
            .O(N__55145),
            .I(N__55139));
    LocalMux I__12975 (
            .O(N__55142),
            .I(sweep_counter_7));
    LocalMux I__12974 (
            .O(N__55139),
            .I(sweep_counter_7));
    InMux I__12973 (
            .O(N__55134),
            .I(n13005));
    InMux I__12972 (
            .O(N__55131),
            .I(N__55127));
    InMux I__12971 (
            .O(N__55130),
            .I(N__55124));
    LocalMux I__12970 (
            .O(N__55127),
            .I(sweep_counter_8));
    LocalMux I__12969 (
            .O(N__55124),
            .I(sweep_counter_8));
    InMux I__12968 (
            .O(N__55119),
            .I(bfn_17_27_0_));
    InMux I__12967 (
            .O(N__55116),
            .I(N__55112));
    InMux I__12966 (
            .O(N__55115),
            .I(N__55109));
    LocalMux I__12965 (
            .O(N__55112),
            .I(sweep_counter_9));
    LocalMux I__12964 (
            .O(N__55109),
            .I(sweep_counter_9));
    InMux I__12963 (
            .O(N__55104),
            .I(n13007));
    InMux I__12962 (
            .O(N__55101),
            .I(N__55097));
    InMux I__12961 (
            .O(N__55100),
            .I(N__55094));
    LocalMux I__12960 (
            .O(N__55097),
            .I(sweep_counter_10));
    LocalMux I__12959 (
            .O(N__55094),
            .I(sweep_counter_10));
    InMux I__12958 (
            .O(N__55089),
            .I(n13008));
    InMux I__12957 (
            .O(N__55086),
            .I(N__55082));
    InMux I__12956 (
            .O(N__55085),
            .I(N__55079));
    LocalMux I__12955 (
            .O(N__55082),
            .I(N__55076));
    LocalMux I__12954 (
            .O(N__55079),
            .I(sweep_counter_11));
    Odrv4 I__12953 (
            .O(N__55076),
            .I(sweep_counter_11));
    InMux I__12952 (
            .O(N__55071),
            .I(n13009));
    InMux I__12951 (
            .O(N__55068),
            .I(N__55064));
    InMux I__12950 (
            .O(N__55067),
            .I(N__55061));
    LocalMux I__12949 (
            .O(N__55064),
            .I(sweep_counter_12));
    LocalMux I__12948 (
            .O(N__55061),
            .I(sweep_counter_12));
    InMux I__12947 (
            .O(N__55056),
            .I(n13010));
    InMux I__12946 (
            .O(N__55053),
            .I(N__55049));
    InMux I__12945 (
            .O(N__55052),
            .I(N__55046));
    LocalMux I__12944 (
            .O(N__55049),
            .I(sweep_counter_13));
    LocalMux I__12943 (
            .O(N__55046),
            .I(sweep_counter_13));
    InMux I__12942 (
            .O(N__55041),
            .I(n13011));
    CascadeMux I__12941 (
            .O(N__55038),
            .I(n5183_cascade_));
    CascadeMux I__12940 (
            .O(N__55035),
            .I(N__55031));
    InMux I__12939 (
            .O(N__55034),
            .I(N__55022));
    InMux I__12938 (
            .O(N__55031),
            .I(N__55022));
    InMux I__12937 (
            .O(N__55030),
            .I(N__55019));
    InMux I__12936 (
            .O(N__55029),
            .I(N__55016));
    InMux I__12935 (
            .O(N__55028),
            .I(N__55011));
    InMux I__12934 (
            .O(N__55027),
            .I(N__55011));
    LocalMux I__12933 (
            .O(N__55022),
            .I(N__55008));
    LocalMux I__12932 (
            .O(N__55019),
            .I(dti));
    LocalMux I__12931 (
            .O(N__55016),
            .I(dti));
    LocalMux I__12930 (
            .O(N__55011),
            .I(dti));
    Odrv4 I__12929 (
            .O(N__55008),
            .I(dti));
    CascadeMux I__12928 (
            .O(N__54999),
            .I(n20_adj_706_cascade_));
    InMux I__12927 (
            .O(N__54996),
            .I(N__54993));
    LocalMux I__12926 (
            .O(N__54993),
            .I(n24_adj_704));
    InMux I__12925 (
            .O(N__54990),
            .I(N__54987));
    LocalMux I__12924 (
            .O(N__54987),
            .I(N__54983));
    InMux I__12923 (
            .O(N__54986),
            .I(N__54980));
    Odrv4 I__12922 (
            .O(N__54983),
            .I(n13187));
    LocalMux I__12921 (
            .O(N__54980),
            .I(n13187));
    InMux I__12920 (
            .O(N__54975),
            .I(N__54971));
    InMux I__12919 (
            .O(N__54974),
            .I(N__54968));
    LocalMux I__12918 (
            .O(N__54971),
            .I(sweep_counter_0));
    LocalMux I__12917 (
            .O(N__54968),
            .I(sweep_counter_0));
    InMux I__12916 (
            .O(N__54963),
            .I(bfn_17_26_0_));
    InMux I__12915 (
            .O(N__54960),
            .I(N__54956));
    InMux I__12914 (
            .O(N__54959),
            .I(N__54953));
    LocalMux I__12913 (
            .O(N__54956),
            .I(sweep_counter_1));
    LocalMux I__12912 (
            .O(N__54953),
            .I(sweep_counter_1));
    InMux I__12911 (
            .O(N__54948),
            .I(n12999));
    InMux I__12910 (
            .O(N__54945),
            .I(N__54941));
    InMux I__12909 (
            .O(N__54944),
            .I(N__54938));
    LocalMux I__12908 (
            .O(N__54941),
            .I(sweep_counter_2));
    LocalMux I__12907 (
            .O(N__54938),
            .I(sweep_counter_2));
    InMux I__12906 (
            .O(N__54933),
            .I(n13000));
    CascadeMux I__12905 (
            .O(N__54930),
            .I(N__54926));
    InMux I__12904 (
            .O(N__54929),
            .I(N__54923));
    InMux I__12903 (
            .O(N__54926),
            .I(N__54920));
    LocalMux I__12902 (
            .O(N__54923),
            .I(sweep_counter_3));
    LocalMux I__12901 (
            .O(N__54920),
            .I(sweep_counter_3));
    InMux I__12900 (
            .O(N__54915),
            .I(n13001));
    InMux I__12899 (
            .O(N__54912),
            .I(N__54908));
    InMux I__12898 (
            .O(N__54911),
            .I(N__54905));
    LocalMux I__12897 (
            .O(N__54908),
            .I(sweep_counter_4));
    LocalMux I__12896 (
            .O(N__54905),
            .I(sweep_counter_4));
    InMux I__12895 (
            .O(N__54900),
            .I(n13002));
    CascadeMux I__12894 (
            .O(N__54897),
            .I(n6_adj_582_cascade_));
    InMux I__12893 (
            .O(N__54894),
            .I(N__54888));
    InMux I__12892 (
            .O(N__54893),
            .I(N__54888));
    LocalMux I__12891 (
            .O(N__54888),
            .I(N__54885));
    Odrv4 I__12890 (
            .O(N__54885),
            .I(n14108));
    CascadeMux I__12889 (
            .O(N__54882),
            .I(N__54878));
    InMux I__12888 (
            .O(N__54881),
            .I(N__54875));
    InMux I__12887 (
            .O(N__54878),
            .I(N__54870));
    LocalMux I__12886 (
            .O(N__54875),
            .I(N__54867));
    InMux I__12885 (
            .O(N__54874),
            .I(N__54864));
    InMux I__12884 (
            .O(N__54873),
            .I(N__54861));
    LocalMux I__12883 (
            .O(N__54870),
            .I(encoder0_position_target_15));
    Odrv12 I__12882 (
            .O(N__54867),
            .I(encoder0_position_target_15));
    LocalMux I__12881 (
            .O(N__54864),
            .I(encoder0_position_target_15));
    LocalMux I__12880 (
            .O(N__54861),
            .I(encoder0_position_target_15));
    CascadeMux I__12879 (
            .O(N__54852),
            .I(N__54849));
    InMux I__12878 (
            .O(N__54849),
            .I(N__54844));
    InMux I__12877 (
            .O(N__54848),
            .I(N__54841));
    CascadeMux I__12876 (
            .O(N__54847),
            .I(N__54838));
    LocalMux I__12875 (
            .O(N__54844),
            .I(N__54835));
    LocalMux I__12874 (
            .O(N__54841),
            .I(N__54831));
    InMux I__12873 (
            .O(N__54838),
            .I(N__54828));
    Span4Mux_h I__12872 (
            .O(N__54835),
            .I(N__54825));
    InMux I__12871 (
            .O(N__54834),
            .I(N__54822));
    Span4Mux_h I__12870 (
            .O(N__54831),
            .I(N__54819));
    LocalMux I__12869 (
            .O(N__54828),
            .I(encoder0_position_target_21));
    Odrv4 I__12868 (
            .O(N__54825),
            .I(encoder0_position_target_21));
    LocalMux I__12867 (
            .O(N__54822),
            .I(encoder0_position_target_21));
    Odrv4 I__12866 (
            .O(N__54819),
            .I(encoder0_position_target_21));
    CascadeMux I__12865 (
            .O(N__54810),
            .I(N__54807));
    InMux I__12864 (
            .O(N__54807),
            .I(N__54802));
    InMux I__12863 (
            .O(N__54806),
            .I(N__54798));
    CascadeMux I__12862 (
            .O(N__54805),
            .I(N__54795));
    LocalMux I__12861 (
            .O(N__54802),
            .I(N__54792));
    CascadeMux I__12860 (
            .O(N__54801),
            .I(N__54789));
    LocalMux I__12859 (
            .O(N__54798),
            .I(N__54786));
    InMux I__12858 (
            .O(N__54795),
            .I(N__54783));
    Span4Mux_v I__12857 (
            .O(N__54792),
            .I(N__54780));
    InMux I__12856 (
            .O(N__54789),
            .I(N__54777));
    Span4Mux_h I__12855 (
            .O(N__54786),
            .I(N__54774));
    LocalMux I__12854 (
            .O(N__54783),
            .I(encoder0_position_target_19));
    Odrv4 I__12853 (
            .O(N__54780),
            .I(encoder0_position_target_19));
    LocalMux I__12852 (
            .O(N__54777),
            .I(encoder0_position_target_19));
    Odrv4 I__12851 (
            .O(N__54774),
            .I(encoder0_position_target_19));
    CascadeMux I__12850 (
            .O(N__54765),
            .I(N__54759));
    InMux I__12849 (
            .O(N__54764),
            .I(N__54756));
    InMux I__12848 (
            .O(N__54763),
            .I(N__54752));
    InMux I__12847 (
            .O(N__54762),
            .I(N__54749));
    InMux I__12846 (
            .O(N__54759),
            .I(N__54745));
    LocalMux I__12845 (
            .O(N__54756),
            .I(N__54742));
    InMux I__12844 (
            .O(N__54755),
            .I(N__54739));
    LocalMux I__12843 (
            .O(N__54752),
            .I(N__54736));
    LocalMux I__12842 (
            .O(N__54749),
            .I(N__54733));
    InMux I__12841 (
            .O(N__54748),
            .I(N__54730));
    LocalMux I__12840 (
            .O(N__54745),
            .I(N__54725));
    Span4Mux_h I__12839 (
            .O(N__54742),
            .I(N__54725));
    LocalMux I__12838 (
            .O(N__54739),
            .I(encoder0_position_target_23));
    Odrv12 I__12837 (
            .O(N__54736),
            .I(encoder0_position_target_23));
    Odrv4 I__12836 (
            .O(N__54733),
            .I(encoder0_position_target_23));
    LocalMux I__12835 (
            .O(N__54730),
            .I(encoder0_position_target_23));
    Odrv4 I__12834 (
            .O(N__54725),
            .I(encoder0_position_target_23));
    InMux I__12833 (
            .O(N__54714),
            .I(N__54711));
    LocalMux I__12832 (
            .O(N__54711),
            .I(N__54708));
    Odrv4 I__12831 (
            .O(N__54708),
            .I(n24_adj_699));
    InMux I__12830 (
            .O(N__54705),
            .I(N__54702));
    LocalMux I__12829 (
            .O(N__54702),
            .I(n16_adj_707));
    CascadeMux I__12828 (
            .O(N__54699),
            .I(N__54694));
    CascadeMux I__12827 (
            .O(N__54698),
            .I(N__54690));
    InMux I__12826 (
            .O(N__54697),
            .I(N__54685));
    InMux I__12825 (
            .O(N__54694),
            .I(N__54679));
    InMux I__12824 (
            .O(N__54693),
            .I(N__54679));
    InMux I__12823 (
            .O(N__54690),
            .I(N__54672));
    InMux I__12822 (
            .O(N__54689),
            .I(N__54672));
    InMux I__12821 (
            .O(N__54688),
            .I(N__54672));
    LocalMux I__12820 (
            .O(N__54685),
            .I(N__54667));
    InMux I__12819 (
            .O(N__54684),
            .I(N__54664));
    LocalMux I__12818 (
            .O(N__54679),
            .I(N__54659));
    LocalMux I__12817 (
            .O(N__54672),
            .I(N__54659));
    InMux I__12816 (
            .O(N__54671),
            .I(N__54656));
    InMux I__12815 (
            .O(N__54670),
            .I(N__54653));
    Odrv4 I__12814 (
            .O(N__54667),
            .I(commutation_state_prev_0));
    LocalMux I__12813 (
            .O(N__54664),
            .I(commutation_state_prev_0));
    Odrv4 I__12812 (
            .O(N__54659),
            .I(commutation_state_prev_0));
    LocalMux I__12811 (
            .O(N__54656),
            .I(commutation_state_prev_0));
    LocalMux I__12810 (
            .O(N__54653),
            .I(commutation_state_prev_0));
    CascadeMux I__12809 (
            .O(N__54642),
            .I(dti_N_333_cascade_));
    CascadeMux I__12808 (
            .O(N__54639),
            .I(N__54631));
    CascadeMux I__12807 (
            .O(N__54638),
            .I(N__54628));
    CascadeMux I__12806 (
            .O(N__54637),
            .I(N__54625));
    CascadeMux I__12805 (
            .O(N__54636),
            .I(N__54620));
    InMux I__12804 (
            .O(N__54635),
            .I(N__54617));
    InMux I__12803 (
            .O(N__54634),
            .I(N__54610));
    InMux I__12802 (
            .O(N__54631),
            .I(N__54610));
    InMux I__12801 (
            .O(N__54628),
            .I(N__54610));
    InMux I__12800 (
            .O(N__54625),
            .I(N__54605));
    InMux I__12799 (
            .O(N__54624),
            .I(N__54605));
    InMux I__12798 (
            .O(N__54623),
            .I(N__54602));
    InMux I__12797 (
            .O(N__54620),
            .I(N__54599));
    LocalMux I__12796 (
            .O(N__54617),
            .I(N__54596));
    LocalMux I__12795 (
            .O(N__54610),
            .I(N__54591));
    LocalMux I__12794 (
            .O(N__54605),
            .I(N__54591));
    LocalMux I__12793 (
            .O(N__54602),
            .I(n4_adj_716));
    LocalMux I__12792 (
            .O(N__54599),
            .I(n4_adj_716));
    Odrv4 I__12791 (
            .O(N__54596),
            .I(n4_adj_716));
    Odrv4 I__12790 (
            .O(N__54591),
            .I(n4_adj_716));
    CEMux I__12789 (
            .O(N__54582),
            .I(N__54579));
    LocalMux I__12788 (
            .O(N__54579),
            .I(n5169));
    CascadeMux I__12787 (
            .O(N__54576),
            .I(N__54573));
    InMux I__12786 (
            .O(N__54573),
            .I(N__54570));
    LocalMux I__12785 (
            .O(N__54570),
            .I(n1377));
    InMux I__12784 (
            .O(N__54567),
            .I(N__54561));
    InMux I__12783 (
            .O(N__54566),
            .I(N__54558));
    InMux I__12782 (
            .O(N__54565),
            .I(N__54553));
    InMux I__12781 (
            .O(N__54564),
            .I(N__54553));
    LocalMux I__12780 (
            .O(N__54561),
            .I(n5119));
    LocalMux I__12779 (
            .O(N__54558),
            .I(n5119));
    LocalMux I__12778 (
            .O(N__54553),
            .I(n5119));
    CascadeMux I__12777 (
            .O(N__54546),
            .I(N__54540));
    CascadeMux I__12776 (
            .O(N__54545),
            .I(N__54536));
    CascadeMux I__12775 (
            .O(N__54544),
            .I(N__54531));
    CascadeMux I__12774 (
            .O(N__54543),
            .I(N__54523));
    InMux I__12773 (
            .O(N__54540),
            .I(N__54491));
    InMux I__12772 (
            .O(N__54539),
            .I(N__54491));
    InMux I__12771 (
            .O(N__54536),
            .I(N__54491));
    InMux I__12770 (
            .O(N__54535),
            .I(N__54491));
    InMux I__12769 (
            .O(N__54534),
            .I(N__54491));
    InMux I__12768 (
            .O(N__54531),
            .I(N__54484));
    InMux I__12767 (
            .O(N__54530),
            .I(N__54484));
    InMux I__12766 (
            .O(N__54529),
            .I(N__54484));
    InMux I__12765 (
            .O(N__54528),
            .I(N__54477));
    InMux I__12764 (
            .O(N__54527),
            .I(N__54477));
    InMux I__12763 (
            .O(N__54526),
            .I(N__54477));
    InMux I__12762 (
            .O(N__54523),
            .I(N__54466));
    InMux I__12761 (
            .O(N__54522),
            .I(N__54466));
    InMux I__12760 (
            .O(N__54521),
            .I(N__54466));
    InMux I__12759 (
            .O(N__54520),
            .I(N__54466));
    InMux I__12758 (
            .O(N__54519),
            .I(N__54466));
    CascadeMux I__12757 (
            .O(N__54518),
            .I(N__54462));
    CascadeMux I__12756 (
            .O(N__54517),
            .I(N__54452));
    CascadeMux I__12755 (
            .O(N__54516),
            .I(N__54449));
    CascadeMux I__12754 (
            .O(N__54515),
            .I(N__54446));
    CascadeMux I__12753 (
            .O(N__54514),
            .I(N__54443));
    CascadeMux I__12752 (
            .O(N__54513),
            .I(N__54440));
    CascadeMux I__12751 (
            .O(N__54512),
            .I(N__54437));
    CascadeMux I__12750 (
            .O(N__54511),
            .I(N__54434));
    CascadeMux I__12749 (
            .O(N__54510),
            .I(N__54431));
    CascadeMux I__12748 (
            .O(N__54509),
            .I(N__54428));
    CascadeMux I__12747 (
            .O(N__54508),
            .I(N__54425));
    CascadeMux I__12746 (
            .O(N__54507),
            .I(N__54419));
    CascadeMux I__12745 (
            .O(N__54506),
            .I(N__54410));
    CascadeMux I__12744 (
            .O(N__54505),
            .I(N__54407));
    CascadeMux I__12743 (
            .O(N__54504),
            .I(N__54396));
    CascadeMux I__12742 (
            .O(N__54503),
            .I(N__54392));
    CascadeMux I__12741 (
            .O(N__54502),
            .I(N__54386));
    LocalMux I__12740 (
            .O(N__54491),
            .I(N__54381));
    LocalMux I__12739 (
            .O(N__54484),
            .I(N__54381));
    LocalMux I__12738 (
            .O(N__54477),
            .I(N__54376));
    LocalMux I__12737 (
            .O(N__54466),
            .I(N__54376));
    InMux I__12736 (
            .O(N__54465),
            .I(N__54371));
    InMux I__12735 (
            .O(N__54462),
            .I(N__54371));
    InMux I__12734 (
            .O(N__54461),
            .I(N__54366));
    InMux I__12733 (
            .O(N__54460),
            .I(N__54366));
    CascadeMux I__12732 (
            .O(N__54459),
            .I(N__54362));
    CascadeMux I__12731 (
            .O(N__54458),
            .I(N__54355));
    CascadeMux I__12730 (
            .O(N__54457),
            .I(N__54347));
    CascadeMux I__12729 (
            .O(N__54456),
            .I(N__54342));
    InMux I__12728 (
            .O(N__54455),
            .I(N__54337));
    InMux I__12727 (
            .O(N__54452),
            .I(N__54337));
    InMux I__12726 (
            .O(N__54449),
            .I(N__54334));
    InMux I__12725 (
            .O(N__54446),
            .I(N__54325));
    InMux I__12724 (
            .O(N__54443),
            .I(N__54325));
    InMux I__12723 (
            .O(N__54440),
            .I(N__54325));
    InMux I__12722 (
            .O(N__54437),
            .I(N__54325));
    InMux I__12721 (
            .O(N__54434),
            .I(N__54316));
    InMux I__12720 (
            .O(N__54431),
            .I(N__54316));
    InMux I__12719 (
            .O(N__54428),
            .I(N__54316));
    InMux I__12718 (
            .O(N__54425),
            .I(N__54316));
    InMux I__12717 (
            .O(N__54424),
            .I(N__54309));
    InMux I__12716 (
            .O(N__54423),
            .I(N__54309));
    InMux I__12715 (
            .O(N__54422),
            .I(N__54309));
    InMux I__12714 (
            .O(N__54419),
            .I(N__54298));
    InMux I__12713 (
            .O(N__54418),
            .I(N__54298));
    InMux I__12712 (
            .O(N__54417),
            .I(N__54298));
    InMux I__12711 (
            .O(N__54416),
            .I(N__54298));
    InMux I__12710 (
            .O(N__54415),
            .I(N__54298));
    InMux I__12709 (
            .O(N__54414),
            .I(N__54259));
    InMux I__12708 (
            .O(N__54413),
            .I(N__54252));
    InMux I__12707 (
            .O(N__54410),
            .I(N__54252));
    InMux I__12706 (
            .O(N__54407),
            .I(N__54252));
    InMux I__12705 (
            .O(N__54406),
            .I(N__54249));
    InMux I__12704 (
            .O(N__54405),
            .I(N__54242));
    InMux I__12703 (
            .O(N__54404),
            .I(N__54242));
    InMux I__12702 (
            .O(N__54403),
            .I(N__54242));
    InMux I__12701 (
            .O(N__54402),
            .I(N__54239));
    InMux I__12700 (
            .O(N__54401),
            .I(N__54232));
    InMux I__12699 (
            .O(N__54400),
            .I(N__54232));
    InMux I__12698 (
            .O(N__54399),
            .I(N__54232));
    InMux I__12697 (
            .O(N__54396),
            .I(N__54219));
    InMux I__12696 (
            .O(N__54395),
            .I(N__54219));
    InMux I__12695 (
            .O(N__54392),
            .I(N__54219));
    InMux I__12694 (
            .O(N__54391),
            .I(N__54219));
    InMux I__12693 (
            .O(N__54390),
            .I(N__54219));
    InMux I__12692 (
            .O(N__54389),
            .I(N__54219));
    InMux I__12691 (
            .O(N__54386),
            .I(N__54216));
    Span4Mux_s3_h I__12690 (
            .O(N__54381),
            .I(N__54207));
    Span4Mux_v I__12689 (
            .O(N__54376),
            .I(N__54207));
    LocalMux I__12688 (
            .O(N__54371),
            .I(N__54207));
    LocalMux I__12687 (
            .O(N__54366),
            .I(N__54207));
    InMux I__12686 (
            .O(N__54365),
            .I(N__54202));
    InMux I__12685 (
            .O(N__54362),
            .I(N__54202));
    CascadeMux I__12684 (
            .O(N__54361),
            .I(N__54198));
    CascadeMux I__12683 (
            .O(N__54360),
            .I(N__54194));
    CascadeMux I__12682 (
            .O(N__54359),
            .I(N__54191));
    InMux I__12681 (
            .O(N__54358),
            .I(N__54169));
    InMux I__12680 (
            .O(N__54355),
            .I(N__54169));
    InMux I__12679 (
            .O(N__54354),
            .I(N__54169));
    InMux I__12678 (
            .O(N__54353),
            .I(N__54164));
    InMux I__12677 (
            .O(N__54352),
            .I(N__54164));
    InMux I__12676 (
            .O(N__54351),
            .I(N__54151));
    InMux I__12675 (
            .O(N__54350),
            .I(N__54151));
    InMux I__12674 (
            .O(N__54347),
            .I(N__54151));
    InMux I__12673 (
            .O(N__54346),
            .I(N__54151));
    InMux I__12672 (
            .O(N__54345),
            .I(N__54151));
    InMux I__12671 (
            .O(N__54342),
            .I(N__54151));
    LocalMux I__12670 (
            .O(N__54337),
            .I(N__54138));
    LocalMux I__12669 (
            .O(N__54334),
            .I(N__54138));
    LocalMux I__12668 (
            .O(N__54325),
            .I(N__54138));
    LocalMux I__12667 (
            .O(N__54316),
            .I(N__54138));
    LocalMux I__12666 (
            .O(N__54309),
            .I(N__54138));
    LocalMux I__12665 (
            .O(N__54298),
            .I(N__54138));
    InMux I__12664 (
            .O(N__54297),
            .I(N__54135));
    CascadeMux I__12663 (
            .O(N__54296),
            .I(N__54131));
    CascadeMux I__12662 (
            .O(N__54295),
            .I(N__54128));
    CascadeMux I__12661 (
            .O(N__54294),
            .I(N__54125));
    CascadeMux I__12660 (
            .O(N__54293),
            .I(N__54122));
    CascadeMux I__12659 (
            .O(N__54292),
            .I(N__54118));
    CascadeMux I__12658 (
            .O(N__54291),
            .I(N__54115));
    CascadeMux I__12657 (
            .O(N__54290),
            .I(N__54112));
    CascadeMux I__12656 (
            .O(N__54289),
            .I(N__54109));
    CascadeMux I__12655 (
            .O(N__54288),
            .I(N__54106));
    CascadeMux I__12654 (
            .O(N__54287),
            .I(N__54103));
    CascadeMux I__12653 (
            .O(N__54286),
            .I(N__54099));
    CascadeMux I__12652 (
            .O(N__54285),
            .I(N__54088));
    CascadeMux I__12651 (
            .O(N__54284),
            .I(N__54085));
    CascadeMux I__12650 (
            .O(N__54283),
            .I(N__54082));
    CascadeMux I__12649 (
            .O(N__54282),
            .I(N__54075));
    CascadeMux I__12648 (
            .O(N__54281),
            .I(N__54072));
    CascadeMux I__12647 (
            .O(N__54280),
            .I(N__54069));
    CascadeMux I__12646 (
            .O(N__54279),
            .I(N__54066));
    CascadeMux I__12645 (
            .O(N__54278),
            .I(N__54063));
    CascadeMux I__12644 (
            .O(N__54277),
            .I(N__54059));
    CascadeMux I__12643 (
            .O(N__54276),
            .I(N__54056));
    CascadeMux I__12642 (
            .O(N__54275),
            .I(N__54053));
    CascadeMux I__12641 (
            .O(N__54274),
            .I(N__54049));
    CascadeMux I__12640 (
            .O(N__54273),
            .I(N__54046));
    CascadeMux I__12639 (
            .O(N__54272),
            .I(N__54043));
    CascadeMux I__12638 (
            .O(N__54271),
            .I(N__54040));
    CascadeMux I__12637 (
            .O(N__54270),
            .I(N__54037));
    CascadeMux I__12636 (
            .O(N__54269),
            .I(N__54034));
    CascadeMux I__12635 (
            .O(N__54268),
            .I(N__54031));
    CascadeMux I__12634 (
            .O(N__54267),
            .I(N__54028));
    CascadeMux I__12633 (
            .O(N__54266),
            .I(N__54025));
    CascadeMux I__12632 (
            .O(N__54265),
            .I(N__54022));
    CascadeMux I__12631 (
            .O(N__54264),
            .I(N__54019));
    CascadeMux I__12630 (
            .O(N__54263),
            .I(N__54015));
    CascadeMux I__12629 (
            .O(N__54262),
            .I(N__54012));
    LocalMux I__12628 (
            .O(N__54259),
            .I(N__53968));
    LocalMux I__12627 (
            .O(N__54252),
            .I(N__53968));
    LocalMux I__12626 (
            .O(N__54249),
            .I(N__53968));
    LocalMux I__12625 (
            .O(N__54242),
            .I(N__53968));
    LocalMux I__12624 (
            .O(N__54239),
            .I(N__53968));
    LocalMux I__12623 (
            .O(N__54232),
            .I(N__53968));
    LocalMux I__12622 (
            .O(N__54219),
            .I(N__53963));
    LocalMux I__12621 (
            .O(N__54216),
            .I(N__53963));
    Span4Mux_h I__12620 (
            .O(N__54207),
            .I(N__53958));
    LocalMux I__12619 (
            .O(N__54202),
            .I(N__53958));
    InMux I__12618 (
            .O(N__54201),
            .I(N__53955));
    InMux I__12617 (
            .O(N__54198),
            .I(N__53948));
    InMux I__12616 (
            .O(N__54197),
            .I(N__53948));
    InMux I__12615 (
            .O(N__54194),
            .I(N__53948));
    InMux I__12614 (
            .O(N__54191),
            .I(N__53943));
    InMux I__12613 (
            .O(N__54190),
            .I(N__53943));
    InMux I__12612 (
            .O(N__54189),
            .I(N__53938));
    InMux I__12611 (
            .O(N__54188),
            .I(N__53938));
    CascadeMux I__12610 (
            .O(N__54187),
            .I(N__53930));
    CascadeMux I__12609 (
            .O(N__54186),
            .I(N__53927));
    CascadeMux I__12608 (
            .O(N__54185),
            .I(N__53922));
    CascadeMux I__12607 (
            .O(N__54184),
            .I(N__53918));
    CascadeMux I__12606 (
            .O(N__54183),
            .I(N__53912));
    CascadeMux I__12605 (
            .O(N__54182),
            .I(N__53909));
    CascadeMux I__12604 (
            .O(N__54181),
            .I(N__53906));
    CascadeMux I__12603 (
            .O(N__54180),
            .I(N__53899));
    CascadeMux I__12602 (
            .O(N__54179),
            .I(N__53893));
    CascadeMux I__12601 (
            .O(N__54178),
            .I(N__53885));
    CascadeMux I__12600 (
            .O(N__54177),
            .I(N__53882));
    CascadeMux I__12599 (
            .O(N__54176),
            .I(N__53879));
    LocalMux I__12598 (
            .O(N__54169),
            .I(N__53872));
    LocalMux I__12597 (
            .O(N__54164),
            .I(N__53872));
    LocalMux I__12596 (
            .O(N__54151),
            .I(N__53872));
    Span4Mux_v I__12595 (
            .O(N__54138),
            .I(N__53867));
    LocalMux I__12594 (
            .O(N__54135),
            .I(N__53867));
    InMux I__12593 (
            .O(N__54134),
            .I(N__53860));
    InMux I__12592 (
            .O(N__54131),
            .I(N__53860));
    InMux I__12591 (
            .O(N__54128),
            .I(N__53860));
    InMux I__12590 (
            .O(N__54125),
            .I(N__53853));
    InMux I__12589 (
            .O(N__54122),
            .I(N__53853));
    InMux I__12588 (
            .O(N__54121),
            .I(N__53853));
    InMux I__12587 (
            .O(N__54118),
            .I(N__53846));
    InMux I__12586 (
            .O(N__54115),
            .I(N__53846));
    InMux I__12585 (
            .O(N__54112),
            .I(N__53846));
    InMux I__12584 (
            .O(N__54109),
            .I(N__53835));
    InMux I__12583 (
            .O(N__54106),
            .I(N__53835));
    InMux I__12582 (
            .O(N__54103),
            .I(N__53835));
    InMux I__12581 (
            .O(N__54102),
            .I(N__53835));
    InMux I__12580 (
            .O(N__54099),
            .I(N__53835));
    InMux I__12579 (
            .O(N__54098),
            .I(N__53828));
    InMux I__12578 (
            .O(N__54097),
            .I(N__53828));
    InMux I__12577 (
            .O(N__54096),
            .I(N__53828));
    CascadeMux I__12576 (
            .O(N__54095),
            .I(N__53825));
    CascadeMux I__12575 (
            .O(N__54094),
            .I(N__53822));
    CascadeMux I__12574 (
            .O(N__54093),
            .I(N__53819));
    CascadeMux I__12573 (
            .O(N__54092),
            .I(N__53815));
    InMux I__12572 (
            .O(N__54091),
            .I(N__53802));
    InMux I__12571 (
            .O(N__54088),
            .I(N__53802));
    InMux I__12570 (
            .O(N__54085),
            .I(N__53797));
    InMux I__12569 (
            .O(N__54082),
            .I(N__53797));
    CascadeMux I__12568 (
            .O(N__54081),
            .I(N__53794));
    CascadeMux I__12567 (
            .O(N__54080),
            .I(N__53789));
    CascadeMux I__12566 (
            .O(N__54079),
            .I(N__53786));
    InMux I__12565 (
            .O(N__54078),
            .I(N__53776));
    InMux I__12564 (
            .O(N__54075),
            .I(N__53776));
    InMux I__12563 (
            .O(N__54072),
            .I(N__53776));
    InMux I__12562 (
            .O(N__54069),
            .I(N__53769));
    InMux I__12561 (
            .O(N__54066),
            .I(N__53769));
    InMux I__12560 (
            .O(N__54063),
            .I(N__53769));
    InMux I__12559 (
            .O(N__54062),
            .I(N__53766));
    InMux I__12558 (
            .O(N__54059),
            .I(N__53758));
    InMux I__12557 (
            .O(N__54056),
            .I(N__53758));
    InMux I__12556 (
            .O(N__54053),
            .I(N__53747));
    InMux I__12555 (
            .O(N__54052),
            .I(N__53747));
    InMux I__12554 (
            .O(N__54049),
            .I(N__53747));
    InMux I__12553 (
            .O(N__54046),
            .I(N__53747));
    InMux I__12552 (
            .O(N__54043),
            .I(N__53747));
    InMux I__12551 (
            .O(N__54040),
            .I(N__53738));
    InMux I__12550 (
            .O(N__54037),
            .I(N__53738));
    InMux I__12549 (
            .O(N__54034),
            .I(N__53738));
    InMux I__12548 (
            .O(N__54031),
            .I(N__53738));
    InMux I__12547 (
            .O(N__54028),
            .I(N__53729));
    InMux I__12546 (
            .O(N__54025),
            .I(N__53729));
    InMux I__12545 (
            .O(N__54022),
            .I(N__53729));
    InMux I__12544 (
            .O(N__54019),
            .I(N__53729));
    InMux I__12543 (
            .O(N__54018),
            .I(N__53718));
    InMux I__12542 (
            .O(N__54015),
            .I(N__53718));
    InMux I__12541 (
            .O(N__54012),
            .I(N__53718));
    InMux I__12540 (
            .O(N__54011),
            .I(N__53718));
    InMux I__12539 (
            .O(N__54010),
            .I(N__53718));
    CascadeMux I__12538 (
            .O(N__54009),
            .I(N__53710));
    CascadeMux I__12537 (
            .O(N__54008),
            .I(N__53704));
    CascadeMux I__12536 (
            .O(N__54007),
            .I(N__53701));
    CascadeMux I__12535 (
            .O(N__54006),
            .I(N__53698));
    CascadeMux I__12534 (
            .O(N__54005),
            .I(N__53695));
    CascadeMux I__12533 (
            .O(N__54004),
            .I(N__53691));
    CascadeMux I__12532 (
            .O(N__54003),
            .I(N__53688));
    CascadeMux I__12531 (
            .O(N__54002),
            .I(N__53685));
    CascadeMux I__12530 (
            .O(N__54001),
            .I(N__53682));
    CascadeMux I__12529 (
            .O(N__54000),
            .I(N__53679));
    CascadeMux I__12528 (
            .O(N__53999),
            .I(N__53676));
    CascadeMux I__12527 (
            .O(N__53998),
            .I(N__53673));
    CascadeMux I__12526 (
            .O(N__53997),
            .I(N__53670));
    CascadeMux I__12525 (
            .O(N__53996),
            .I(N__53667));
    CascadeMux I__12524 (
            .O(N__53995),
            .I(N__53664));
    CascadeMux I__12523 (
            .O(N__53994),
            .I(N__53661));
    CascadeMux I__12522 (
            .O(N__53993),
            .I(N__53658));
    CascadeMux I__12521 (
            .O(N__53992),
            .I(N__53655));
    CascadeMux I__12520 (
            .O(N__53991),
            .I(N__53652));
    CascadeMux I__12519 (
            .O(N__53990),
            .I(N__53649));
    CascadeMux I__12518 (
            .O(N__53989),
            .I(N__53646));
    CascadeMux I__12517 (
            .O(N__53988),
            .I(N__53643));
    CascadeMux I__12516 (
            .O(N__53987),
            .I(N__53640));
    CascadeMux I__12515 (
            .O(N__53986),
            .I(N__53633));
    CascadeMux I__12514 (
            .O(N__53985),
            .I(N__53630));
    CascadeMux I__12513 (
            .O(N__53984),
            .I(N__53627));
    CascadeMux I__12512 (
            .O(N__53983),
            .I(N__53624));
    CascadeMux I__12511 (
            .O(N__53982),
            .I(N__53621));
    CascadeMux I__12510 (
            .O(N__53981),
            .I(N__53617));
    Span4Mux_h I__12509 (
            .O(N__53968),
            .I(N__53596));
    Span4Mux_v I__12508 (
            .O(N__53963),
            .I(N__53596));
    Span4Mux_v I__12507 (
            .O(N__53958),
            .I(N__53596));
    LocalMux I__12506 (
            .O(N__53955),
            .I(N__53596));
    LocalMux I__12505 (
            .O(N__53948),
            .I(N__53596));
    LocalMux I__12504 (
            .O(N__53943),
            .I(N__53593));
    LocalMux I__12503 (
            .O(N__53938),
            .I(N__53590));
    InMux I__12502 (
            .O(N__53937),
            .I(N__53587));
    CascadeMux I__12501 (
            .O(N__53936),
            .I(N__53580));
    CascadeMux I__12500 (
            .O(N__53935),
            .I(N__53573));
    CascadeMux I__12499 (
            .O(N__53934),
            .I(N__53568));
    CascadeMux I__12498 (
            .O(N__53933),
            .I(N__53565));
    InMux I__12497 (
            .O(N__53930),
            .I(N__53547));
    InMux I__12496 (
            .O(N__53927),
            .I(N__53547));
    InMux I__12495 (
            .O(N__53926),
            .I(N__53547));
    InMux I__12494 (
            .O(N__53925),
            .I(N__53547));
    InMux I__12493 (
            .O(N__53922),
            .I(N__53547));
    CascadeMux I__12492 (
            .O(N__53921),
            .I(N__53543));
    InMux I__12491 (
            .O(N__53918),
            .I(N__53536));
    InMux I__12490 (
            .O(N__53917),
            .I(N__53536));
    InMux I__12489 (
            .O(N__53916),
            .I(N__53536));
    InMux I__12488 (
            .O(N__53915),
            .I(N__53531));
    InMux I__12487 (
            .O(N__53912),
            .I(N__53531));
    InMux I__12486 (
            .O(N__53909),
            .I(N__53526));
    InMux I__12485 (
            .O(N__53906),
            .I(N__53526));
    InMux I__12484 (
            .O(N__53905),
            .I(N__53523));
    InMux I__12483 (
            .O(N__53904),
            .I(N__53516));
    InMux I__12482 (
            .O(N__53903),
            .I(N__53516));
    InMux I__12481 (
            .O(N__53902),
            .I(N__53516));
    InMux I__12480 (
            .O(N__53899),
            .I(N__53507));
    InMux I__12479 (
            .O(N__53898),
            .I(N__53507));
    InMux I__12478 (
            .O(N__53897),
            .I(N__53507));
    InMux I__12477 (
            .O(N__53896),
            .I(N__53507));
    InMux I__12476 (
            .O(N__53893),
            .I(N__53498));
    InMux I__12475 (
            .O(N__53892),
            .I(N__53498));
    InMux I__12474 (
            .O(N__53891),
            .I(N__53498));
    InMux I__12473 (
            .O(N__53890),
            .I(N__53498));
    CascadeMux I__12472 (
            .O(N__53889),
            .I(N__53495));
    CascadeMux I__12471 (
            .O(N__53888),
            .I(N__53492));
    InMux I__12470 (
            .O(N__53885),
            .I(N__53484));
    InMux I__12469 (
            .O(N__53882),
            .I(N__53484));
    InMux I__12468 (
            .O(N__53879),
            .I(N__53484));
    Span4Mux_h I__12467 (
            .O(N__53872),
            .I(N__53471));
    Span4Mux_h I__12466 (
            .O(N__53867),
            .I(N__53471));
    LocalMux I__12465 (
            .O(N__53860),
            .I(N__53471));
    LocalMux I__12464 (
            .O(N__53853),
            .I(N__53471));
    LocalMux I__12463 (
            .O(N__53846),
            .I(N__53471));
    LocalMux I__12462 (
            .O(N__53835),
            .I(N__53471));
    LocalMux I__12461 (
            .O(N__53828),
            .I(N__53468));
    InMux I__12460 (
            .O(N__53825),
            .I(N__53457));
    InMux I__12459 (
            .O(N__53822),
            .I(N__53457));
    InMux I__12458 (
            .O(N__53819),
            .I(N__53457));
    InMux I__12457 (
            .O(N__53818),
            .I(N__53457));
    InMux I__12456 (
            .O(N__53815),
            .I(N__53457));
    InMux I__12455 (
            .O(N__53814),
            .I(N__53454));
    CascadeMux I__12454 (
            .O(N__53813),
            .I(N__53446));
    CascadeMux I__12453 (
            .O(N__53812),
            .I(N__53442));
    CascadeMux I__12452 (
            .O(N__53811),
            .I(N__53429));
    CascadeMux I__12451 (
            .O(N__53810),
            .I(N__53426));
    CascadeMux I__12450 (
            .O(N__53809),
            .I(N__53422));
    CascadeMux I__12449 (
            .O(N__53808),
            .I(N__53419));
    CascadeMux I__12448 (
            .O(N__53807),
            .I(N__53414));
    LocalMux I__12447 (
            .O(N__53802),
            .I(N__53406));
    LocalMux I__12446 (
            .O(N__53797),
            .I(N__53406));
    InMux I__12445 (
            .O(N__53794),
            .I(N__53399));
    InMux I__12444 (
            .O(N__53793),
            .I(N__53399));
    InMux I__12443 (
            .O(N__53792),
            .I(N__53399));
    InMux I__12442 (
            .O(N__53789),
            .I(N__53388));
    InMux I__12441 (
            .O(N__53786),
            .I(N__53388));
    InMux I__12440 (
            .O(N__53785),
            .I(N__53388));
    InMux I__12439 (
            .O(N__53784),
            .I(N__53388));
    InMux I__12438 (
            .O(N__53783),
            .I(N__53388));
    LocalMux I__12437 (
            .O(N__53776),
            .I(N__53380));
    LocalMux I__12436 (
            .O(N__53769),
            .I(N__53380));
    LocalMux I__12435 (
            .O(N__53766),
            .I(N__53377));
    InMux I__12434 (
            .O(N__53765),
            .I(N__53370));
    InMux I__12433 (
            .O(N__53764),
            .I(N__53370));
    InMux I__12432 (
            .O(N__53763),
            .I(N__53370));
    LocalMux I__12431 (
            .O(N__53758),
            .I(N__53359));
    LocalMux I__12430 (
            .O(N__53747),
            .I(N__53359));
    LocalMux I__12429 (
            .O(N__53738),
            .I(N__53359));
    LocalMux I__12428 (
            .O(N__53729),
            .I(N__53359));
    LocalMux I__12427 (
            .O(N__53718),
            .I(N__53359));
    InMux I__12426 (
            .O(N__53717),
            .I(N__53356));
    InMux I__12425 (
            .O(N__53716),
            .I(N__53349));
    InMux I__12424 (
            .O(N__53715),
            .I(N__53349));
    InMux I__12423 (
            .O(N__53714),
            .I(N__53349));
    InMux I__12422 (
            .O(N__53713),
            .I(N__53340));
    InMux I__12421 (
            .O(N__53710),
            .I(N__53340));
    InMux I__12420 (
            .O(N__53709),
            .I(N__53340));
    InMux I__12419 (
            .O(N__53708),
            .I(N__53340));
    InMux I__12418 (
            .O(N__53707),
            .I(N__53330));
    InMux I__12417 (
            .O(N__53704),
            .I(N__53330));
    InMux I__12416 (
            .O(N__53701),
            .I(N__53330));
    InMux I__12415 (
            .O(N__53698),
            .I(N__53330));
    InMux I__12414 (
            .O(N__53695),
            .I(N__53319));
    InMux I__12413 (
            .O(N__53694),
            .I(N__53319));
    InMux I__12412 (
            .O(N__53691),
            .I(N__53319));
    InMux I__12411 (
            .O(N__53688),
            .I(N__53319));
    InMux I__12410 (
            .O(N__53685),
            .I(N__53319));
    InMux I__12409 (
            .O(N__53682),
            .I(N__53310));
    InMux I__12408 (
            .O(N__53679),
            .I(N__53310));
    InMux I__12407 (
            .O(N__53676),
            .I(N__53310));
    InMux I__12406 (
            .O(N__53673),
            .I(N__53310));
    InMux I__12405 (
            .O(N__53670),
            .I(N__53301));
    InMux I__12404 (
            .O(N__53667),
            .I(N__53301));
    InMux I__12403 (
            .O(N__53664),
            .I(N__53301));
    InMux I__12402 (
            .O(N__53661),
            .I(N__53301));
    InMux I__12401 (
            .O(N__53658),
            .I(N__53292));
    InMux I__12400 (
            .O(N__53655),
            .I(N__53292));
    InMux I__12399 (
            .O(N__53652),
            .I(N__53292));
    InMux I__12398 (
            .O(N__53649),
            .I(N__53292));
    InMux I__12397 (
            .O(N__53646),
            .I(N__53285));
    InMux I__12396 (
            .O(N__53643),
            .I(N__53285));
    InMux I__12395 (
            .O(N__53640),
            .I(N__53285));
    CascadeMux I__12394 (
            .O(N__53639),
            .I(N__53282));
    CascadeMux I__12393 (
            .O(N__53638),
            .I(N__53279));
    CascadeMux I__12392 (
            .O(N__53637),
            .I(N__53276));
    CascadeMux I__12391 (
            .O(N__53636),
            .I(N__53273));
    InMux I__12390 (
            .O(N__53633),
            .I(N__53268));
    InMux I__12389 (
            .O(N__53630),
            .I(N__53268));
    InMux I__12388 (
            .O(N__53627),
            .I(N__53255));
    InMux I__12387 (
            .O(N__53624),
            .I(N__53255));
    InMux I__12386 (
            .O(N__53621),
            .I(N__53255));
    InMux I__12385 (
            .O(N__53620),
            .I(N__53255));
    InMux I__12384 (
            .O(N__53617),
            .I(N__53255));
    InMux I__12383 (
            .O(N__53616),
            .I(N__53255));
    InMux I__12382 (
            .O(N__53615),
            .I(N__53248));
    InMux I__12381 (
            .O(N__53614),
            .I(N__53241));
    InMux I__12380 (
            .O(N__53613),
            .I(N__53241));
    InMux I__12379 (
            .O(N__53612),
            .I(N__53241));
    InMux I__12378 (
            .O(N__53611),
            .I(N__53234));
    InMux I__12377 (
            .O(N__53610),
            .I(N__53234));
    InMux I__12376 (
            .O(N__53609),
            .I(N__53234));
    InMux I__12375 (
            .O(N__53608),
            .I(N__53229));
    InMux I__12374 (
            .O(N__53607),
            .I(N__53229));
    Span4Mux_h I__12373 (
            .O(N__53596),
            .I(N__53220));
    Span4Mux_v I__12372 (
            .O(N__53593),
            .I(N__53220));
    Span4Mux_v I__12371 (
            .O(N__53590),
            .I(N__53220));
    LocalMux I__12370 (
            .O(N__53587),
            .I(N__53220));
    InMux I__12369 (
            .O(N__53586),
            .I(N__53213));
    InMux I__12368 (
            .O(N__53585),
            .I(N__53213));
    InMux I__12367 (
            .O(N__53584),
            .I(N__53213));
    InMux I__12366 (
            .O(N__53583),
            .I(N__53202));
    InMux I__12365 (
            .O(N__53580),
            .I(N__53202));
    InMux I__12364 (
            .O(N__53579),
            .I(N__53202));
    InMux I__12363 (
            .O(N__53578),
            .I(N__53202));
    InMux I__12362 (
            .O(N__53577),
            .I(N__53202));
    CascadeMux I__12361 (
            .O(N__53576),
            .I(N__53199));
    InMux I__12360 (
            .O(N__53573),
            .I(N__53180));
    InMux I__12359 (
            .O(N__53572),
            .I(N__53180));
    InMux I__12358 (
            .O(N__53571),
            .I(N__53180));
    InMux I__12357 (
            .O(N__53568),
            .I(N__53169));
    InMux I__12356 (
            .O(N__53565),
            .I(N__53169));
    InMux I__12355 (
            .O(N__53564),
            .I(N__53169));
    InMux I__12354 (
            .O(N__53563),
            .I(N__53169));
    InMux I__12353 (
            .O(N__53562),
            .I(N__53169));
    InMux I__12352 (
            .O(N__53561),
            .I(N__53164));
    InMux I__12351 (
            .O(N__53560),
            .I(N__53164));
    CascadeMux I__12350 (
            .O(N__53559),
            .I(N__53161));
    CascadeMux I__12349 (
            .O(N__53558),
            .I(N__53155));
    LocalMux I__12348 (
            .O(N__53547),
            .I(N__53149));
    InMux I__12347 (
            .O(N__53546),
            .I(N__53144));
    InMux I__12346 (
            .O(N__53543),
            .I(N__53144));
    LocalMux I__12345 (
            .O(N__53536),
            .I(N__53141));
    LocalMux I__12344 (
            .O(N__53531),
            .I(N__53128));
    LocalMux I__12343 (
            .O(N__53526),
            .I(N__53128));
    LocalMux I__12342 (
            .O(N__53523),
            .I(N__53128));
    LocalMux I__12341 (
            .O(N__53516),
            .I(N__53128));
    LocalMux I__12340 (
            .O(N__53507),
            .I(N__53128));
    LocalMux I__12339 (
            .O(N__53498),
            .I(N__53128));
    InMux I__12338 (
            .O(N__53495),
            .I(N__53121));
    InMux I__12337 (
            .O(N__53492),
            .I(N__53121));
    InMux I__12336 (
            .O(N__53491),
            .I(N__53121));
    LocalMux I__12335 (
            .O(N__53484),
            .I(N__53116));
    Span4Mux_v I__12334 (
            .O(N__53471),
            .I(N__53116));
    Span4Mux_v I__12333 (
            .O(N__53468),
            .I(N__53109));
    LocalMux I__12332 (
            .O(N__53457),
            .I(N__53109));
    LocalMux I__12331 (
            .O(N__53454),
            .I(N__53109));
    InMux I__12330 (
            .O(N__53453),
            .I(N__53104));
    InMux I__12329 (
            .O(N__53452),
            .I(N__53104));
    CascadeMux I__12328 (
            .O(N__53451),
            .I(N__53096));
    CascadeMux I__12327 (
            .O(N__53450),
            .I(N__53092));
    CascadeMux I__12326 (
            .O(N__53449),
            .I(N__53087));
    InMux I__12325 (
            .O(N__53446),
            .I(N__53082));
    InMux I__12324 (
            .O(N__53445),
            .I(N__53075));
    InMux I__12323 (
            .O(N__53442),
            .I(N__53075));
    InMux I__12322 (
            .O(N__53441),
            .I(N__53075));
    InMux I__12321 (
            .O(N__53440),
            .I(N__53066));
    InMux I__12320 (
            .O(N__53439),
            .I(N__53066));
    InMux I__12319 (
            .O(N__53438),
            .I(N__53066));
    InMux I__12318 (
            .O(N__53437),
            .I(N__53066));
    InMux I__12317 (
            .O(N__53436),
            .I(N__53057));
    InMux I__12316 (
            .O(N__53435),
            .I(N__53057));
    InMux I__12315 (
            .O(N__53434),
            .I(N__53057));
    InMux I__12314 (
            .O(N__53433),
            .I(N__53057));
    InMux I__12313 (
            .O(N__53432),
            .I(N__53048));
    InMux I__12312 (
            .O(N__53429),
            .I(N__53048));
    InMux I__12311 (
            .O(N__53426),
            .I(N__53048));
    InMux I__12310 (
            .O(N__53425),
            .I(N__53048));
    InMux I__12309 (
            .O(N__53422),
            .I(N__53041));
    InMux I__12308 (
            .O(N__53419),
            .I(N__53041));
    InMux I__12307 (
            .O(N__53418),
            .I(N__53041));
    InMux I__12306 (
            .O(N__53417),
            .I(N__53032));
    InMux I__12305 (
            .O(N__53414),
            .I(N__53032));
    InMux I__12304 (
            .O(N__53413),
            .I(N__53032));
    InMux I__12303 (
            .O(N__53412),
            .I(N__53032));
    CascadeMux I__12302 (
            .O(N__53411),
            .I(N__53025));
    Span4Mux_s2_v I__12301 (
            .O(N__53406),
            .I(N__53022));
    LocalMux I__12300 (
            .O(N__53399),
            .I(N__53017));
    LocalMux I__12299 (
            .O(N__53388),
            .I(N__53017));
    CascadeMux I__12298 (
            .O(N__53387),
            .I(N__53013));
    CascadeMux I__12297 (
            .O(N__53386),
            .I(N__53009));
    CascadeMux I__12296 (
            .O(N__53385),
            .I(N__53005));
    Span4Mux_s3_v I__12295 (
            .O(N__53380),
            .I(N__52993));
    Span4Mux_s2_h I__12294 (
            .O(N__53377),
            .I(N__52993));
    LocalMux I__12293 (
            .O(N__53370),
            .I(N__52993));
    Span4Mux_s3_v I__12292 (
            .O(N__53359),
            .I(N__52986));
    LocalMux I__12291 (
            .O(N__53356),
            .I(N__52986));
    LocalMux I__12290 (
            .O(N__53349),
            .I(N__52986));
    LocalMux I__12289 (
            .O(N__53340),
            .I(N__52983));
    CascadeMux I__12288 (
            .O(N__53339),
            .I(N__52976));
    LocalMux I__12287 (
            .O(N__53330),
            .I(N__52966));
    LocalMux I__12286 (
            .O(N__53319),
            .I(N__52966));
    LocalMux I__12285 (
            .O(N__53310),
            .I(N__52957));
    LocalMux I__12284 (
            .O(N__53301),
            .I(N__52957));
    LocalMux I__12283 (
            .O(N__53292),
            .I(N__52957));
    LocalMux I__12282 (
            .O(N__53285),
            .I(N__52957));
    InMux I__12281 (
            .O(N__53282),
            .I(N__52954));
    InMux I__12280 (
            .O(N__53279),
            .I(N__52947));
    InMux I__12279 (
            .O(N__53276),
            .I(N__52947));
    InMux I__12278 (
            .O(N__53273),
            .I(N__52947));
    LocalMux I__12277 (
            .O(N__53268),
            .I(N__52942));
    LocalMux I__12276 (
            .O(N__53255),
            .I(N__52942));
    InMux I__12275 (
            .O(N__53254),
            .I(N__52939));
    InMux I__12274 (
            .O(N__53253),
            .I(N__52932));
    InMux I__12273 (
            .O(N__53252),
            .I(N__52932));
    InMux I__12272 (
            .O(N__53251),
            .I(N__52932));
    LocalMux I__12271 (
            .O(N__53248),
            .I(N__52927));
    LocalMux I__12270 (
            .O(N__53241),
            .I(N__52927));
    LocalMux I__12269 (
            .O(N__53234),
            .I(N__52922));
    LocalMux I__12268 (
            .O(N__53229),
            .I(N__52922));
    Span4Mux_h I__12267 (
            .O(N__53220),
            .I(N__52915));
    LocalMux I__12266 (
            .O(N__53213),
            .I(N__52915));
    LocalMux I__12265 (
            .O(N__53202),
            .I(N__52915));
    InMux I__12264 (
            .O(N__53199),
            .I(N__52910));
    InMux I__12263 (
            .O(N__53198),
            .I(N__52910));
    InMux I__12262 (
            .O(N__53197),
            .I(N__52905));
    InMux I__12261 (
            .O(N__53196),
            .I(N__52905));
    CascadeMux I__12260 (
            .O(N__53195),
            .I(N__52887));
    CascadeMux I__12259 (
            .O(N__53194),
            .I(N__52883));
    CascadeMux I__12258 (
            .O(N__53193),
            .I(N__52880));
    CascadeMux I__12257 (
            .O(N__53192),
            .I(N__52877));
    CascadeMux I__12256 (
            .O(N__53191),
            .I(N__52874));
    CascadeMux I__12255 (
            .O(N__53190),
            .I(N__52871));
    CascadeMux I__12254 (
            .O(N__53189),
            .I(N__52868));
    CascadeMux I__12253 (
            .O(N__53188),
            .I(N__52865));
    CascadeMux I__12252 (
            .O(N__53187),
            .I(N__52862));
    LocalMux I__12251 (
            .O(N__53180),
            .I(N__52855));
    LocalMux I__12250 (
            .O(N__53169),
            .I(N__52855));
    LocalMux I__12249 (
            .O(N__53164),
            .I(N__52855));
    InMux I__12248 (
            .O(N__53161),
            .I(N__52846));
    InMux I__12247 (
            .O(N__53160),
            .I(N__52846));
    InMux I__12246 (
            .O(N__53159),
            .I(N__52846));
    InMux I__12245 (
            .O(N__53158),
            .I(N__52846));
    InMux I__12244 (
            .O(N__53155),
            .I(N__52837));
    InMux I__12243 (
            .O(N__53154),
            .I(N__52837));
    InMux I__12242 (
            .O(N__53153),
            .I(N__52837));
    InMux I__12241 (
            .O(N__53152),
            .I(N__52837));
    Span4Mux_h I__12240 (
            .O(N__53149),
            .I(N__52832));
    LocalMux I__12239 (
            .O(N__53144),
            .I(N__52832));
    Span4Mux_v I__12238 (
            .O(N__53141),
            .I(N__52821));
    Span4Mux_v I__12237 (
            .O(N__53128),
            .I(N__52821));
    LocalMux I__12236 (
            .O(N__53121),
            .I(N__52821));
    Span4Mux_v I__12235 (
            .O(N__53116),
            .I(N__52821));
    Span4Mux_v I__12234 (
            .O(N__53109),
            .I(N__52821));
    LocalMux I__12233 (
            .O(N__53104),
            .I(N__52818));
    InMux I__12232 (
            .O(N__53103),
            .I(N__52811));
    InMux I__12231 (
            .O(N__53102),
            .I(N__52811));
    InMux I__12230 (
            .O(N__53101),
            .I(N__52811));
    InMux I__12229 (
            .O(N__53100),
            .I(N__52801));
    InMux I__12228 (
            .O(N__53099),
            .I(N__52801));
    InMux I__12227 (
            .O(N__53096),
            .I(N__52801));
    InMux I__12226 (
            .O(N__53095),
            .I(N__52801));
    InMux I__12225 (
            .O(N__53092),
            .I(N__52794));
    InMux I__12224 (
            .O(N__53091),
            .I(N__52794));
    InMux I__12223 (
            .O(N__53090),
            .I(N__52794));
    InMux I__12222 (
            .O(N__53087),
            .I(N__52787));
    InMux I__12221 (
            .O(N__53086),
            .I(N__52787));
    InMux I__12220 (
            .O(N__53085),
            .I(N__52787));
    LocalMux I__12219 (
            .O(N__53082),
            .I(N__52771));
    LocalMux I__12218 (
            .O(N__53075),
            .I(N__52771));
    LocalMux I__12217 (
            .O(N__53066),
            .I(N__52771));
    LocalMux I__12216 (
            .O(N__53057),
            .I(N__52771));
    LocalMux I__12215 (
            .O(N__53048),
            .I(N__52771));
    LocalMux I__12214 (
            .O(N__53041),
            .I(N__52771));
    LocalMux I__12213 (
            .O(N__53032),
            .I(N__52771));
    InMux I__12212 (
            .O(N__53031),
            .I(N__52768));
    InMux I__12211 (
            .O(N__53030),
            .I(N__52761));
    InMux I__12210 (
            .O(N__53029),
            .I(N__52761));
    InMux I__12209 (
            .O(N__53028),
            .I(N__52761));
    InMux I__12208 (
            .O(N__53025),
            .I(N__52758));
    Span4Mux_v I__12207 (
            .O(N__53022),
            .I(N__52753));
    Span4Mux_v I__12206 (
            .O(N__53017),
            .I(N__52753));
    InMux I__12205 (
            .O(N__53016),
            .I(N__52742));
    InMux I__12204 (
            .O(N__53013),
            .I(N__52742));
    InMux I__12203 (
            .O(N__53012),
            .I(N__52742));
    InMux I__12202 (
            .O(N__53009),
            .I(N__52742));
    InMux I__12201 (
            .O(N__53008),
            .I(N__52742));
    InMux I__12200 (
            .O(N__53005),
            .I(N__52735));
    InMux I__12199 (
            .O(N__53004),
            .I(N__52735));
    InMux I__12198 (
            .O(N__53003),
            .I(N__52735));
    CascadeMux I__12197 (
            .O(N__53002),
            .I(N__52727));
    CascadeMux I__12196 (
            .O(N__53001),
            .I(N__52718));
    CascadeMux I__12195 (
            .O(N__53000),
            .I(N__52714));
    Span4Mux_v I__12194 (
            .O(N__52993),
            .I(N__52704));
    Span4Mux_v I__12193 (
            .O(N__52986),
            .I(N__52704));
    Span4Mux_v I__12192 (
            .O(N__52983),
            .I(N__52704));
    InMux I__12191 (
            .O(N__52982),
            .I(N__52697));
    InMux I__12190 (
            .O(N__52981),
            .I(N__52697));
    InMux I__12189 (
            .O(N__52980),
            .I(N__52697));
    InMux I__12188 (
            .O(N__52979),
            .I(N__52694));
    InMux I__12187 (
            .O(N__52976),
            .I(N__52689));
    InMux I__12186 (
            .O(N__52975),
            .I(N__52689));
    InMux I__12185 (
            .O(N__52974),
            .I(N__52684));
    InMux I__12184 (
            .O(N__52973),
            .I(N__52684));
    InMux I__12183 (
            .O(N__52972),
            .I(N__52679));
    InMux I__12182 (
            .O(N__52971),
            .I(N__52679));
    Span4Mux_s3_v I__12181 (
            .O(N__52966),
            .I(N__52672));
    Span4Mux_s3_v I__12180 (
            .O(N__52957),
            .I(N__52672));
    LocalMux I__12179 (
            .O(N__52954),
            .I(N__52672));
    LocalMux I__12178 (
            .O(N__52947),
            .I(N__52669));
    Span4Mux_s3_h I__12177 (
            .O(N__52942),
            .I(N__52662));
    LocalMux I__12176 (
            .O(N__52939),
            .I(N__52662));
    LocalMux I__12175 (
            .O(N__52932),
            .I(N__52662));
    Span4Mux_v I__12174 (
            .O(N__52927),
            .I(N__52651));
    Span4Mux_v I__12173 (
            .O(N__52922),
            .I(N__52651));
    Span4Mux_v I__12172 (
            .O(N__52915),
            .I(N__52651));
    LocalMux I__12171 (
            .O(N__52910),
            .I(N__52651));
    LocalMux I__12170 (
            .O(N__52905),
            .I(N__52651));
    InMux I__12169 (
            .O(N__52904),
            .I(N__52646));
    InMux I__12168 (
            .O(N__52903),
            .I(N__52646));
    InMux I__12167 (
            .O(N__52902),
            .I(N__52641));
    InMux I__12166 (
            .O(N__52901),
            .I(N__52641));
    InMux I__12165 (
            .O(N__52900),
            .I(N__52634));
    InMux I__12164 (
            .O(N__52899),
            .I(N__52634));
    InMux I__12163 (
            .O(N__52898),
            .I(N__52634));
    InMux I__12162 (
            .O(N__52897),
            .I(N__52631));
    InMux I__12161 (
            .O(N__52896),
            .I(N__52624));
    InMux I__12160 (
            .O(N__52895),
            .I(N__52624));
    InMux I__12159 (
            .O(N__52894),
            .I(N__52624));
    InMux I__12158 (
            .O(N__52893),
            .I(N__52619));
    InMux I__12157 (
            .O(N__52892),
            .I(N__52619));
    InMux I__12156 (
            .O(N__52891),
            .I(N__52616));
    InMux I__12155 (
            .O(N__52890),
            .I(N__52609));
    InMux I__12154 (
            .O(N__52887),
            .I(N__52609));
    InMux I__12153 (
            .O(N__52886),
            .I(N__52609));
    InMux I__12152 (
            .O(N__52883),
            .I(N__52600));
    InMux I__12151 (
            .O(N__52880),
            .I(N__52600));
    InMux I__12150 (
            .O(N__52877),
            .I(N__52600));
    InMux I__12149 (
            .O(N__52874),
            .I(N__52600));
    InMux I__12148 (
            .O(N__52871),
            .I(N__52591));
    InMux I__12147 (
            .O(N__52868),
            .I(N__52591));
    InMux I__12146 (
            .O(N__52865),
            .I(N__52591));
    InMux I__12145 (
            .O(N__52862),
            .I(N__52591));
    Span4Mux_h I__12144 (
            .O(N__52855),
            .I(N__52583));
    LocalMux I__12143 (
            .O(N__52846),
            .I(N__52583));
    LocalMux I__12142 (
            .O(N__52837),
            .I(N__52583));
    Span4Mux_h I__12141 (
            .O(N__52832),
            .I(N__52576));
    Span4Mux_h I__12140 (
            .O(N__52821),
            .I(N__52576));
    Span4Mux_v I__12139 (
            .O(N__52818),
            .I(N__52576));
    LocalMux I__12138 (
            .O(N__52811),
            .I(N__52573));
    InMux I__12137 (
            .O(N__52810),
            .I(N__52570));
    LocalMux I__12136 (
            .O(N__52801),
            .I(N__52563));
    LocalMux I__12135 (
            .O(N__52794),
            .I(N__52563));
    LocalMux I__12134 (
            .O(N__52787),
            .I(N__52563));
    InMux I__12133 (
            .O(N__52786),
            .I(N__52560));
    Span12Mux_v I__12132 (
            .O(N__52771),
            .I(N__52542));
    LocalMux I__12131 (
            .O(N__52768),
            .I(N__52542));
    LocalMux I__12130 (
            .O(N__52761),
            .I(N__52542));
    LocalMux I__12129 (
            .O(N__52758),
            .I(N__52542));
    Sp12to4 I__12128 (
            .O(N__52753),
            .I(N__52542));
    LocalMux I__12127 (
            .O(N__52742),
            .I(N__52542));
    LocalMux I__12126 (
            .O(N__52735),
            .I(N__52542));
    InMux I__12125 (
            .O(N__52734),
            .I(N__52539));
    InMux I__12124 (
            .O(N__52733),
            .I(N__52532));
    InMux I__12123 (
            .O(N__52732),
            .I(N__52532));
    InMux I__12122 (
            .O(N__52731),
            .I(N__52532));
    InMux I__12121 (
            .O(N__52730),
            .I(N__52521));
    InMux I__12120 (
            .O(N__52727),
            .I(N__52521));
    InMux I__12119 (
            .O(N__52726),
            .I(N__52521));
    InMux I__12118 (
            .O(N__52725),
            .I(N__52521));
    InMux I__12117 (
            .O(N__52724),
            .I(N__52521));
    InMux I__12116 (
            .O(N__52723),
            .I(N__52514));
    InMux I__12115 (
            .O(N__52722),
            .I(N__52514));
    InMux I__12114 (
            .O(N__52721),
            .I(N__52514));
    InMux I__12113 (
            .O(N__52718),
            .I(N__52505));
    InMux I__12112 (
            .O(N__52717),
            .I(N__52505));
    InMux I__12111 (
            .O(N__52714),
            .I(N__52505));
    InMux I__12110 (
            .O(N__52713),
            .I(N__52505));
    InMux I__12109 (
            .O(N__52712),
            .I(N__52500));
    InMux I__12108 (
            .O(N__52711),
            .I(N__52500));
    Span4Mux_h I__12107 (
            .O(N__52704),
            .I(N__52497));
    LocalMux I__12106 (
            .O(N__52697),
            .I(N__52494));
    LocalMux I__12105 (
            .O(N__52694),
            .I(N__52485));
    LocalMux I__12104 (
            .O(N__52689),
            .I(N__52485));
    LocalMux I__12103 (
            .O(N__52684),
            .I(N__52485));
    LocalMux I__12102 (
            .O(N__52679),
            .I(N__52485));
    Span4Mux_v I__12101 (
            .O(N__52672),
            .I(N__52478));
    Span4Mux_v I__12100 (
            .O(N__52669),
            .I(N__52478));
    Span4Mux_h I__12099 (
            .O(N__52662),
            .I(N__52478));
    Span4Mux_h I__12098 (
            .O(N__52651),
            .I(N__52471));
    LocalMux I__12097 (
            .O(N__52646),
            .I(N__52471));
    LocalMux I__12096 (
            .O(N__52641),
            .I(N__52471));
    LocalMux I__12095 (
            .O(N__52634),
            .I(N__52460));
    LocalMux I__12094 (
            .O(N__52631),
            .I(N__52460));
    LocalMux I__12093 (
            .O(N__52624),
            .I(N__52460));
    LocalMux I__12092 (
            .O(N__52619),
            .I(N__52460));
    LocalMux I__12091 (
            .O(N__52616),
            .I(N__52460));
    LocalMux I__12090 (
            .O(N__52609),
            .I(N__52453));
    LocalMux I__12089 (
            .O(N__52600),
            .I(N__52453));
    LocalMux I__12088 (
            .O(N__52591),
            .I(N__52453));
    InMux I__12087 (
            .O(N__52590),
            .I(N__52450));
    Span4Mux_h I__12086 (
            .O(N__52583),
            .I(N__52437));
    Span4Mux_h I__12085 (
            .O(N__52576),
            .I(N__52437));
    Span4Mux_v I__12084 (
            .O(N__52573),
            .I(N__52437));
    LocalMux I__12083 (
            .O(N__52570),
            .I(N__52437));
    Span4Mux_h I__12082 (
            .O(N__52563),
            .I(N__52437));
    LocalMux I__12081 (
            .O(N__52560),
            .I(N__52437));
    InMux I__12080 (
            .O(N__52559),
            .I(N__52430));
    InMux I__12079 (
            .O(N__52558),
            .I(N__52430));
    InMux I__12078 (
            .O(N__52557),
            .I(N__52430));
    Span12Mux_h I__12077 (
            .O(N__52542),
            .I(N__52412));
    LocalMux I__12076 (
            .O(N__52539),
            .I(N__52412));
    LocalMux I__12075 (
            .O(N__52532),
            .I(N__52412));
    LocalMux I__12074 (
            .O(N__52521),
            .I(N__52412));
    LocalMux I__12073 (
            .O(N__52514),
            .I(N__52412));
    LocalMux I__12072 (
            .O(N__52505),
            .I(N__52412));
    LocalMux I__12071 (
            .O(N__52500),
            .I(N__52412));
    Span4Mux_h I__12070 (
            .O(N__52497),
            .I(N__52405));
    Span4Mux_v I__12069 (
            .O(N__52494),
            .I(N__52405));
    Span4Mux_v I__12068 (
            .O(N__52485),
            .I(N__52405));
    Span4Mux_h I__12067 (
            .O(N__52478),
            .I(N__52398));
    Span4Mux_v I__12066 (
            .O(N__52471),
            .I(N__52398));
    Span4Mux_v I__12065 (
            .O(N__52460),
            .I(N__52398));
    Span12Mux_h I__12064 (
            .O(N__52453),
            .I(N__52393));
    LocalMux I__12063 (
            .O(N__52450),
            .I(N__52393));
    Span4Mux_v I__12062 (
            .O(N__52437),
            .I(N__52388));
    LocalMux I__12061 (
            .O(N__52430),
            .I(N__52388));
    InMux I__12060 (
            .O(N__52429),
            .I(N__52385));
    InMux I__12059 (
            .O(N__52428),
            .I(N__52380));
    InMux I__12058 (
            .O(N__52427),
            .I(N__52380));
    Odrv12 I__12057 (
            .O(N__52412),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12056 (
            .O(N__52405),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12055 (
            .O(N__52398),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__12054 (
            .O(N__52393),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12053 (
            .O(N__52388),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12052 (
            .O(N__52385),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12051 (
            .O(N__52380),
            .I(CONSTANT_ONE_NET));
    InMux I__12050 (
            .O(N__52365),
            .I(N__52362));
    LocalMux I__12049 (
            .O(N__52362),
            .I(N__52359));
    Span4Mux_v I__12048 (
            .O(N__52359),
            .I(N__52356));
    Sp12to4 I__12047 (
            .O(N__52356),
            .I(N__52352));
    InMux I__12046 (
            .O(N__52355),
            .I(N__52349));
    Odrv12 I__12045 (
            .O(N__52352),
            .I(n15513));
    LocalMux I__12044 (
            .O(N__52349),
            .I(n15513));
    CascadeMux I__12043 (
            .O(N__52344),
            .I(N__52341));
    InMux I__12042 (
            .O(N__52341),
            .I(N__52338));
    LocalMux I__12041 (
            .O(N__52338),
            .I(N__52334));
    InMux I__12040 (
            .O(N__52337),
            .I(N__52331));
    Odrv4 I__12039 (
            .O(N__52334),
            .I(n1125));
    LocalMux I__12038 (
            .O(N__52331),
            .I(n1125));
    InMux I__12037 (
            .O(N__52326),
            .I(n12516));
    CascadeMux I__12036 (
            .O(N__52323),
            .I(N__52319));
    InMux I__12035 (
            .O(N__52322),
            .I(N__52316));
    InMux I__12034 (
            .O(N__52319),
            .I(N__52313));
    LocalMux I__12033 (
            .O(N__52316),
            .I(N__52310));
    LocalMux I__12032 (
            .O(N__52313),
            .I(n1224));
    Odrv4 I__12031 (
            .O(N__52310),
            .I(n1224));
    CascadeMux I__12030 (
            .O(N__52305),
            .I(N__52301));
    InMux I__12029 (
            .O(N__52304),
            .I(N__52296));
    InMux I__12028 (
            .O(N__52301),
            .I(N__52296));
    LocalMux I__12027 (
            .O(N__52296),
            .I(N__52293));
    Span4Mux_h I__12026 (
            .O(N__52293),
            .I(N__52290));
    Odrv4 I__12025 (
            .O(N__52290),
            .I(n1126));
    CascadeMux I__12024 (
            .O(N__52287),
            .I(N__52284));
    InMux I__12023 (
            .O(N__52284),
            .I(N__52281));
    LocalMux I__12022 (
            .O(N__52281),
            .I(n1193));
    CascadeMux I__12021 (
            .O(N__52278),
            .I(N__52271));
    CascadeMux I__12020 (
            .O(N__52277),
            .I(N__52268));
    CascadeMux I__12019 (
            .O(N__52276),
            .I(N__52265));
    InMux I__12018 (
            .O(N__52275),
            .I(N__52261));
    InMux I__12017 (
            .O(N__52274),
            .I(N__52258));
    InMux I__12016 (
            .O(N__52271),
            .I(N__52249));
    InMux I__12015 (
            .O(N__52268),
            .I(N__52249));
    InMux I__12014 (
            .O(N__52265),
            .I(N__52249));
    InMux I__12013 (
            .O(N__52264),
            .I(N__52249));
    LocalMux I__12012 (
            .O(N__52261),
            .I(N__52246));
    LocalMux I__12011 (
            .O(N__52258),
            .I(N__52242));
    LocalMux I__12010 (
            .O(N__52249),
            .I(N__52236));
    Span12Mux_s9_v I__12009 (
            .O(N__52246),
            .I(N__52233));
    InMux I__12008 (
            .O(N__52245),
            .I(N__52230));
    Span4Mux_h I__12007 (
            .O(N__52242),
            .I(N__52227));
    InMux I__12006 (
            .O(N__52241),
            .I(N__52224));
    InMux I__12005 (
            .O(N__52240),
            .I(N__52221));
    InMux I__12004 (
            .O(N__52239),
            .I(N__52218));
    Span4Mux_h I__12003 (
            .O(N__52236),
            .I(N__52215));
    Odrv12 I__12002 (
            .O(N__52233),
            .I(n1158));
    LocalMux I__12001 (
            .O(N__52230),
            .I(n1158));
    Odrv4 I__12000 (
            .O(N__52227),
            .I(n1158));
    LocalMux I__11999 (
            .O(N__52224),
            .I(n1158));
    LocalMux I__11998 (
            .O(N__52221),
            .I(n1158));
    LocalMux I__11997 (
            .O(N__52218),
            .I(n1158));
    Odrv4 I__11996 (
            .O(N__52215),
            .I(n1158));
    InMux I__11995 (
            .O(N__52200),
            .I(N__52197));
    LocalMux I__11994 (
            .O(N__52197),
            .I(N__52192));
    CascadeMux I__11993 (
            .O(N__52196),
            .I(N__52189));
    InMux I__11992 (
            .O(N__52195),
            .I(N__52186));
    Span4Mux_h I__11991 (
            .O(N__52192),
            .I(N__52183));
    InMux I__11990 (
            .O(N__52189),
            .I(N__52180));
    LocalMux I__11989 (
            .O(N__52186),
            .I(N__52177));
    Odrv4 I__11988 (
            .O(N__52183),
            .I(n1225));
    LocalMux I__11987 (
            .O(N__52180),
            .I(n1225));
    Odrv12 I__11986 (
            .O(N__52177),
            .I(n1225));
    InMux I__11985 (
            .O(N__52170),
            .I(N__52167));
    LocalMux I__11984 (
            .O(N__52167),
            .I(N__52164));
    Odrv12 I__11983 (
            .O(N__52164),
            .I(n23_adj_700));
    CascadeMux I__11982 (
            .O(N__52161),
            .I(N__52158));
    InMux I__11981 (
            .O(N__52158),
            .I(N__52155));
    LocalMux I__11980 (
            .O(N__52155),
            .I(N__52152));
    Odrv4 I__11979 (
            .O(N__52152),
            .I(n25_adj_698));
    CascadeMux I__11978 (
            .O(N__52149),
            .I(direction_N_342_cascade_));
    CascadeMux I__11977 (
            .O(N__52146),
            .I(N__52143));
    InMux I__11976 (
            .O(N__52143),
            .I(N__52140));
    LocalMux I__11975 (
            .O(N__52140),
            .I(n1693));
    InMux I__11974 (
            .O(N__52137),
            .I(N__52133));
    InMux I__11973 (
            .O(N__52136),
            .I(N__52130));
    LocalMux I__11972 (
            .O(N__52133),
            .I(N__52125));
    LocalMux I__11971 (
            .O(N__52130),
            .I(N__52125));
    Span4Mux_h I__11970 (
            .O(N__52125),
            .I(N__52122));
    Odrv4 I__11969 (
            .O(N__52122),
            .I(direction_N_340));
    InMux I__11968 (
            .O(N__52119),
            .I(N__52116));
    LocalMux I__11967 (
            .O(N__52116),
            .I(direction_N_342));
    CascadeMux I__11966 (
            .O(N__52113),
            .I(n13661_cascade_));
    InMux I__11965 (
            .O(N__52110),
            .I(N__52103));
    CascadeMux I__11964 (
            .O(N__52109),
            .I(N__52100));
    CascadeMux I__11963 (
            .O(N__52108),
            .I(N__52096));
    CascadeMux I__11962 (
            .O(N__52107),
            .I(N__52092));
    CascadeMux I__11961 (
            .O(N__52106),
            .I(N__52088));
    LocalMux I__11960 (
            .O(N__52103),
            .I(N__52078));
    InMux I__11959 (
            .O(N__52100),
            .I(N__52061));
    InMux I__11958 (
            .O(N__52099),
            .I(N__52061));
    InMux I__11957 (
            .O(N__52096),
            .I(N__52061));
    InMux I__11956 (
            .O(N__52095),
            .I(N__52061));
    InMux I__11955 (
            .O(N__52092),
            .I(N__52061));
    InMux I__11954 (
            .O(N__52091),
            .I(N__52061));
    InMux I__11953 (
            .O(N__52088),
            .I(N__52061));
    InMux I__11952 (
            .O(N__52087),
            .I(N__52061));
    CascadeMux I__11951 (
            .O(N__52086),
            .I(N__52058));
    CascadeMux I__11950 (
            .O(N__52085),
            .I(N__52054));
    CascadeMux I__11949 (
            .O(N__52084),
            .I(N__52050));
    CascadeMux I__11948 (
            .O(N__52083),
            .I(N__52046));
    CascadeMux I__11947 (
            .O(N__52082),
            .I(N__52039));
    InMux I__11946 (
            .O(N__52081),
            .I(N__52030));
    Span4Mux_v I__11945 (
            .O(N__52078),
            .I(N__52025));
    LocalMux I__11944 (
            .O(N__52061),
            .I(N__52025));
    InMux I__11943 (
            .O(N__52058),
            .I(N__52008));
    InMux I__11942 (
            .O(N__52057),
            .I(N__52008));
    InMux I__11941 (
            .O(N__52054),
            .I(N__52008));
    InMux I__11940 (
            .O(N__52053),
            .I(N__52008));
    InMux I__11939 (
            .O(N__52050),
            .I(N__52008));
    InMux I__11938 (
            .O(N__52049),
            .I(N__52008));
    InMux I__11937 (
            .O(N__52046),
            .I(N__52008));
    InMux I__11936 (
            .O(N__52045),
            .I(N__52008));
    InMux I__11935 (
            .O(N__52044),
            .I(N__51999));
    InMux I__11934 (
            .O(N__52043),
            .I(N__51999));
    InMux I__11933 (
            .O(N__52042),
            .I(N__51999));
    InMux I__11932 (
            .O(N__52039),
            .I(N__51999));
    InMux I__11931 (
            .O(N__52038),
            .I(N__51990));
    InMux I__11930 (
            .O(N__52037),
            .I(N__51990));
    InMux I__11929 (
            .O(N__52036),
            .I(N__51990));
    InMux I__11928 (
            .O(N__52035),
            .I(N__51990));
    InMux I__11927 (
            .O(N__52034),
            .I(N__51985));
    InMux I__11926 (
            .O(N__52033),
            .I(N__51985));
    LocalMux I__11925 (
            .O(N__52030),
            .I(direction_c));
    Odrv4 I__11924 (
            .O(N__52025),
            .I(direction_c));
    LocalMux I__11923 (
            .O(N__52008),
            .I(direction_c));
    LocalMux I__11922 (
            .O(N__51999),
            .I(direction_c));
    LocalMux I__11921 (
            .O(N__51990),
            .I(direction_c));
    LocalMux I__11920 (
            .O(N__51985),
            .I(direction_c));
    CascadeMux I__11919 (
            .O(N__51972),
            .I(n22_adj_705_cascade_));
    InMux I__11918 (
            .O(N__51969),
            .I(N__51966));
    LocalMux I__11917 (
            .O(N__51966),
            .I(N__51963));
    Odrv4 I__11916 (
            .O(N__51963),
            .I(n1200));
    InMux I__11915 (
            .O(N__51960),
            .I(n12508));
    InMux I__11914 (
            .O(N__51957),
            .I(N__51954));
    LocalMux I__11913 (
            .O(N__51954),
            .I(N__51950));
    InMux I__11912 (
            .O(N__51953),
            .I(N__51947));
    Span4Mux_v I__11911 (
            .O(N__51950),
            .I(N__51944));
    LocalMux I__11910 (
            .O(N__51947),
            .I(n1132));
    Odrv4 I__11909 (
            .O(N__51944),
            .I(n1132));
    InMux I__11908 (
            .O(N__51939),
            .I(N__51936));
    LocalMux I__11907 (
            .O(N__51936),
            .I(N__51933));
    Span4Mux_h I__11906 (
            .O(N__51933),
            .I(N__51930));
    Odrv4 I__11905 (
            .O(N__51930),
            .I(n1199));
    InMux I__11904 (
            .O(N__51927),
            .I(n12509));
    CascadeMux I__11903 (
            .O(N__51924),
            .I(N__51921));
    InMux I__11902 (
            .O(N__51921),
            .I(N__51917));
    InMux I__11901 (
            .O(N__51920),
            .I(N__51914));
    LocalMux I__11900 (
            .O(N__51917),
            .I(N__51910));
    LocalMux I__11899 (
            .O(N__51914),
            .I(N__51907));
    InMux I__11898 (
            .O(N__51913),
            .I(N__51904));
    Span4Mux_h I__11897 (
            .O(N__51910),
            .I(N__51901));
    Odrv4 I__11896 (
            .O(N__51907),
            .I(n1131));
    LocalMux I__11895 (
            .O(N__51904),
            .I(n1131));
    Odrv4 I__11894 (
            .O(N__51901),
            .I(n1131));
    CascadeMux I__11893 (
            .O(N__51894),
            .I(N__51891));
    InMux I__11892 (
            .O(N__51891),
            .I(N__51888));
    LocalMux I__11891 (
            .O(N__51888),
            .I(n1198));
    InMux I__11890 (
            .O(N__51885),
            .I(n12510));
    InMux I__11889 (
            .O(N__51882),
            .I(N__51878));
    CascadeMux I__11888 (
            .O(N__51881),
            .I(N__51875));
    LocalMux I__11887 (
            .O(N__51878),
            .I(N__51871));
    InMux I__11886 (
            .O(N__51875),
            .I(N__51868));
    CascadeMux I__11885 (
            .O(N__51874),
            .I(N__51865));
    Span4Mux_v I__11884 (
            .O(N__51871),
            .I(N__51860));
    LocalMux I__11883 (
            .O(N__51868),
            .I(N__51860));
    InMux I__11882 (
            .O(N__51865),
            .I(N__51857));
    Odrv4 I__11881 (
            .O(N__51860),
            .I(n1130));
    LocalMux I__11880 (
            .O(N__51857),
            .I(n1130));
    InMux I__11879 (
            .O(N__51852),
            .I(N__51849));
    LocalMux I__11878 (
            .O(N__51849),
            .I(n1197));
    InMux I__11877 (
            .O(N__51846),
            .I(n12511));
    InMux I__11876 (
            .O(N__51843),
            .I(N__51839));
    CascadeMux I__11875 (
            .O(N__51842),
            .I(N__51836));
    LocalMux I__11874 (
            .O(N__51839),
            .I(N__51833));
    InMux I__11873 (
            .O(N__51836),
            .I(N__51830));
    Span4Mux_v I__11872 (
            .O(N__51833),
            .I(N__51825));
    LocalMux I__11871 (
            .O(N__51830),
            .I(N__51825));
    Span4Mux_h I__11870 (
            .O(N__51825),
            .I(N__51821));
    InMux I__11869 (
            .O(N__51824),
            .I(N__51818));
    Odrv4 I__11868 (
            .O(N__51821),
            .I(n1129));
    LocalMux I__11867 (
            .O(N__51818),
            .I(n1129));
    InMux I__11866 (
            .O(N__51813),
            .I(N__51810));
    LocalMux I__11865 (
            .O(N__51810),
            .I(n1196));
    InMux I__11864 (
            .O(N__51807),
            .I(n12512));
    CascadeMux I__11863 (
            .O(N__51804),
            .I(N__51800));
    CascadeMux I__11862 (
            .O(N__51803),
            .I(N__51797));
    InMux I__11861 (
            .O(N__51800),
            .I(N__51794));
    InMux I__11860 (
            .O(N__51797),
            .I(N__51791));
    LocalMux I__11859 (
            .O(N__51794),
            .I(N__51788));
    LocalMux I__11858 (
            .O(N__51791),
            .I(N__51784));
    Span4Mux_h I__11857 (
            .O(N__51788),
            .I(N__51781));
    InMux I__11856 (
            .O(N__51787),
            .I(N__51778));
    Odrv12 I__11855 (
            .O(N__51784),
            .I(n1128));
    Odrv4 I__11854 (
            .O(N__51781),
            .I(n1128));
    LocalMux I__11853 (
            .O(N__51778),
            .I(n1128));
    InMux I__11852 (
            .O(N__51771),
            .I(N__51768));
    LocalMux I__11851 (
            .O(N__51768),
            .I(n1195));
    InMux I__11850 (
            .O(N__51765),
            .I(n12513));
    InMux I__11849 (
            .O(N__51762),
            .I(N__51758));
    CascadeMux I__11848 (
            .O(N__51761),
            .I(N__51755));
    LocalMux I__11847 (
            .O(N__51758),
            .I(N__51752));
    InMux I__11846 (
            .O(N__51755),
            .I(N__51749));
    Span4Mux_h I__11845 (
            .O(N__51752),
            .I(N__51745));
    LocalMux I__11844 (
            .O(N__51749),
            .I(N__51742));
    InMux I__11843 (
            .O(N__51748),
            .I(N__51739));
    Odrv4 I__11842 (
            .O(N__51745),
            .I(n1127));
    Odrv12 I__11841 (
            .O(N__51742),
            .I(n1127));
    LocalMux I__11840 (
            .O(N__51739),
            .I(n1127));
    InMux I__11839 (
            .O(N__51732),
            .I(N__51729));
    LocalMux I__11838 (
            .O(N__51729),
            .I(n1194));
    InMux I__11837 (
            .O(N__51726),
            .I(n12514));
    InMux I__11836 (
            .O(N__51723),
            .I(bfn_16_24_0_));
    CascadeMux I__11835 (
            .O(N__51720),
            .I(N__51716));
    CascadeMux I__11834 (
            .O(N__51719),
            .I(N__51713));
    InMux I__11833 (
            .O(N__51716),
            .I(N__51710));
    InMux I__11832 (
            .O(N__51713),
            .I(N__51707));
    LocalMux I__11831 (
            .O(N__51710),
            .I(N__51704));
    LocalMux I__11830 (
            .O(N__51707),
            .I(n1226));
    Odrv4 I__11829 (
            .O(N__51704),
            .I(n1226));
    CascadeMux I__11828 (
            .O(N__51699),
            .I(n1226_cascade_));
    InMux I__11827 (
            .O(N__51696),
            .I(N__51693));
    LocalMux I__11826 (
            .O(N__51693),
            .I(N__51690));
    Odrv4 I__11825 (
            .O(N__51690),
            .I(n1293));
    CascadeMux I__11824 (
            .O(N__51687),
            .I(N__51684));
    InMux I__11823 (
            .O(N__51684),
            .I(N__51679));
    InMux I__11822 (
            .O(N__51683),
            .I(N__51674));
    InMux I__11821 (
            .O(N__51682),
            .I(N__51674));
    LocalMux I__11820 (
            .O(N__51679),
            .I(n1325));
    LocalMux I__11819 (
            .O(N__51674),
            .I(n1325));
    CascadeMux I__11818 (
            .O(N__51669),
            .I(N__51665));
    InMux I__11817 (
            .O(N__51668),
            .I(N__51662));
    InMux I__11816 (
            .O(N__51665),
            .I(N__51659));
    LocalMux I__11815 (
            .O(N__51662),
            .I(n1229));
    LocalMux I__11814 (
            .O(N__51659),
            .I(n1229));
    InMux I__11813 (
            .O(N__51654),
            .I(N__51651));
    LocalMux I__11812 (
            .O(N__51651),
            .I(N__51648));
    Span4Mux_h I__11811 (
            .O(N__51648),
            .I(N__51645));
    Odrv4 I__11810 (
            .O(N__51645),
            .I(n11910));
    CascadeMux I__11809 (
            .O(N__51642),
            .I(n1229_cascade_));
    InMux I__11808 (
            .O(N__51639),
            .I(N__51634));
    InMux I__11807 (
            .O(N__51638),
            .I(N__51631));
    CascadeMux I__11806 (
            .O(N__51637),
            .I(N__51628));
    LocalMux I__11805 (
            .O(N__51634),
            .I(N__51625));
    LocalMux I__11804 (
            .O(N__51631),
            .I(N__51622));
    InMux I__11803 (
            .O(N__51628),
            .I(N__51619));
    Span4Mux_h I__11802 (
            .O(N__51625),
            .I(N__51616));
    Odrv4 I__11801 (
            .O(N__51622),
            .I(n1231));
    LocalMux I__11800 (
            .O(N__51619),
            .I(n1231));
    Odrv4 I__11799 (
            .O(N__51616),
            .I(n1231));
    InMux I__11798 (
            .O(N__51609),
            .I(N__51606));
    LocalMux I__11797 (
            .O(N__51606),
            .I(n13711));
    InMux I__11796 (
            .O(N__51603),
            .I(N__51598));
    CascadeMux I__11795 (
            .O(N__51602),
            .I(N__51594));
    CascadeMux I__11794 (
            .O(N__51601),
            .I(N__51591));
    LocalMux I__11793 (
            .O(N__51598),
            .I(N__51586));
    CascadeMux I__11792 (
            .O(N__51597),
            .I(N__51583));
    InMux I__11791 (
            .O(N__51594),
            .I(N__51576));
    InMux I__11790 (
            .O(N__51591),
            .I(N__51576));
    InMux I__11789 (
            .O(N__51590),
            .I(N__51573));
    CascadeMux I__11788 (
            .O(N__51589),
            .I(N__51570));
    Span12Mux_h I__11787 (
            .O(N__51586),
            .I(N__51564));
    InMux I__11786 (
            .O(N__51583),
            .I(N__51557));
    InMux I__11785 (
            .O(N__51582),
            .I(N__51557));
    InMux I__11784 (
            .O(N__51581),
            .I(N__51557));
    LocalMux I__11783 (
            .O(N__51576),
            .I(N__51552));
    LocalMux I__11782 (
            .O(N__51573),
            .I(N__51552));
    InMux I__11781 (
            .O(N__51570),
            .I(N__51547));
    InMux I__11780 (
            .O(N__51569),
            .I(N__51547));
    InMux I__11779 (
            .O(N__51568),
            .I(N__51542));
    InMux I__11778 (
            .O(N__51567),
            .I(N__51542));
    Odrv12 I__11777 (
            .O(N__51564),
            .I(n1257));
    LocalMux I__11776 (
            .O(N__51557),
            .I(n1257));
    Odrv4 I__11775 (
            .O(N__51552),
            .I(n1257));
    LocalMux I__11774 (
            .O(N__51547),
            .I(n1257));
    LocalMux I__11773 (
            .O(N__51542),
            .I(n1257));
    InMux I__11772 (
            .O(N__51531),
            .I(N__51528));
    LocalMux I__11771 (
            .O(N__51528),
            .I(N__51525));
    Span4Mux_h I__11770 (
            .O(N__51525),
            .I(N__51522));
    Span4Mux_h I__11769 (
            .O(N__51522),
            .I(N__51518));
    InMux I__11768 (
            .O(N__51521),
            .I(N__51515));
    Span4Mux_h I__11767 (
            .O(N__51518),
            .I(N__51510));
    LocalMux I__11766 (
            .O(N__51515),
            .I(N__51510));
    Odrv4 I__11765 (
            .O(N__51510),
            .I(n15528));
    CascadeMux I__11764 (
            .O(N__51507),
            .I(N__51502));
    InMux I__11763 (
            .O(N__51506),
            .I(N__51497));
    InMux I__11762 (
            .O(N__51505),
            .I(N__51497));
    InMux I__11761 (
            .O(N__51502),
            .I(N__51494));
    LocalMux I__11760 (
            .O(N__51497),
            .I(n1228));
    LocalMux I__11759 (
            .O(N__51494),
            .I(n1228));
    CascadeMux I__11758 (
            .O(N__51489),
            .I(N__51484));
    InMux I__11757 (
            .O(N__51488),
            .I(N__51481));
    InMux I__11756 (
            .O(N__51487),
            .I(N__51478));
    InMux I__11755 (
            .O(N__51484),
            .I(N__51475));
    LocalMux I__11754 (
            .O(N__51481),
            .I(n1230));
    LocalMux I__11753 (
            .O(N__51478),
            .I(n1230));
    LocalMux I__11752 (
            .O(N__51475),
            .I(n1230));
    CascadeMux I__11751 (
            .O(N__51468),
            .I(N__51465));
    InMux I__11750 (
            .O(N__51465),
            .I(N__51460));
    InMux I__11749 (
            .O(N__51464),
            .I(N__51455));
    InMux I__11748 (
            .O(N__51463),
            .I(N__51455));
    LocalMux I__11747 (
            .O(N__51460),
            .I(N__51452));
    LocalMux I__11746 (
            .O(N__51455),
            .I(N__51449));
    Span4Mux_h I__11745 (
            .O(N__51452),
            .I(N__51446));
    Odrv4 I__11744 (
            .O(N__51449),
            .I(n297));
    Odrv4 I__11743 (
            .O(N__51446),
            .I(n297));
    InMux I__11742 (
            .O(N__51441),
            .I(N__51438));
    LocalMux I__11741 (
            .O(N__51438),
            .I(N__51435));
    Odrv12 I__11740 (
            .O(N__51435),
            .I(n1201));
    InMux I__11739 (
            .O(N__51432),
            .I(bfn_16_23_0_));
    CascadeMux I__11738 (
            .O(N__51429),
            .I(N__51425));
    CascadeMux I__11737 (
            .O(N__51428),
            .I(N__51422));
    InMux I__11736 (
            .O(N__51425),
            .I(N__51419));
    InMux I__11735 (
            .O(N__51422),
            .I(N__51416));
    LocalMux I__11734 (
            .O(N__51419),
            .I(N__51413));
    LocalMux I__11733 (
            .O(N__51416),
            .I(N__51410));
    Odrv4 I__11732 (
            .O(N__51413),
            .I(n1133));
    Odrv4 I__11731 (
            .O(N__51410),
            .I(n1133));
    InMux I__11730 (
            .O(N__51405),
            .I(N__51402));
    LocalMux I__11729 (
            .O(N__51402),
            .I(N__51394));
    CascadeMux I__11728 (
            .O(N__51401),
            .I(N__51388));
    CascadeMux I__11727 (
            .O(N__51400),
            .I(N__51383));
    CascadeMux I__11726 (
            .O(N__51399),
            .I(N__51380));
    CascadeMux I__11725 (
            .O(N__51398),
            .I(N__51376));
    InMux I__11724 (
            .O(N__51397),
            .I(N__51372));
    Span12Mux_h I__11723 (
            .O(N__51394),
            .I(N__51369));
    InMux I__11722 (
            .O(N__51393),
            .I(N__51366));
    InMux I__11721 (
            .O(N__51392),
            .I(N__51363));
    InMux I__11720 (
            .O(N__51391),
            .I(N__51358));
    InMux I__11719 (
            .O(N__51388),
            .I(N__51358));
    InMux I__11718 (
            .O(N__51387),
            .I(N__51351));
    InMux I__11717 (
            .O(N__51386),
            .I(N__51351));
    InMux I__11716 (
            .O(N__51383),
            .I(N__51351));
    InMux I__11715 (
            .O(N__51380),
            .I(N__51342));
    InMux I__11714 (
            .O(N__51379),
            .I(N__51342));
    InMux I__11713 (
            .O(N__51376),
            .I(N__51342));
    InMux I__11712 (
            .O(N__51375),
            .I(N__51342));
    LocalMux I__11711 (
            .O(N__51372),
            .I(N__51339));
    Odrv12 I__11710 (
            .O(N__51369),
            .I(n1455));
    LocalMux I__11709 (
            .O(N__51366),
            .I(n1455));
    LocalMux I__11708 (
            .O(N__51363),
            .I(n1455));
    LocalMux I__11707 (
            .O(N__51358),
            .I(n1455));
    LocalMux I__11706 (
            .O(N__51351),
            .I(n1455));
    LocalMux I__11705 (
            .O(N__51342),
            .I(n1455));
    Odrv4 I__11704 (
            .O(N__51339),
            .I(n1455));
    InMux I__11703 (
            .O(N__51324),
            .I(N__51321));
    LocalMux I__11702 (
            .O(N__51321),
            .I(N__51318));
    Span12Mux_h I__11701 (
            .O(N__51318),
            .I(N__51314));
    InMux I__11700 (
            .O(N__51317),
            .I(N__51311));
    Odrv12 I__11699 (
            .O(N__51314),
            .I(n15562));
    LocalMux I__11698 (
            .O(N__51311),
            .I(n15562));
    InMux I__11697 (
            .O(N__51306),
            .I(N__51303));
    LocalMux I__11696 (
            .O(N__51303),
            .I(n1392));
    InMux I__11695 (
            .O(N__51300),
            .I(N__51297));
    LocalMux I__11694 (
            .O(N__51297),
            .I(N__51291));
    InMux I__11693 (
            .O(N__51296),
            .I(N__51288));
    CascadeMux I__11692 (
            .O(N__51295),
            .I(N__51284));
    InMux I__11691 (
            .O(N__51294),
            .I(N__51278));
    Span4Mux_h I__11690 (
            .O(N__51291),
            .I(N__51274));
    LocalMux I__11689 (
            .O(N__51288),
            .I(N__51271));
    CascadeMux I__11688 (
            .O(N__51287),
            .I(N__51267));
    InMux I__11687 (
            .O(N__51284),
            .I(N__51261));
    InMux I__11686 (
            .O(N__51283),
            .I(N__51261));
    InMux I__11685 (
            .O(N__51282),
            .I(N__51258));
    InMux I__11684 (
            .O(N__51281),
            .I(N__51255));
    LocalMux I__11683 (
            .O(N__51278),
            .I(N__51252));
    CascadeMux I__11682 (
            .O(N__51277),
            .I(N__51249));
    Span4Mux_h I__11681 (
            .O(N__51274),
            .I(N__51243));
    Span4Mux_h I__11680 (
            .O(N__51271),
            .I(N__51243));
    InMux I__11679 (
            .O(N__51270),
            .I(N__51236));
    InMux I__11678 (
            .O(N__51267),
            .I(N__51236));
    InMux I__11677 (
            .O(N__51266),
            .I(N__51236));
    LocalMux I__11676 (
            .O(N__51261),
            .I(N__51227));
    LocalMux I__11675 (
            .O(N__51258),
            .I(N__51227));
    LocalMux I__11674 (
            .O(N__51255),
            .I(N__51227));
    Span4Mux_h I__11673 (
            .O(N__51252),
            .I(N__51227));
    InMux I__11672 (
            .O(N__51249),
            .I(N__51222));
    InMux I__11671 (
            .O(N__51248),
            .I(N__51222));
    Odrv4 I__11670 (
            .O(N__51243),
            .I(n1356));
    LocalMux I__11669 (
            .O(N__51236),
            .I(n1356));
    Odrv4 I__11668 (
            .O(N__51227),
            .I(n1356));
    LocalMux I__11667 (
            .O(N__51222),
            .I(n1356));
    CascadeMux I__11666 (
            .O(N__51213),
            .I(N__51208));
    InMux I__11665 (
            .O(N__51212),
            .I(N__51205));
    InMux I__11664 (
            .O(N__51211),
            .I(N__51202));
    InMux I__11663 (
            .O(N__51208),
            .I(N__51199));
    LocalMux I__11662 (
            .O(N__51205),
            .I(N__51194));
    LocalMux I__11661 (
            .O(N__51202),
            .I(N__51194));
    LocalMux I__11660 (
            .O(N__51199),
            .I(n1424));
    Odrv4 I__11659 (
            .O(N__51194),
            .I(n1424));
    InMux I__11658 (
            .O(N__51189),
            .I(N__51186));
    LocalMux I__11657 (
            .O(N__51186),
            .I(N__51183));
    Odrv4 I__11656 (
            .O(N__51183),
            .I(n1294));
    CascadeMux I__11655 (
            .O(N__51180),
            .I(N__51177));
    InMux I__11654 (
            .O(N__51177),
            .I(N__51174));
    LocalMux I__11653 (
            .O(N__51174),
            .I(N__51171));
    Odrv4 I__11652 (
            .O(N__51171),
            .I(n1295));
    InMux I__11651 (
            .O(N__51168),
            .I(N__51161));
    InMux I__11650 (
            .O(N__51167),
            .I(N__51161));
    InMux I__11649 (
            .O(N__51166),
            .I(N__51158));
    LocalMux I__11648 (
            .O(N__51161),
            .I(n1227));
    LocalMux I__11647 (
            .O(N__51158),
            .I(n1227));
    CascadeMux I__11646 (
            .O(N__51153),
            .I(n14482_cascade_));
    InMux I__11645 (
            .O(N__51150),
            .I(N__51147));
    LocalMux I__11644 (
            .O(N__51147),
            .I(N__51144));
    Odrv4 I__11643 (
            .O(N__51144),
            .I(n1296));
    CascadeMux I__11642 (
            .O(N__51141),
            .I(n1257_cascade_));
    InMux I__11641 (
            .O(N__51138),
            .I(N__51134));
    CascadeMux I__11640 (
            .O(N__51137),
            .I(N__51131));
    LocalMux I__11639 (
            .O(N__51134),
            .I(N__51128));
    InMux I__11638 (
            .O(N__51131),
            .I(N__51125));
    Odrv4 I__11637 (
            .O(N__51128),
            .I(n1328));
    LocalMux I__11636 (
            .O(N__51125),
            .I(n1328));
    InMux I__11635 (
            .O(N__51120),
            .I(N__51115));
    InMux I__11634 (
            .O(N__51119),
            .I(N__51112));
    InMux I__11633 (
            .O(N__51118),
            .I(N__51109));
    LocalMux I__11632 (
            .O(N__51115),
            .I(n1327));
    LocalMux I__11631 (
            .O(N__51112),
            .I(n1327));
    LocalMux I__11630 (
            .O(N__51109),
            .I(n1327));
    CascadeMux I__11629 (
            .O(N__51102),
            .I(n1328_cascade_));
    CascadeMux I__11628 (
            .O(N__51099),
            .I(N__51095));
    CascadeMux I__11627 (
            .O(N__51098),
            .I(N__51092));
    InMux I__11626 (
            .O(N__51095),
            .I(N__51088));
    InMux I__11625 (
            .O(N__51092),
            .I(N__51085));
    InMux I__11624 (
            .O(N__51091),
            .I(N__51082));
    LocalMux I__11623 (
            .O(N__51088),
            .I(n1326));
    LocalMux I__11622 (
            .O(N__51085),
            .I(n1326));
    LocalMux I__11621 (
            .O(N__51082),
            .I(n1326));
    InMux I__11620 (
            .O(N__51075),
            .I(N__51072));
    LocalMux I__11619 (
            .O(N__51072),
            .I(N__51069));
    Span4Mux_h I__11618 (
            .O(N__51069),
            .I(N__51066));
    Odrv4 I__11617 (
            .O(N__51066),
            .I(n14282));
    CascadeMux I__11616 (
            .O(N__51063),
            .I(N__51060));
    InMux I__11615 (
            .O(N__51060),
            .I(N__51057));
    LocalMux I__11614 (
            .O(N__51057),
            .I(N__51052));
    InMux I__11613 (
            .O(N__51056),
            .I(N__51049));
    InMux I__11612 (
            .O(N__51055),
            .I(N__51046));
    Span4Mux_h I__11611 (
            .O(N__51052),
            .I(N__51043));
    LocalMux I__11610 (
            .O(N__51049),
            .I(n1429));
    LocalMux I__11609 (
            .O(N__51046),
            .I(n1429));
    Odrv4 I__11608 (
            .O(N__51043),
            .I(n1429));
    InMux I__11607 (
            .O(N__51036),
            .I(N__51033));
    LocalMux I__11606 (
            .O(N__51033),
            .I(N__51030));
    Odrv4 I__11605 (
            .O(N__51030),
            .I(n1496));
    InMux I__11604 (
            .O(N__51027),
            .I(n12542));
    CascadeMux I__11603 (
            .O(N__51024),
            .I(N__51021));
    InMux I__11602 (
            .O(N__51021),
            .I(N__51017));
    CascadeMux I__11601 (
            .O(N__51020),
            .I(N__51013));
    LocalMux I__11600 (
            .O(N__51017),
            .I(N__51010));
    InMux I__11599 (
            .O(N__51016),
            .I(N__51007));
    InMux I__11598 (
            .O(N__51013),
            .I(N__51004));
    Span4Mux_v I__11597 (
            .O(N__51010),
            .I(N__51001));
    LocalMux I__11596 (
            .O(N__51007),
            .I(n1428));
    LocalMux I__11595 (
            .O(N__51004),
            .I(n1428));
    Odrv4 I__11594 (
            .O(N__51001),
            .I(n1428));
    InMux I__11593 (
            .O(N__50994),
            .I(N__50991));
    LocalMux I__11592 (
            .O(N__50991),
            .I(N__50988));
    Span4Mux_h I__11591 (
            .O(N__50988),
            .I(N__50985));
    Odrv4 I__11590 (
            .O(N__50985),
            .I(n1495));
    InMux I__11589 (
            .O(N__50982),
            .I(n12543));
    CascadeMux I__11588 (
            .O(N__50979),
            .I(N__50975));
    InMux I__11587 (
            .O(N__50978),
            .I(N__50972));
    InMux I__11586 (
            .O(N__50975),
            .I(N__50969));
    LocalMux I__11585 (
            .O(N__50972),
            .I(N__50966));
    LocalMux I__11584 (
            .O(N__50969),
            .I(n1427));
    Odrv4 I__11583 (
            .O(N__50966),
            .I(n1427));
    InMux I__11582 (
            .O(N__50961),
            .I(N__50958));
    LocalMux I__11581 (
            .O(N__50958),
            .I(n1494));
    InMux I__11580 (
            .O(N__50955),
            .I(n12544));
    CascadeMux I__11579 (
            .O(N__50952),
            .I(N__50949));
    InMux I__11578 (
            .O(N__50949),
            .I(N__50944));
    InMux I__11577 (
            .O(N__50948),
            .I(N__50939));
    InMux I__11576 (
            .O(N__50947),
            .I(N__50939));
    LocalMux I__11575 (
            .O(N__50944),
            .I(n1426));
    LocalMux I__11574 (
            .O(N__50939),
            .I(n1426));
    InMux I__11573 (
            .O(N__50934),
            .I(N__50931));
    LocalMux I__11572 (
            .O(N__50931),
            .I(n1493));
    InMux I__11571 (
            .O(N__50928),
            .I(bfn_16_20_0_));
    CascadeMux I__11570 (
            .O(N__50925),
            .I(N__50922));
    InMux I__11569 (
            .O(N__50922),
            .I(N__50917));
    InMux I__11568 (
            .O(N__50921),
            .I(N__50912));
    InMux I__11567 (
            .O(N__50920),
            .I(N__50912));
    LocalMux I__11566 (
            .O(N__50917),
            .I(n1425));
    LocalMux I__11565 (
            .O(N__50912),
            .I(n1425));
    CascadeMux I__11564 (
            .O(N__50907),
            .I(N__50904));
    InMux I__11563 (
            .O(N__50904),
            .I(N__50901));
    LocalMux I__11562 (
            .O(N__50901),
            .I(n1492));
    InMux I__11561 (
            .O(N__50898),
            .I(n12546));
    InMux I__11560 (
            .O(N__50895),
            .I(N__50892));
    LocalMux I__11559 (
            .O(N__50892),
            .I(n1491));
    InMux I__11558 (
            .O(N__50889),
            .I(n12547));
    CascadeMux I__11557 (
            .O(N__50886),
            .I(N__50883));
    InMux I__11556 (
            .O(N__50883),
            .I(N__50880));
    LocalMux I__11555 (
            .O(N__50880),
            .I(N__50876));
    InMux I__11554 (
            .O(N__50879),
            .I(N__50872));
    Span4Mux_h I__11553 (
            .O(N__50876),
            .I(N__50869));
    InMux I__11552 (
            .O(N__50875),
            .I(N__50866));
    LocalMux I__11551 (
            .O(N__50872),
            .I(n1423));
    Odrv4 I__11550 (
            .O(N__50869),
            .I(n1423));
    LocalMux I__11549 (
            .O(N__50866),
            .I(n1423));
    CascadeMux I__11548 (
            .O(N__50859),
            .I(N__50856));
    InMux I__11547 (
            .O(N__50856),
            .I(N__50853));
    LocalMux I__11546 (
            .O(N__50853),
            .I(N__50850));
    Odrv4 I__11545 (
            .O(N__50850),
            .I(n1490));
    InMux I__11544 (
            .O(N__50847),
            .I(n12548));
    CascadeMux I__11543 (
            .O(N__50844),
            .I(N__50841));
    InMux I__11542 (
            .O(N__50841),
            .I(N__50837));
    InMux I__11541 (
            .O(N__50840),
            .I(N__50834));
    LocalMux I__11540 (
            .O(N__50837),
            .I(N__50831));
    LocalMux I__11539 (
            .O(N__50834),
            .I(N__50828));
    Odrv4 I__11538 (
            .O(N__50831),
            .I(n1422));
    Odrv4 I__11537 (
            .O(N__50828),
            .I(n1422));
    InMux I__11536 (
            .O(N__50823),
            .I(n12549));
    CascadeMux I__11535 (
            .O(N__50820),
            .I(N__50817));
    InMux I__11534 (
            .O(N__50817),
            .I(N__50814));
    LocalMux I__11533 (
            .O(N__50814),
            .I(N__50810));
    InMux I__11532 (
            .O(N__50813),
            .I(N__50807));
    Odrv4 I__11531 (
            .O(N__50810),
            .I(n1521));
    LocalMux I__11530 (
            .O(N__50807),
            .I(n1521));
    InMux I__11529 (
            .O(N__50802),
            .I(N__50799));
    LocalMux I__11528 (
            .O(N__50799),
            .I(N__50795));
    CascadeMux I__11527 (
            .O(N__50798),
            .I(N__50792));
    Span4Mux_h I__11526 (
            .O(N__50795),
            .I(N__50789));
    InMux I__11525 (
            .O(N__50792),
            .I(N__50786));
    Odrv4 I__11524 (
            .O(N__50789),
            .I(n1527));
    LocalMux I__11523 (
            .O(N__50786),
            .I(n1527));
    InMux I__11522 (
            .O(N__50781),
            .I(N__50778));
    LocalMux I__11521 (
            .O(N__50778),
            .I(N__50775));
    Span4Mux_h I__11520 (
            .O(N__50775),
            .I(N__50772));
    Odrv4 I__11519 (
            .O(N__50772),
            .I(n1594));
    CascadeMux I__11518 (
            .O(N__50769),
            .I(N__50766));
    InMux I__11517 (
            .O(N__50766),
            .I(N__50761));
    InMux I__11516 (
            .O(N__50765),
            .I(N__50756));
    InMux I__11515 (
            .O(N__50764),
            .I(N__50756));
    LocalMux I__11514 (
            .O(N__50761),
            .I(n1626_adj_613));
    LocalMux I__11513 (
            .O(N__50756),
            .I(n1626_adj_613));
    CascadeMux I__11512 (
            .O(N__50751),
            .I(N__50748));
    InMux I__11511 (
            .O(N__50748),
            .I(N__50743));
    InMux I__11510 (
            .O(N__50747),
            .I(N__50740));
    InMux I__11509 (
            .O(N__50746),
            .I(N__50737));
    LocalMux I__11508 (
            .O(N__50743),
            .I(N__50734));
    LocalMux I__11507 (
            .O(N__50740),
            .I(n1529));
    LocalMux I__11506 (
            .O(N__50737),
            .I(n1529));
    Odrv4 I__11505 (
            .O(N__50734),
            .I(n1529));
    CascadeMux I__11504 (
            .O(N__50727),
            .I(N__50724));
    InMux I__11503 (
            .O(N__50724),
            .I(N__50721));
    LocalMux I__11502 (
            .O(N__50721),
            .I(N__50718));
    Span4Mux_h I__11501 (
            .O(N__50718),
            .I(N__50715));
    Odrv4 I__11500 (
            .O(N__50715),
            .I(n1596));
    CascadeMux I__11499 (
            .O(N__50712),
            .I(N__50708));
    CascadeMux I__11498 (
            .O(N__50711),
            .I(N__50705));
    InMux I__11497 (
            .O(N__50708),
            .I(N__50701));
    InMux I__11496 (
            .O(N__50705),
            .I(N__50698));
    InMux I__11495 (
            .O(N__50704),
            .I(N__50695));
    LocalMux I__11494 (
            .O(N__50701),
            .I(n1628_adj_615));
    LocalMux I__11493 (
            .O(N__50698),
            .I(n1628_adj_615));
    LocalMux I__11492 (
            .O(N__50695),
            .I(n1628_adj_615));
    InMux I__11491 (
            .O(N__50688),
            .I(N__50685));
    LocalMux I__11490 (
            .O(N__50685),
            .I(N__50682));
    Span4Mux_h I__11489 (
            .O(N__50682),
            .I(N__50679));
    Odrv4 I__11488 (
            .O(N__50679),
            .I(n1597));
    InMux I__11487 (
            .O(N__50676),
            .I(N__50673));
    LocalMux I__11486 (
            .O(N__50673),
            .I(N__50669));
    InMux I__11485 (
            .O(N__50672),
            .I(N__50663));
    Sp12to4 I__11484 (
            .O(N__50669),
            .I(N__50658));
    InMux I__11483 (
            .O(N__50668),
            .I(N__50655));
    CascadeMux I__11482 (
            .O(N__50667),
            .I(N__50649));
    CascadeMux I__11481 (
            .O(N__50666),
            .I(N__50643));
    LocalMux I__11480 (
            .O(N__50663),
            .I(N__50640));
    CascadeMux I__11479 (
            .O(N__50662),
            .I(N__50637));
    CascadeMux I__11478 (
            .O(N__50661),
            .I(N__50634));
    Span12Mux_v I__11477 (
            .O(N__50658),
            .I(N__50629));
    LocalMux I__11476 (
            .O(N__50655),
            .I(N__50626));
    InMux I__11475 (
            .O(N__50654),
            .I(N__50623));
    InMux I__11474 (
            .O(N__50653),
            .I(N__50618));
    InMux I__11473 (
            .O(N__50652),
            .I(N__50618));
    InMux I__11472 (
            .O(N__50649),
            .I(N__50607));
    InMux I__11471 (
            .O(N__50648),
            .I(N__50607));
    InMux I__11470 (
            .O(N__50647),
            .I(N__50607));
    InMux I__11469 (
            .O(N__50646),
            .I(N__50607));
    InMux I__11468 (
            .O(N__50643),
            .I(N__50607));
    Span4Mux_h I__11467 (
            .O(N__50640),
            .I(N__50604));
    InMux I__11466 (
            .O(N__50637),
            .I(N__50595));
    InMux I__11465 (
            .O(N__50634),
            .I(N__50595));
    InMux I__11464 (
            .O(N__50633),
            .I(N__50595));
    InMux I__11463 (
            .O(N__50632),
            .I(N__50595));
    Odrv12 I__11462 (
            .O(N__50629),
            .I(n1554));
    Odrv4 I__11461 (
            .O(N__50626),
            .I(n1554));
    LocalMux I__11460 (
            .O(N__50623),
            .I(n1554));
    LocalMux I__11459 (
            .O(N__50618),
            .I(n1554));
    LocalMux I__11458 (
            .O(N__50607),
            .I(n1554));
    Odrv4 I__11457 (
            .O(N__50604),
            .I(n1554));
    LocalMux I__11456 (
            .O(N__50595),
            .I(n1554));
    CascadeMux I__11455 (
            .O(N__50580),
            .I(N__50577));
    InMux I__11454 (
            .O(N__50577),
            .I(N__50572));
    InMux I__11453 (
            .O(N__50576),
            .I(N__50569));
    InMux I__11452 (
            .O(N__50575),
            .I(N__50566));
    LocalMux I__11451 (
            .O(N__50572),
            .I(N__50563));
    LocalMux I__11450 (
            .O(N__50569),
            .I(n1530));
    LocalMux I__11449 (
            .O(N__50566),
            .I(n1530));
    Odrv4 I__11448 (
            .O(N__50563),
            .I(n1530));
    CascadeMux I__11447 (
            .O(N__50556),
            .I(N__50551));
    CascadeMux I__11446 (
            .O(N__50555),
            .I(N__50548));
    InMux I__11445 (
            .O(N__50554),
            .I(N__50545));
    InMux I__11444 (
            .O(N__50551),
            .I(N__50542));
    InMux I__11443 (
            .O(N__50548),
            .I(N__50539));
    LocalMux I__11442 (
            .O(N__50545),
            .I(N__50536));
    LocalMux I__11441 (
            .O(N__50542),
            .I(n1629_adj_616));
    LocalMux I__11440 (
            .O(N__50539),
            .I(n1629_adj_616));
    Odrv4 I__11439 (
            .O(N__50536),
            .I(n1629_adj_616));
    InMux I__11438 (
            .O(N__50529),
            .I(N__50525));
    InMux I__11437 (
            .O(N__50528),
            .I(N__50522));
    LocalMux I__11436 (
            .O(N__50525),
            .I(N__50516));
    LocalMux I__11435 (
            .O(N__50522),
            .I(N__50516));
    InMux I__11434 (
            .O(N__50521),
            .I(N__50513));
    Span4Mux_h I__11433 (
            .O(N__50516),
            .I(N__50510));
    LocalMux I__11432 (
            .O(N__50513),
            .I(N__50507));
    Odrv4 I__11431 (
            .O(N__50510),
            .I(n300));
    Odrv4 I__11430 (
            .O(N__50507),
            .I(n300));
    InMux I__11429 (
            .O(N__50502),
            .I(N__50499));
    LocalMux I__11428 (
            .O(N__50499),
            .I(N__50496));
    Odrv12 I__11427 (
            .O(N__50496),
            .I(n1501));
    InMux I__11426 (
            .O(N__50493),
            .I(bfn_16_19_0_));
    CascadeMux I__11425 (
            .O(N__50490),
            .I(N__50486));
    CascadeMux I__11424 (
            .O(N__50489),
            .I(N__50483));
    InMux I__11423 (
            .O(N__50486),
            .I(N__50480));
    InMux I__11422 (
            .O(N__50483),
            .I(N__50477));
    LocalMux I__11421 (
            .O(N__50480),
            .I(N__50472));
    LocalMux I__11420 (
            .O(N__50477),
            .I(N__50472));
    Span4Mux_h I__11419 (
            .O(N__50472),
            .I(N__50469));
    Odrv4 I__11418 (
            .O(N__50469),
            .I(n1433));
    InMux I__11417 (
            .O(N__50466),
            .I(N__50463));
    LocalMux I__11416 (
            .O(N__50463),
            .I(n1500));
    InMux I__11415 (
            .O(N__50460),
            .I(n12538));
    CascadeMux I__11414 (
            .O(N__50457),
            .I(N__50454));
    InMux I__11413 (
            .O(N__50454),
            .I(N__50450));
    InMux I__11412 (
            .O(N__50453),
            .I(N__50447));
    LocalMux I__11411 (
            .O(N__50450),
            .I(N__50444));
    LocalMux I__11410 (
            .O(N__50447),
            .I(N__50440));
    Span4Mux_v I__11409 (
            .O(N__50444),
            .I(N__50437));
    InMux I__11408 (
            .O(N__50443),
            .I(N__50434));
    Odrv4 I__11407 (
            .O(N__50440),
            .I(n1432));
    Odrv4 I__11406 (
            .O(N__50437),
            .I(n1432));
    LocalMux I__11405 (
            .O(N__50434),
            .I(n1432));
    InMux I__11404 (
            .O(N__50427),
            .I(N__50424));
    LocalMux I__11403 (
            .O(N__50424),
            .I(N__50421));
    Odrv4 I__11402 (
            .O(N__50421),
            .I(n1499));
    InMux I__11401 (
            .O(N__50418),
            .I(n12539));
    CascadeMux I__11400 (
            .O(N__50415),
            .I(N__50411));
    InMux I__11399 (
            .O(N__50414),
            .I(N__50407));
    InMux I__11398 (
            .O(N__50411),
            .I(N__50404));
    InMux I__11397 (
            .O(N__50410),
            .I(N__50401));
    LocalMux I__11396 (
            .O(N__50407),
            .I(n1431));
    LocalMux I__11395 (
            .O(N__50404),
            .I(n1431));
    LocalMux I__11394 (
            .O(N__50401),
            .I(n1431));
    InMux I__11393 (
            .O(N__50394),
            .I(N__50391));
    LocalMux I__11392 (
            .O(N__50391),
            .I(n1498));
    InMux I__11391 (
            .O(N__50388),
            .I(n12540));
    CascadeMux I__11390 (
            .O(N__50385),
            .I(N__50381));
    CascadeMux I__11389 (
            .O(N__50384),
            .I(N__50378));
    InMux I__11388 (
            .O(N__50381),
            .I(N__50375));
    InMux I__11387 (
            .O(N__50378),
            .I(N__50372));
    LocalMux I__11386 (
            .O(N__50375),
            .I(N__50366));
    LocalMux I__11385 (
            .O(N__50372),
            .I(N__50366));
    InMux I__11384 (
            .O(N__50371),
            .I(N__50363));
    Span4Mux_h I__11383 (
            .O(N__50366),
            .I(N__50360));
    LocalMux I__11382 (
            .O(N__50363),
            .I(n1430));
    Odrv4 I__11381 (
            .O(N__50360),
            .I(n1430));
    InMux I__11380 (
            .O(N__50355),
            .I(N__50352));
    LocalMux I__11379 (
            .O(N__50352),
            .I(n1497));
    InMux I__11378 (
            .O(N__50349),
            .I(n12541));
    CascadeMux I__11377 (
            .O(N__50346),
            .I(n1727_cascade_));
    InMux I__11376 (
            .O(N__50343),
            .I(N__50340));
    LocalMux I__11375 (
            .O(N__50340),
            .I(N__50335));
    CascadeMux I__11374 (
            .O(N__50339),
            .I(N__50332));
    InMux I__11373 (
            .O(N__50338),
            .I(N__50329));
    Span4Mux_h I__11372 (
            .O(N__50335),
            .I(N__50326));
    InMux I__11371 (
            .O(N__50332),
            .I(N__50323));
    LocalMux I__11370 (
            .O(N__50329),
            .I(N__50320));
    Odrv4 I__11369 (
            .O(N__50326),
            .I(n1726));
    LocalMux I__11368 (
            .O(N__50323),
            .I(n1726));
    Odrv4 I__11367 (
            .O(N__50320),
            .I(n1726));
    InMux I__11366 (
            .O(N__50313),
            .I(N__50309));
    CascadeMux I__11365 (
            .O(N__50312),
            .I(N__50306));
    LocalMux I__11364 (
            .O(N__50309),
            .I(N__50303));
    InMux I__11363 (
            .O(N__50306),
            .I(N__50300));
    Span4Mux_h I__11362 (
            .O(N__50303),
            .I(N__50294));
    LocalMux I__11361 (
            .O(N__50300),
            .I(N__50294));
    InMux I__11360 (
            .O(N__50299),
            .I(N__50291));
    Odrv4 I__11359 (
            .O(N__50294),
            .I(n1724));
    LocalMux I__11358 (
            .O(N__50291),
            .I(n1724));
    InMux I__11357 (
            .O(N__50286),
            .I(N__50282));
    CascadeMux I__11356 (
            .O(N__50285),
            .I(N__50279));
    LocalMux I__11355 (
            .O(N__50282),
            .I(N__50276));
    InMux I__11354 (
            .O(N__50279),
            .I(N__50273));
    Span4Mux_h I__11353 (
            .O(N__50276),
            .I(N__50268));
    LocalMux I__11352 (
            .O(N__50273),
            .I(N__50268));
    Span4Mux_h I__11351 (
            .O(N__50268),
            .I(N__50264));
    InMux I__11350 (
            .O(N__50267),
            .I(N__50261));
    Odrv4 I__11349 (
            .O(N__50264),
            .I(n1725));
    LocalMux I__11348 (
            .O(N__50261),
            .I(n1725));
    CascadeMux I__11347 (
            .O(N__50256),
            .I(n14166_cascade_));
    InMux I__11346 (
            .O(N__50253),
            .I(N__50250));
    LocalMux I__11345 (
            .O(N__50250),
            .I(N__50245));
    CascadeMux I__11344 (
            .O(N__50249),
            .I(N__50242));
    InMux I__11343 (
            .O(N__50248),
            .I(N__50239));
    Span4Mux_h I__11342 (
            .O(N__50245),
            .I(N__50236));
    InMux I__11341 (
            .O(N__50242),
            .I(N__50233));
    LocalMux I__11340 (
            .O(N__50239),
            .I(N__50230));
    Odrv4 I__11339 (
            .O(N__50236),
            .I(n1723));
    LocalMux I__11338 (
            .O(N__50233),
            .I(n1723));
    Odrv4 I__11337 (
            .O(N__50230),
            .I(n1723));
    InMux I__11336 (
            .O(N__50223),
            .I(N__50220));
    LocalMux I__11335 (
            .O(N__50220),
            .I(N__50217));
    Span4Mux_v I__11334 (
            .O(N__50217),
            .I(N__50214));
    Span4Mux_h I__11333 (
            .O(N__50214),
            .I(N__50211));
    Odrv4 I__11332 (
            .O(N__50211),
            .I(n14172));
    InMux I__11331 (
            .O(N__50208),
            .I(N__50205));
    LocalMux I__11330 (
            .O(N__50205),
            .I(n1696));
    InMux I__11329 (
            .O(N__50202),
            .I(N__50199));
    LocalMux I__11328 (
            .O(N__50199),
            .I(N__50196));
    Span4Mux_h I__11327 (
            .O(N__50196),
            .I(N__50192));
    CascadeMux I__11326 (
            .O(N__50195),
            .I(N__50189));
    Span4Mux_h I__11325 (
            .O(N__50192),
            .I(N__50183));
    InMux I__11324 (
            .O(N__50189),
            .I(N__50176));
    InMux I__11323 (
            .O(N__50188),
            .I(N__50176));
    InMux I__11322 (
            .O(N__50187),
            .I(N__50176));
    CascadeMux I__11321 (
            .O(N__50186),
            .I(N__50172));
    Span4Mux_v I__11320 (
            .O(N__50183),
            .I(N__50160));
    LocalMux I__11319 (
            .O(N__50176),
            .I(N__50160));
    InMux I__11318 (
            .O(N__50175),
            .I(N__50153));
    InMux I__11317 (
            .O(N__50172),
            .I(N__50153));
    InMux I__11316 (
            .O(N__50171),
            .I(N__50153));
    CascadeMux I__11315 (
            .O(N__50170),
            .I(N__50150));
    CascadeMux I__11314 (
            .O(N__50169),
            .I(N__50147));
    InMux I__11313 (
            .O(N__50168),
            .I(N__50137));
    InMux I__11312 (
            .O(N__50167),
            .I(N__50137));
    InMux I__11311 (
            .O(N__50166),
            .I(N__50137));
    InMux I__11310 (
            .O(N__50165),
            .I(N__50134));
    Span4Mux_v I__11309 (
            .O(N__50160),
            .I(N__50129));
    LocalMux I__11308 (
            .O(N__50153),
            .I(N__50129));
    InMux I__11307 (
            .O(N__50150),
            .I(N__50118));
    InMux I__11306 (
            .O(N__50147),
            .I(N__50118));
    InMux I__11305 (
            .O(N__50146),
            .I(N__50118));
    InMux I__11304 (
            .O(N__50145),
            .I(N__50118));
    InMux I__11303 (
            .O(N__50144),
            .I(N__50118));
    LocalMux I__11302 (
            .O(N__50137),
            .I(n1653));
    LocalMux I__11301 (
            .O(N__50134),
            .I(n1653));
    Odrv4 I__11300 (
            .O(N__50129),
            .I(n1653));
    LocalMux I__11299 (
            .O(N__50118),
            .I(n1653));
    CascadeMux I__11298 (
            .O(N__50109),
            .I(N__50106));
    InMux I__11297 (
            .O(N__50106),
            .I(N__50102));
    CascadeMux I__11296 (
            .O(N__50105),
            .I(N__50099));
    LocalMux I__11295 (
            .O(N__50102),
            .I(N__50096));
    InMux I__11294 (
            .O(N__50099),
            .I(N__50093));
    Span4Mux_v I__11293 (
            .O(N__50096),
            .I(N__50087));
    LocalMux I__11292 (
            .O(N__50093),
            .I(N__50087));
    InMux I__11291 (
            .O(N__50092),
            .I(N__50084));
    Odrv4 I__11290 (
            .O(N__50087),
            .I(n1728));
    LocalMux I__11289 (
            .O(N__50084),
            .I(n1728));
    InMux I__11288 (
            .O(N__50079),
            .I(N__50076));
    LocalMux I__11287 (
            .O(N__50076),
            .I(N__50073));
    Odrv4 I__11286 (
            .O(N__50073),
            .I(n14508));
    CascadeMux I__11285 (
            .O(N__50070),
            .I(N__50067));
    InMux I__11284 (
            .O(N__50067),
            .I(N__50064));
    LocalMux I__11283 (
            .O(N__50064),
            .I(N__50061));
    Span4Mux_h I__11282 (
            .O(N__50061),
            .I(N__50058));
    Odrv4 I__11281 (
            .O(N__50058),
            .I(n1395));
    CascadeMux I__11280 (
            .O(N__50055),
            .I(n1427_cascade_));
    CascadeMux I__11279 (
            .O(N__50052),
            .I(N__50048));
    CascadeMux I__11278 (
            .O(N__50051),
            .I(N__50045));
    InMux I__11277 (
            .O(N__50048),
            .I(N__50042));
    InMux I__11276 (
            .O(N__50045),
            .I(N__50039));
    LocalMux I__11275 (
            .O(N__50042),
            .I(N__50034));
    LocalMux I__11274 (
            .O(N__50039),
            .I(N__50034));
    Span4Mux_h I__11273 (
            .O(N__50034),
            .I(N__50031));
    Odrv4 I__11272 (
            .O(N__50031),
            .I(n1526));
    CascadeMux I__11271 (
            .O(N__50028),
            .I(n1526_cascade_));
    InMux I__11270 (
            .O(N__50025),
            .I(N__50022));
    LocalMux I__11269 (
            .O(N__50022),
            .I(N__50019));
    Span4Mux_h I__11268 (
            .O(N__50019),
            .I(N__50016));
    Odrv4 I__11267 (
            .O(N__50016),
            .I(n1593));
    CascadeMux I__11266 (
            .O(N__50013),
            .I(N__50009));
    CascadeMux I__11265 (
            .O(N__50012),
            .I(N__50006));
    InMux I__11264 (
            .O(N__50009),
            .I(N__50000));
    InMux I__11263 (
            .O(N__50006),
            .I(N__50000));
    InMux I__11262 (
            .O(N__50005),
            .I(N__49997));
    LocalMux I__11261 (
            .O(N__50000),
            .I(n1625_adj_612));
    LocalMux I__11260 (
            .O(N__49997),
            .I(n1625_adj_612));
    InMux I__11259 (
            .O(N__49992),
            .I(N__49988));
    InMux I__11258 (
            .O(N__49991),
            .I(N__49984));
    LocalMux I__11257 (
            .O(N__49988),
            .I(N__49981));
    CascadeMux I__11256 (
            .O(N__49987),
            .I(N__49978));
    LocalMux I__11255 (
            .O(N__49984),
            .I(N__49974));
    Span4Mux_v I__11254 (
            .O(N__49981),
            .I(N__49971));
    InMux I__11253 (
            .O(N__49978),
            .I(N__49968));
    InMux I__11252 (
            .O(N__49977),
            .I(N__49965));
    Odrv4 I__11251 (
            .O(N__49974),
            .I(n1528));
    Odrv4 I__11250 (
            .O(N__49971),
            .I(n1528));
    LocalMux I__11249 (
            .O(N__49968),
            .I(n1528));
    LocalMux I__11248 (
            .O(N__49965),
            .I(n1528));
    CascadeMux I__11247 (
            .O(N__49956),
            .I(N__49952));
    CascadeMux I__11246 (
            .O(N__49955),
            .I(N__49949));
    InMux I__11245 (
            .O(N__49952),
            .I(N__49946));
    InMux I__11244 (
            .O(N__49949),
            .I(N__49943));
    LocalMux I__11243 (
            .O(N__49946),
            .I(N__49940));
    LocalMux I__11242 (
            .O(N__49943),
            .I(N__49937));
    Span4Mux_h I__11241 (
            .O(N__49940),
            .I(N__49934));
    Odrv4 I__11240 (
            .O(N__49937),
            .I(n1595));
    Odrv4 I__11239 (
            .O(N__49934),
            .I(n1595));
    CascadeMux I__11238 (
            .O(N__49929),
            .I(N__49925));
    InMux I__11237 (
            .O(N__49928),
            .I(N__49922));
    InMux I__11236 (
            .O(N__49925),
            .I(N__49919));
    LocalMux I__11235 (
            .O(N__49922),
            .I(n1627_adj_614));
    LocalMux I__11234 (
            .O(N__49919),
            .I(n1627_adj_614));
    InMux I__11233 (
            .O(N__49914),
            .I(n12966));
    CascadeMux I__11232 (
            .O(N__49911),
            .I(N__49904));
    CascadeMux I__11231 (
            .O(N__49910),
            .I(N__49900));
    CascadeMux I__11230 (
            .O(N__49909),
            .I(N__49896));
    InMux I__11229 (
            .O(N__49908),
            .I(N__49881));
    InMux I__11228 (
            .O(N__49907),
            .I(N__49881));
    InMux I__11227 (
            .O(N__49904),
            .I(N__49881));
    InMux I__11226 (
            .O(N__49903),
            .I(N__49881));
    InMux I__11225 (
            .O(N__49900),
            .I(N__49881));
    InMux I__11224 (
            .O(N__49899),
            .I(N__49881));
    InMux I__11223 (
            .O(N__49896),
            .I(N__49881));
    LocalMux I__11222 (
            .O(N__49881),
            .I(n11514));
    InMux I__11221 (
            .O(N__49878),
            .I(N__49875));
    LocalMux I__11220 (
            .O(N__49875),
            .I(n15089));
    InMux I__11219 (
            .O(N__49872),
            .I(n12967));
    CascadeMux I__11218 (
            .O(N__49869),
            .I(N__49866));
    InMux I__11217 (
            .O(N__49866),
            .I(N__49863));
    LocalMux I__11216 (
            .O(N__49863),
            .I(N__49858));
    InMux I__11215 (
            .O(N__49862),
            .I(N__49853));
    InMux I__11214 (
            .O(N__49861),
            .I(N__49853));
    Odrv4 I__11213 (
            .O(N__49858),
            .I(dti_counter_7));
    LocalMux I__11212 (
            .O(N__49853),
            .I(dti_counter_7));
    CascadeMux I__11211 (
            .O(N__49848),
            .I(n4_adj_716_cascade_));
    CascadeMux I__11210 (
            .O(N__49845),
            .I(N__49842));
    InMux I__11209 (
            .O(N__49842),
            .I(N__49837));
    InMux I__11208 (
            .O(N__49841),
            .I(N__49834));
    InMux I__11207 (
            .O(N__49840),
            .I(N__49831));
    LocalMux I__11206 (
            .O(N__49837),
            .I(dti_counter_6));
    LocalMux I__11205 (
            .O(N__49834),
            .I(dti_counter_6));
    LocalMux I__11204 (
            .O(N__49831),
            .I(dti_counter_6));
    InMux I__11203 (
            .O(N__49824),
            .I(N__49821));
    LocalMux I__11202 (
            .O(N__49821),
            .I(n15090));
    InMux I__11201 (
            .O(N__49818),
            .I(N__49815));
    LocalMux I__11200 (
            .O(N__49815),
            .I(commutation_state_prev_1));
    InMux I__11199 (
            .O(N__49812),
            .I(N__49809));
    LocalMux I__11198 (
            .O(N__49809),
            .I(commutation_state_prev_2));
    InMux I__11197 (
            .O(N__49806),
            .I(N__49803));
    LocalMux I__11196 (
            .O(N__49803),
            .I(n1693_adj_621));
    InMux I__11195 (
            .O(N__49800),
            .I(N__49797));
    LocalMux I__11194 (
            .O(N__49797),
            .I(N__49794));
    Odrv4 I__11193 (
            .O(N__49794),
            .I(n1695));
    CascadeMux I__11192 (
            .O(N__49791),
            .I(N__49787));
    InMux I__11191 (
            .O(N__49790),
            .I(N__49784));
    InMux I__11190 (
            .O(N__49787),
            .I(N__49781));
    LocalMux I__11189 (
            .O(N__49784),
            .I(N__49776));
    LocalMux I__11188 (
            .O(N__49781),
            .I(N__49776));
    Odrv12 I__11187 (
            .O(N__49776),
            .I(n1727));
    InMux I__11186 (
            .O(N__49773),
            .I(N__49770));
    LocalMux I__11185 (
            .O(N__49770),
            .I(N__49767));
    Odrv4 I__11184 (
            .O(N__49767),
            .I(n15088));
    InMux I__11183 (
            .O(N__49764),
            .I(N__49759));
    InMux I__11182 (
            .O(N__49763),
            .I(N__49756));
    InMux I__11181 (
            .O(N__49762),
            .I(N__49753));
    LocalMux I__11180 (
            .O(N__49759),
            .I(dti_counter_0));
    LocalMux I__11179 (
            .O(N__49756),
            .I(dti_counter_0));
    LocalMux I__11178 (
            .O(N__49753),
            .I(dti_counter_0));
    InMux I__11177 (
            .O(N__49746),
            .I(bfn_15_31_0_));
    InMux I__11176 (
            .O(N__49743),
            .I(N__49740));
    LocalMux I__11175 (
            .O(N__49740),
            .I(n15095));
    InMux I__11174 (
            .O(N__49737),
            .I(N__49732));
    InMux I__11173 (
            .O(N__49736),
            .I(N__49729));
    InMux I__11172 (
            .O(N__49735),
            .I(N__49726));
    LocalMux I__11171 (
            .O(N__49732),
            .I(N__49723));
    LocalMux I__11170 (
            .O(N__49729),
            .I(N__49720));
    LocalMux I__11169 (
            .O(N__49726),
            .I(dti_counter_1));
    Odrv4 I__11168 (
            .O(N__49723),
            .I(dti_counter_1));
    Odrv4 I__11167 (
            .O(N__49720),
            .I(dti_counter_1));
    InMux I__11166 (
            .O(N__49713),
            .I(n12961));
    InMux I__11165 (
            .O(N__49710),
            .I(N__49707));
    LocalMux I__11164 (
            .O(N__49707),
            .I(n15094));
    CascadeMux I__11163 (
            .O(N__49704),
            .I(N__49700));
    CascadeMux I__11162 (
            .O(N__49703),
            .I(N__49696));
    InMux I__11161 (
            .O(N__49700),
            .I(N__49693));
    InMux I__11160 (
            .O(N__49699),
            .I(N__49690));
    InMux I__11159 (
            .O(N__49696),
            .I(N__49687));
    LocalMux I__11158 (
            .O(N__49693),
            .I(N__49682));
    LocalMux I__11157 (
            .O(N__49690),
            .I(N__49682));
    LocalMux I__11156 (
            .O(N__49687),
            .I(dti_counter_2));
    Odrv4 I__11155 (
            .O(N__49682),
            .I(dti_counter_2));
    InMux I__11154 (
            .O(N__49677),
            .I(n12962));
    InMux I__11153 (
            .O(N__49674),
            .I(N__49671));
    LocalMux I__11152 (
            .O(N__49671),
            .I(n15093));
    InMux I__11151 (
            .O(N__49668),
            .I(N__49663));
    InMux I__11150 (
            .O(N__49667),
            .I(N__49658));
    InMux I__11149 (
            .O(N__49666),
            .I(N__49658));
    LocalMux I__11148 (
            .O(N__49663),
            .I(dti_counter_3));
    LocalMux I__11147 (
            .O(N__49658),
            .I(dti_counter_3));
    InMux I__11146 (
            .O(N__49653),
            .I(n12963));
    InMux I__11145 (
            .O(N__49650),
            .I(N__49647));
    LocalMux I__11144 (
            .O(N__49647),
            .I(n15092));
    CascadeMux I__11143 (
            .O(N__49644),
            .I(N__49640));
    CascadeMux I__11142 (
            .O(N__49643),
            .I(N__49636));
    InMux I__11141 (
            .O(N__49640),
            .I(N__49633));
    InMux I__11140 (
            .O(N__49639),
            .I(N__49630));
    InMux I__11139 (
            .O(N__49636),
            .I(N__49627));
    LocalMux I__11138 (
            .O(N__49633),
            .I(dti_counter_4));
    LocalMux I__11137 (
            .O(N__49630),
            .I(dti_counter_4));
    LocalMux I__11136 (
            .O(N__49627),
            .I(dti_counter_4));
    InMux I__11135 (
            .O(N__49620),
            .I(n12964));
    InMux I__11134 (
            .O(N__49617),
            .I(N__49614));
    LocalMux I__11133 (
            .O(N__49614),
            .I(n15091));
    InMux I__11132 (
            .O(N__49611),
            .I(N__49606));
    InMux I__11131 (
            .O(N__49610),
            .I(N__49603));
    InMux I__11130 (
            .O(N__49609),
            .I(N__49600));
    LocalMux I__11129 (
            .O(N__49606),
            .I(dti_counter_5));
    LocalMux I__11128 (
            .O(N__49603),
            .I(dti_counter_5));
    LocalMux I__11127 (
            .O(N__49600),
            .I(dti_counter_5));
    InMux I__11126 (
            .O(N__49593),
            .I(n12965));
    InMux I__11125 (
            .O(N__49590),
            .I(N__49586));
    CascadeMux I__11124 (
            .O(N__49589),
            .I(N__49582));
    LocalMux I__11123 (
            .O(N__49586),
            .I(N__49578));
    InMux I__11122 (
            .O(N__49585),
            .I(N__49575));
    InMux I__11121 (
            .O(N__49582),
            .I(N__49572));
    InMux I__11120 (
            .O(N__49581),
            .I(N__49569));
    Span4Mux_v I__11119 (
            .O(N__49578),
            .I(N__49566));
    LocalMux I__11118 (
            .O(N__49575),
            .I(N__49561));
    LocalMux I__11117 (
            .O(N__49572),
            .I(N__49561));
    LocalMux I__11116 (
            .O(N__49569),
            .I(encoder0_position_target_20));
    Odrv4 I__11115 (
            .O(N__49566),
            .I(encoder0_position_target_20));
    Odrv4 I__11114 (
            .O(N__49561),
            .I(encoder0_position_target_20));
    InMux I__11113 (
            .O(N__49554),
            .I(n12455));
    InMux I__11112 (
            .O(N__49551),
            .I(n12456));
    CascadeMux I__11111 (
            .O(N__49548),
            .I(N__49544));
    InMux I__11110 (
            .O(N__49547),
            .I(N__49541));
    InMux I__11109 (
            .O(N__49544),
            .I(N__49538));
    LocalMux I__11108 (
            .O(N__49541),
            .I(N__49534));
    LocalMux I__11107 (
            .O(N__49538),
            .I(N__49530));
    InMux I__11106 (
            .O(N__49537),
            .I(N__49527));
    Span4Mux_h I__11105 (
            .O(N__49534),
            .I(N__49524));
    InMux I__11104 (
            .O(N__49533),
            .I(N__49521));
    Span4Mux_h I__11103 (
            .O(N__49530),
            .I(N__49516));
    LocalMux I__11102 (
            .O(N__49527),
            .I(N__49516));
    Span4Mux_h I__11101 (
            .O(N__49524),
            .I(N__49513));
    LocalMux I__11100 (
            .O(N__49521),
            .I(encoder0_position_target_22));
    Odrv4 I__11099 (
            .O(N__49516),
            .I(encoder0_position_target_22));
    Odrv4 I__11098 (
            .O(N__49513),
            .I(encoder0_position_target_22));
    InMux I__11097 (
            .O(N__49506),
            .I(n12457));
    InMux I__11096 (
            .O(N__49503),
            .I(bfn_15_28_0_));
    CascadeMux I__11095 (
            .O(N__49500),
            .I(n14_adj_718_cascade_));
    InMux I__11094 (
            .O(N__49497),
            .I(N__49494));
    LocalMux I__11093 (
            .O(N__49494),
            .I(n10_adj_719));
    CascadeMux I__11092 (
            .O(N__49491),
            .I(n5119_cascade_));
    CascadeMux I__11091 (
            .O(N__49488),
            .I(N__49485));
    InMux I__11090 (
            .O(N__49485),
            .I(N__49480));
    InMux I__11089 (
            .O(N__49484),
            .I(N__49477));
    CascadeMux I__11088 (
            .O(N__49483),
            .I(N__49474));
    LocalMux I__11087 (
            .O(N__49480),
            .I(N__49471));
    LocalMux I__11086 (
            .O(N__49477),
            .I(N__49467));
    InMux I__11085 (
            .O(N__49474),
            .I(N__49464));
    Span4Mux_v I__11084 (
            .O(N__49471),
            .I(N__49461));
    InMux I__11083 (
            .O(N__49470),
            .I(N__49458));
    Span4Mux_v I__11082 (
            .O(N__49467),
            .I(N__49455));
    LocalMux I__11081 (
            .O(N__49464),
            .I(encoder0_position_target_11));
    Odrv4 I__11080 (
            .O(N__49461),
            .I(encoder0_position_target_11));
    LocalMux I__11079 (
            .O(N__49458),
            .I(encoder0_position_target_11));
    Odrv4 I__11078 (
            .O(N__49455),
            .I(encoder0_position_target_11));
    InMux I__11077 (
            .O(N__49446),
            .I(n12446));
    CascadeMux I__11076 (
            .O(N__49443),
            .I(N__49439));
    CascadeMux I__11075 (
            .O(N__49442),
            .I(N__49436));
    InMux I__11074 (
            .O(N__49439),
            .I(N__49432));
    InMux I__11073 (
            .O(N__49436),
            .I(N__49429));
    InMux I__11072 (
            .O(N__49435),
            .I(N__49426));
    LocalMux I__11071 (
            .O(N__49432),
            .I(N__49422));
    LocalMux I__11070 (
            .O(N__49429),
            .I(N__49419));
    LocalMux I__11069 (
            .O(N__49426),
            .I(N__49416));
    InMux I__11068 (
            .O(N__49425),
            .I(N__49413));
    Span4Mux_v I__11067 (
            .O(N__49422),
            .I(N__49410));
    Span4Mux_h I__11066 (
            .O(N__49419),
            .I(N__49407));
    Span4Mux_h I__11065 (
            .O(N__49416),
            .I(N__49404));
    LocalMux I__11064 (
            .O(N__49413),
            .I(encoder0_position_target_12));
    Odrv4 I__11063 (
            .O(N__49410),
            .I(encoder0_position_target_12));
    Odrv4 I__11062 (
            .O(N__49407),
            .I(encoder0_position_target_12));
    Odrv4 I__11061 (
            .O(N__49404),
            .I(encoder0_position_target_12));
    InMux I__11060 (
            .O(N__49395),
            .I(n12447));
    CascadeMux I__11059 (
            .O(N__49392),
            .I(N__49389));
    InMux I__11058 (
            .O(N__49389),
            .I(N__49384));
    InMux I__11057 (
            .O(N__49388),
            .I(N__49381));
    CascadeMux I__11056 (
            .O(N__49387),
            .I(N__49377));
    LocalMux I__11055 (
            .O(N__49384),
            .I(N__49374));
    LocalMux I__11054 (
            .O(N__49381),
            .I(N__49371));
    InMux I__11053 (
            .O(N__49380),
            .I(N__49368));
    InMux I__11052 (
            .O(N__49377),
            .I(N__49365));
    Span4Mux_h I__11051 (
            .O(N__49374),
            .I(N__49362));
    Span4Mux_h I__11050 (
            .O(N__49371),
            .I(N__49359));
    LocalMux I__11049 (
            .O(N__49368),
            .I(N__49356));
    LocalMux I__11048 (
            .O(N__49365),
            .I(encoder0_position_target_13));
    Odrv4 I__11047 (
            .O(N__49362),
            .I(encoder0_position_target_13));
    Odrv4 I__11046 (
            .O(N__49359),
            .I(encoder0_position_target_13));
    Odrv12 I__11045 (
            .O(N__49356),
            .I(encoder0_position_target_13));
    InMux I__11044 (
            .O(N__49347),
            .I(n12448));
    CascadeMux I__11043 (
            .O(N__49344),
            .I(N__49341));
    InMux I__11042 (
            .O(N__49341),
            .I(N__49337));
    InMux I__11041 (
            .O(N__49340),
            .I(N__49334));
    LocalMux I__11040 (
            .O(N__49337),
            .I(N__49329));
    LocalMux I__11039 (
            .O(N__49334),
            .I(N__49326));
    CascadeMux I__11038 (
            .O(N__49333),
            .I(N__49323));
    InMux I__11037 (
            .O(N__49332),
            .I(N__49320));
    Span4Mux_h I__11036 (
            .O(N__49329),
            .I(N__49317));
    Span4Mux_h I__11035 (
            .O(N__49326),
            .I(N__49314));
    InMux I__11034 (
            .O(N__49323),
            .I(N__49311));
    LocalMux I__11033 (
            .O(N__49320),
            .I(encoder0_position_target_14));
    Odrv4 I__11032 (
            .O(N__49317),
            .I(encoder0_position_target_14));
    Odrv4 I__11031 (
            .O(N__49314),
            .I(encoder0_position_target_14));
    LocalMux I__11030 (
            .O(N__49311),
            .I(encoder0_position_target_14));
    InMux I__11029 (
            .O(N__49302),
            .I(n12449));
    InMux I__11028 (
            .O(N__49299),
            .I(bfn_15_27_0_));
    CascadeMux I__11027 (
            .O(N__49296),
            .I(N__49293));
    InMux I__11026 (
            .O(N__49293),
            .I(N__49290));
    LocalMux I__11025 (
            .O(N__49290),
            .I(N__49285));
    InMux I__11024 (
            .O(N__49289),
            .I(N__49282));
    InMux I__11023 (
            .O(N__49288),
            .I(N__49278));
    Span4Mux_h I__11022 (
            .O(N__49285),
            .I(N__49275));
    LocalMux I__11021 (
            .O(N__49282),
            .I(N__49272));
    InMux I__11020 (
            .O(N__49281),
            .I(N__49269));
    LocalMux I__11019 (
            .O(N__49278),
            .I(encoder0_position_target_16));
    Odrv4 I__11018 (
            .O(N__49275),
            .I(encoder0_position_target_16));
    Odrv4 I__11017 (
            .O(N__49272),
            .I(encoder0_position_target_16));
    LocalMux I__11016 (
            .O(N__49269),
            .I(encoder0_position_target_16));
    InMux I__11015 (
            .O(N__49260),
            .I(n12451));
    CascadeMux I__11014 (
            .O(N__49257),
            .I(N__49254));
    InMux I__11013 (
            .O(N__49254),
            .I(N__49250));
    CascadeMux I__11012 (
            .O(N__49253),
            .I(N__49246));
    LocalMux I__11011 (
            .O(N__49250),
            .I(N__49243));
    InMux I__11010 (
            .O(N__49249),
            .I(N__49239));
    InMux I__11009 (
            .O(N__49246),
            .I(N__49236));
    Span4Mux_h I__11008 (
            .O(N__49243),
            .I(N__49233));
    InMux I__11007 (
            .O(N__49242),
            .I(N__49230));
    LocalMux I__11006 (
            .O(N__49239),
            .I(N__49227));
    LocalMux I__11005 (
            .O(N__49236),
            .I(encoder0_position_target_17));
    Odrv4 I__11004 (
            .O(N__49233),
            .I(encoder0_position_target_17));
    LocalMux I__11003 (
            .O(N__49230),
            .I(encoder0_position_target_17));
    Odrv4 I__11002 (
            .O(N__49227),
            .I(encoder0_position_target_17));
    InMux I__11001 (
            .O(N__49218),
            .I(n12452));
    CascadeMux I__11000 (
            .O(N__49215),
            .I(N__49212));
    InMux I__10999 (
            .O(N__49212),
            .I(N__49208));
    InMux I__10998 (
            .O(N__49211),
            .I(N__49204));
    LocalMux I__10997 (
            .O(N__49208),
            .I(N__49201));
    InMux I__10996 (
            .O(N__49207),
            .I(N__49198));
    LocalMux I__10995 (
            .O(N__49204),
            .I(N__49195));
    Span4Mux_h I__10994 (
            .O(N__49201),
            .I(N__49191));
    LocalMux I__10993 (
            .O(N__49198),
            .I(N__49186));
    Span4Mux_v I__10992 (
            .O(N__49195),
            .I(N__49186));
    InMux I__10991 (
            .O(N__49194),
            .I(N__49183));
    Odrv4 I__10990 (
            .O(N__49191),
            .I(encoder0_position_target_18));
    Odrv4 I__10989 (
            .O(N__49186),
            .I(encoder0_position_target_18));
    LocalMux I__10988 (
            .O(N__49183),
            .I(encoder0_position_target_18));
    InMux I__10987 (
            .O(N__49176),
            .I(n12453));
    InMux I__10986 (
            .O(N__49173),
            .I(n12454));
    CascadeMux I__10985 (
            .O(N__49170),
            .I(N__49167));
    InMux I__10984 (
            .O(N__49167),
            .I(N__49163));
    CascadeMux I__10983 (
            .O(N__49166),
            .I(N__49160));
    LocalMux I__10982 (
            .O(N__49163),
            .I(N__49157));
    InMux I__10981 (
            .O(N__49160),
            .I(N__49153));
    Span4Mux_v I__10980 (
            .O(N__49157),
            .I(N__49150));
    InMux I__10979 (
            .O(N__49156),
            .I(N__49147));
    LocalMux I__10978 (
            .O(N__49153),
            .I(encoder0_position_target_3));
    Odrv4 I__10977 (
            .O(N__49150),
            .I(encoder0_position_target_3));
    LocalMux I__10976 (
            .O(N__49147),
            .I(encoder0_position_target_3));
    InMux I__10975 (
            .O(N__49140),
            .I(n12438));
    InMux I__10974 (
            .O(N__49137),
            .I(N__49133));
    CascadeMux I__10973 (
            .O(N__49136),
            .I(N__49130));
    LocalMux I__10972 (
            .O(N__49133),
            .I(N__49127));
    InMux I__10971 (
            .O(N__49130),
            .I(N__49122));
    Span4Mux_v I__10970 (
            .O(N__49127),
            .I(N__49119));
    InMux I__10969 (
            .O(N__49126),
            .I(N__49114));
    InMux I__10968 (
            .O(N__49125),
            .I(N__49114));
    LocalMux I__10967 (
            .O(N__49122),
            .I(encoder0_position_target_4));
    Odrv4 I__10966 (
            .O(N__49119),
            .I(encoder0_position_target_4));
    LocalMux I__10965 (
            .O(N__49114),
            .I(encoder0_position_target_4));
    InMux I__10964 (
            .O(N__49107),
            .I(n12439));
    CascadeMux I__10963 (
            .O(N__49104),
            .I(N__49101));
    InMux I__10962 (
            .O(N__49101),
            .I(N__49097));
    CascadeMux I__10961 (
            .O(N__49100),
            .I(N__49094));
    LocalMux I__10960 (
            .O(N__49097),
            .I(N__49091));
    InMux I__10959 (
            .O(N__49094),
            .I(N__49086));
    Span4Mux_h I__10958 (
            .O(N__49091),
            .I(N__49083));
    InMux I__10957 (
            .O(N__49090),
            .I(N__49078));
    InMux I__10956 (
            .O(N__49089),
            .I(N__49078));
    LocalMux I__10955 (
            .O(N__49086),
            .I(encoder0_position_target_5));
    Odrv4 I__10954 (
            .O(N__49083),
            .I(encoder0_position_target_5));
    LocalMux I__10953 (
            .O(N__49078),
            .I(encoder0_position_target_5));
    InMux I__10952 (
            .O(N__49071),
            .I(n12440));
    CascadeMux I__10951 (
            .O(N__49068),
            .I(N__49064));
    CascadeMux I__10950 (
            .O(N__49067),
            .I(N__49061));
    InMux I__10949 (
            .O(N__49064),
            .I(N__49058));
    InMux I__10948 (
            .O(N__49061),
            .I(N__49053));
    LocalMux I__10947 (
            .O(N__49058),
            .I(N__49050));
    CascadeMux I__10946 (
            .O(N__49057),
            .I(N__49047));
    CascadeMux I__10945 (
            .O(N__49056),
            .I(N__49044));
    LocalMux I__10944 (
            .O(N__49053),
            .I(N__49039));
    Span4Mux_h I__10943 (
            .O(N__49050),
            .I(N__49039));
    InMux I__10942 (
            .O(N__49047),
            .I(N__49036));
    InMux I__10941 (
            .O(N__49044),
            .I(N__49033));
    Span4Mux_h I__10940 (
            .O(N__49039),
            .I(N__49030));
    LocalMux I__10939 (
            .O(N__49036),
            .I(encoder0_position_target_6));
    LocalMux I__10938 (
            .O(N__49033),
            .I(encoder0_position_target_6));
    Odrv4 I__10937 (
            .O(N__49030),
            .I(encoder0_position_target_6));
    InMux I__10936 (
            .O(N__49023),
            .I(n12441));
    InMux I__10935 (
            .O(N__49020),
            .I(N__49015));
    InMux I__10934 (
            .O(N__49019),
            .I(N__49012));
    CascadeMux I__10933 (
            .O(N__49018),
            .I(N__49009));
    LocalMux I__10932 (
            .O(N__49015),
            .I(N__49003));
    LocalMux I__10931 (
            .O(N__49012),
            .I(N__49003));
    InMux I__10930 (
            .O(N__49009),
            .I(N__49000));
    InMux I__10929 (
            .O(N__49008),
            .I(N__48997));
    Span4Mux_h I__10928 (
            .O(N__49003),
            .I(N__48994));
    LocalMux I__10927 (
            .O(N__49000),
            .I(encoder0_position_target_7));
    LocalMux I__10926 (
            .O(N__48997),
            .I(encoder0_position_target_7));
    Odrv4 I__10925 (
            .O(N__48994),
            .I(encoder0_position_target_7));
    InMux I__10924 (
            .O(N__48987),
            .I(bfn_15_26_0_));
    CascadeMux I__10923 (
            .O(N__48984),
            .I(N__48981));
    InMux I__10922 (
            .O(N__48981),
            .I(N__48978));
    LocalMux I__10921 (
            .O(N__48978),
            .I(N__48973));
    InMux I__10920 (
            .O(N__48977),
            .I(N__48969));
    InMux I__10919 (
            .O(N__48976),
            .I(N__48966));
    Span4Mux_h I__10918 (
            .O(N__48973),
            .I(N__48963));
    InMux I__10917 (
            .O(N__48972),
            .I(N__48960));
    LocalMux I__10916 (
            .O(N__48969),
            .I(N__48957));
    LocalMux I__10915 (
            .O(N__48966),
            .I(encoder0_position_target_8));
    Odrv4 I__10914 (
            .O(N__48963),
            .I(encoder0_position_target_8));
    LocalMux I__10913 (
            .O(N__48960),
            .I(encoder0_position_target_8));
    Odrv12 I__10912 (
            .O(N__48957),
            .I(encoder0_position_target_8));
    InMux I__10911 (
            .O(N__48948),
            .I(n12443));
    CascadeMux I__10910 (
            .O(N__48945),
            .I(N__48942));
    InMux I__10909 (
            .O(N__48942),
            .I(N__48937));
    CascadeMux I__10908 (
            .O(N__48941),
            .I(N__48934));
    InMux I__10907 (
            .O(N__48940),
            .I(N__48931));
    LocalMux I__10906 (
            .O(N__48937),
            .I(N__48928));
    InMux I__10905 (
            .O(N__48934),
            .I(N__48924));
    LocalMux I__10904 (
            .O(N__48931),
            .I(N__48921));
    Span4Mux_h I__10903 (
            .O(N__48928),
            .I(N__48918));
    InMux I__10902 (
            .O(N__48927),
            .I(N__48915));
    LocalMux I__10901 (
            .O(N__48924),
            .I(N__48910));
    Span4Mux_h I__10900 (
            .O(N__48921),
            .I(N__48910));
    Odrv4 I__10899 (
            .O(N__48918),
            .I(encoder0_position_target_9));
    LocalMux I__10898 (
            .O(N__48915),
            .I(encoder0_position_target_9));
    Odrv4 I__10897 (
            .O(N__48910),
            .I(encoder0_position_target_9));
    InMux I__10896 (
            .O(N__48903),
            .I(n12444));
    CascadeMux I__10895 (
            .O(N__48900),
            .I(N__48897));
    InMux I__10894 (
            .O(N__48897),
            .I(N__48893));
    InMux I__10893 (
            .O(N__48896),
            .I(N__48890));
    LocalMux I__10892 (
            .O(N__48893),
            .I(N__48885));
    LocalMux I__10891 (
            .O(N__48890),
            .I(N__48882));
    InMux I__10890 (
            .O(N__48889),
            .I(N__48879));
    InMux I__10889 (
            .O(N__48888),
            .I(N__48876));
    Span4Mux_v I__10888 (
            .O(N__48885),
            .I(N__48871));
    Span4Mux_h I__10887 (
            .O(N__48882),
            .I(N__48871));
    LocalMux I__10886 (
            .O(N__48879),
            .I(encoder0_position_target_10));
    LocalMux I__10885 (
            .O(N__48876),
            .I(encoder0_position_target_10));
    Odrv4 I__10884 (
            .O(N__48871),
            .I(encoder0_position_target_10));
    InMux I__10883 (
            .O(N__48864),
            .I(n12445));
    InMux I__10882 (
            .O(N__48861),
            .I(n12523));
    InMux I__10881 (
            .O(N__48858),
            .I(bfn_15_24_0_));
    InMux I__10880 (
            .O(N__48855),
            .I(N__48852));
    LocalMux I__10879 (
            .O(N__48852),
            .I(N__48849));
    Odrv4 I__10878 (
            .O(N__48849),
            .I(n1292));
    InMux I__10877 (
            .O(N__48846),
            .I(n12525));
    InMux I__10876 (
            .O(N__48843),
            .I(n12526));
    InMux I__10875 (
            .O(N__48840),
            .I(N__48836));
    InMux I__10874 (
            .O(N__48839),
            .I(N__48833));
    LocalMux I__10873 (
            .O(N__48836),
            .I(N__48828));
    LocalMux I__10872 (
            .O(N__48833),
            .I(N__48828));
    Odrv4 I__10871 (
            .O(N__48828),
            .I(n1323));
    CascadeMux I__10870 (
            .O(N__48825),
            .I(N__48822));
    InMux I__10869 (
            .O(N__48822),
            .I(N__48819));
    LocalMux I__10868 (
            .O(N__48819),
            .I(N__48816));
    Span4Mux_h I__10867 (
            .O(N__48816),
            .I(N__48812));
    InMux I__10866 (
            .O(N__48815),
            .I(N__48808));
    Span4Mux_h I__10865 (
            .O(N__48812),
            .I(N__48805));
    InMux I__10864 (
            .O(N__48811),
            .I(N__48802));
    LocalMux I__10863 (
            .O(N__48808),
            .I(encoder0_position_target_0));
    Odrv4 I__10862 (
            .O(N__48805),
            .I(encoder0_position_target_0));
    LocalMux I__10861 (
            .O(N__48802),
            .I(encoder0_position_target_0));
    InMux I__10860 (
            .O(N__48795),
            .I(n12435));
    CascadeMux I__10859 (
            .O(N__48792),
            .I(N__48789));
    InMux I__10858 (
            .O(N__48789),
            .I(N__48785));
    CascadeMux I__10857 (
            .O(N__48788),
            .I(N__48781));
    LocalMux I__10856 (
            .O(N__48785),
            .I(N__48778));
    CascadeMux I__10855 (
            .O(N__48784),
            .I(N__48775));
    InMux I__10854 (
            .O(N__48781),
            .I(N__48772));
    Span4Mux_h I__10853 (
            .O(N__48778),
            .I(N__48769));
    InMux I__10852 (
            .O(N__48775),
            .I(N__48766));
    LocalMux I__10851 (
            .O(N__48772),
            .I(encoder0_position_target_1));
    Odrv4 I__10850 (
            .O(N__48769),
            .I(encoder0_position_target_1));
    LocalMux I__10849 (
            .O(N__48766),
            .I(encoder0_position_target_1));
    InMux I__10848 (
            .O(N__48759),
            .I(n12436));
    InMux I__10847 (
            .O(N__48756),
            .I(N__48752));
    CascadeMux I__10846 (
            .O(N__48755),
            .I(N__48749));
    LocalMux I__10845 (
            .O(N__48752),
            .I(N__48746));
    InMux I__10844 (
            .O(N__48749),
            .I(N__48742));
    Span4Mux_h I__10843 (
            .O(N__48746),
            .I(N__48739));
    InMux I__10842 (
            .O(N__48745),
            .I(N__48736));
    LocalMux I__10841 (
            .O(N__48742),
            .I(encoder0_position_target_2));
    Odrv4 I__10840 (
            .O(N__48739),
            .I(encoder0_position_target_2));
    LocalMux I__10839 (
            .O(N__48736),
            .I(encoder0_position_target_2));
    InMux I__10838 (
            .O(N__48729),
            .I(n12437));
    CascadeMux I__10837 (
            .O(N__48726),
            .I(N__48722));
    InMux I__10836 (
            .O(N__48725),
            .I(N__48718));
    InMux I__10835 (
            .O(N__48722),
            .I(N__48715));
    InMux I__10834 (
            .O(N__48721),
            .I(N__48712));
    LocalMux I__10833 (
            .O(N__48718),
            .I(n1329));
    LocalMux I__10832 (
            .O(N__48715),
            .I(n1329));
    LocalMux I__10831 (
            .O(N__48712),
            .I(n1329));
    CascadeMux I__10830 (
            .O(N__48705),
            .I(N__48700));
    InMux I__10829 (
            .O(N__48704),
            .I(N__48695));
    InMux I__10828 (
            .O(N__48703),
            .I(N__48695));
    InMux I__10827 (
            .O(N__48700),
            .I(N__48692));
    LocalMux I__10826 (
            .O(N__48695),
            .I(n1333));
    LocalMux I__10825 (
            .O(N__48692),
            .I(n1333));
    InMux I__10824 (
            .O(N__48687),
            .I(N__48682));
    InMux I__10823 (
            .O(N__48686),
            .I(N__48679));
    InMux I__10822 (
            .O(N__48685),
            .I(N__48676));
    LocalMux I__10821 (
            .O(N__48682),
            .I(n298));
    LocalMux I__10820 (
            .O(N__48679),
            .I(n298));
    LocalMux I__10819 (
            .O(N__48676),
            .I(n298));
    InMux I__10818 (
            .O(N__48669),
            .I(N__48666));
    LocalMux I__10817 (
            .O(N__48666),
            .I(n1301));
    InMux I__10816 (
            .O(N__48663),
            .I(bfn_15_23_0_));
    CascadeMux I__10815 (
            .O(N__48660),
            .I(N__48656));
    InMux I__10814 (
            .O(N__48659),
            .I(N__48652));
    InMux I__10813 (
            .O(N__48656),
            .I(N__48649));
    InMux I__10812 (
            .O(N__48655),
            .I(N__48646));
    LocalMux I__10811 (
            .O(N__48652),
            .I(n1233));
    LocalMux I__10810 (
            .O(N__48649),
            .I(n1233));
    LocalMux I__10809 (
            .O(N__48646),
            .I(n1233));
    CascadeMux I__10808 (
            .O(N__48639),
            .I(N__48636));
    InMux I__10807 (
            .O(N__48636),
            .I(N__48633));
    LocalMux I__10806 (
            .O(N__48633),
            .I(n1300));
    InMux I__10805 (
            .O(N__48630),
            .I(n12517));
    CascadeMux I__10804 (
            .O(N__48627),
            .I(N__48624));
    InMux I__10803 (
            .O(N__48624),
            .I(N__48620));
    CascadeMux I__10802 (
            .O(N__48623),
            .I(N__48617));
    LocalMux I__10801 (
            .O(N__48620),
            .I(N__48614));
    InMux I__10800 (
            .O(N__48617),
            .I(N__48611));
    Odrv4 I__10799 (
            .O(N__48614),
            .I(n1232));
    LocalMux I__10798 (
            .O(N__48611),
            .I(n1232));
    InMux I__10797 (
            .O(N__48606),
            .I(N__48603));
    LocalMux I__10796 (
            .O(N__48603),
            .I(N__48600));
    Span4Mux_v I__10795 (
            .O(N__48600),
            .I(N__48597));
    Odrv4 I__10794 (
            .O(N__48597),
            .I(n1299));
    InMux I__10793 (
            .O(N__48594),
            .I(n12518));
    InMux I__10792 (
            .O(N__48591),
            .I(N__48588));
    LocalMux I__10791 (
            .O(N__48588),
            .I(N__48585));
    Odrv4 I__10790 (
            .O(N__48585),
            .I(n1298));
    InMux I__10789 (
            .O(N__48582),
            .I(n12519));
    InMux I__10788 (
            .O(N__48579),
            .I(N__48576));
    LocalMux I__10787 (
            .O(N__48576),
            .I(n1297));
    InMux I__10786 (
            .O(N__48573),
            .I(n12520));
    InMux I__10785 (
            .O(N__48570),
            .I(n12521));
    InMux I__10784 (
            .O(N__48567),
            .I(n12522));
    InMux I__10783 (
            .O(N__48564),
            .I(n12532));
    InMux I__10782 (
            .O(N__48561),
            .I(N__48558));
    LocalMux I__10781 (
            .O(N__48558),
            .I(n1394));
    InMux I__10780 (
            .O(N__48555),
            .I(n12533));
    InMux I__10779 (
            .O(N__48552),
            .I(N__48549));
    LocalMux I__10778 (
            .O(N__48549),
            .I(N__48546));
    Odrv12 I__10777 (
            .O(N__48546),
            .I(n1393));
    InMux I__10776 (
            .O(N__48543),
            .I(bfn_15_22_0_));
    InMux I__10775 (
            .O(N__48540),
            .I(n12535));
    CascadeMux I__10774 (
            .O(N__48537),
            .I(N__48534));
    InMux I__10773 (
            .O(N__48534),
            .I(N__48530));
    InMux I__10772 (
            .O(N__48533),
            .I(N__48527));
    LocalMux I__10771 (
            .O(N__48530),
            .I(n1324));
    LocalMux I__10770 (
            .O(N__48527),
            .I(n1324));
    InMux I__10769 (
            .O(N__48522),
            .I(N__48519));
    LocalMux I__10768 (
            .O(N__48519),
            .I(n1391));
    InMux I__10767 (
            .O(N__48516),
            .I(n12536));
    InMux I__10766 (
            .O(N__48513),
            .I(N__48510));
    LocalMux I__10765 (
            .O(N__48510),
            .I(N__48507));
    Span4Mux_h I__10764 (
            .O(N__48507),
            .I(N__48503));
    CascadeMux I__10763 (
            .O(N__48506),
            .I(N__48500));
    Span4Mux_h I__10762 (
            .O(N__48503),
            .I(N__48497));
    InMux I__10761 (
            .O(N__48500),
            .I(N__48494));
    Odrv4 I__10760 (
            .O(N__48497),
            .I(n15544));
    LocalMux I__10759 (
            .O(N__48494),
            .I(n15544));
    InMux I__10758 (
            .O(N__48489),
            .I(n12537));
    CascadeMux I__10757 (
            .O(N__48486),
            .I(N__48483));
    InMux I__10756 (
            .O(N__48483),
            .I(N__48478));
    CascadeMux I__10755 (
            .O(N__48482),
            .I(N__48475));
    CascadeMux I__10754 (
            .O(N__48481),
            .I(N__48472));
    LocalMux I__10753 (
            .O(N__48478),
            .I(N__48469));
    InMux I__10752 (
            .O(N__48475),
            .I(N__48466));
    InMux I__10751 (
            .O(N__48472),
            .I(N__48463));
    Odrv4 I__10750 (
            .O(N__48469),
            .I(n1332));
    LocalMux I__10749 (
            .O(N__48466),
            .I(n1332));
    LocalMux I__10748 (
            .O(N__48463),
            .I(n1332));
    InMux I__10747 (
            .O(N__48456),
            .I(N__48453));
    LocalMux I__10746 (
            .O(N__48453),
            .I(n13727));
    CascadeMux I__10745 (
            .O(N__48450),
            .I(n14496_cascade_));
    CascadeMux I__10744 (
            .O(N__48447),
            .I(n1455_cascade_));
    CascadeMux I__10743 (
            .O(N__48444),
            .I(N__48441));
    InMux I__10742 (
            .O(N__48441),
            .I(N__48437));
    InMux I__10741 (
            .O(N__48440),
            .I(N__48433));
    LocalMux I__10740 (
            .O(N__48437),
            .I(N__48430));
    InMux I__10739 (
            .O(N__48436),
            .I(N__48427));
    LocalMux I__10738 (
            .O(N__48433),
            .I(n1525));
    Odrv4 I__10737 (
            .O(N__48430),
            .I(n1525));
    LocalMux I__10736 (
            .O(N__48427),
            .I(n1525));
    CascadeMux I__10735 (
            .O(N__48420),
            .I(N__48417));
    InMux I__10734 (
            .O(N__48417),
            .I(N__48413));
    InMux I__10733 (
            .O(N__48416),
            .I(N__48410));
    LocalMux I__10732 (
            .O(N__48413),
            .I(N__48406));
    LocalMux I__10731 (
            .O(N__48410),
            .I(N__48403));
    InMux I__10730 (
            .O(N__48409),
            .I(N__48400));
    Odrv4 I__10729 (
            .O(N__48406),
            .I(n1524));
    Odrv4 I__10728 (
            .O(N__48403),
            .I(n1524));
    LocalMux I__10727 (
            .O(N__48400),
            .I(n1524));
    InMux I__10726 (
            .O(N__48393),
            .I(N__48388));
    InMux I__10725 (
            .O(N__48392),
            .I(N__48383));
    InMux I__10724 (
            .O(N__48391),
            .I(N__48383));
    LocalMux I__10723 (
            .O(N__48388),
            .I(N__48380));
    LocalMux I__10722 (
            .O(N__48383),
            .I(n299));
    Odrv4 I__10721 (
            .O(N__48380),
            .I(n299));
    CascadeMux I__10720 (
            .O(N__48375),
            .I(N__48372));
    InMux I__10719 (
            .O(N__48372),
            .I(N__48369));
    LocalMux I__10718 (
            .O(N__48369),
            .I(n1401));
    InMux I__10717 (
            .O(N__48366),
            .I(bfn_15_21_0_));
    InMux I__10716 (
            .O(N__48363),
            .I(N__48360));
    LocalMux I__10715 (
            .O(N__48360),
            .I(n1400));
    InMux I__10714 (
            .O(N__48357),
            .I(n12527));
    InMux I__10713 (
            .O(N__48354),
            .I(N__48351));
    LocalMux I__10712 (
            .O(N__48351),
            .I(N__48348));
    Odrv4 I__10711 (
            .O(N__48348),
            .I(n1399));
    InMux I__10710 (
            .O(N__48345),
            .I(n12528));
    CascadeMux I__10709 (
            .O(N__48342),
            .I(N__48338));
    CascadeMux I__10708 (
            .O(N__48341),
            .I(N__48335));
    InMux I__10707 (
            .O(N__48338),
            .I(N__48331));
    InMux I__10706 (
            .O(N__48335),
            .I(N__48328));
    InMux I__10705 (
            .O(N__48334),
            .I(N__48325));
    LocalMux I__10704 (
            .O(N__48331),
            .I(N__48322));
    LocalMux I__10703 (
            .O(N__48328),
            .I(n1331));
    LocalMux I__10702 (
            .O(N__48325),
            .I(n1331));
    Odrv4 I__10701 (
            .O(N__48322),
            .I(n1331));
    InMux I__10700 (
            .O(N__48315),
            .I(N__48312));
    LocalMux I__10699 (
            .O(N__48312),
            .I(n1398));
    InMux I__10698 (
            .O(N__48309),
            .I(n12529));
    CascadeMux I__10697 (
            .O(N__48306),
            .I(N__48301));
    InMux I__10696 (
            .O(N__48305),
            .I(N__48298));
    InMux I__10695 (
            .O(N__48304),
            .I(N__48295));
    InMux I__10694 (
            .O(N__48301),
            .I(N__48292));
    LocalMux I__10693 (
            .O(N__48298),
            .I(n1330));
    LocalMux I__10692 (
            .O(N__48295),
            .I(n1330));
    LocalMux I__10691 (
            .O(N__48292),
            .I(n1330));
    CascadeMux I__10690 (
            .O(N__48285),
            .I(N__48282));
    InMux I__10689 (
            .O(N__48282),
            .I(N__48279));
    LocalMux I__10688 (
            .O(N__48279),
            .I(n1397));
    InMux I__10687 (
            .O(N__48276),
            .I(n12530));
    InMux I__10686 (
            .O(N__48273),
            .I(N__48270));
    LocalMux I__10685 (
            .O(N__48270),
            .I(n1396));
    InMux I__10684 (
            .O(N__48267),
            .I(n12531));
    InMux I__10683 (
            .O(N__48264),
            .I(N__48259));
    InMux I__10682 (
            .O(N__48263),
            .I(N__48256));
    InMux I__10681 (
            .O(N__48262),
            .I(N__48253));
    LocalMux I__10680 (
            .O(N__48259),
            .I(n1522));
    LocalMux I__10679 (
            .O(N__48256),
            .I(n1522));
    LocalMux I__10678 (
            .O(N__48253),
            .I(n1522));
    CascadeMux I__10677 (
            .O(N__48246),
            .I(n1523_cascade_));
    InMux I__10676 (
            .O(N__48243),
            .I(N__48240));
    LocalMux I__10675 (
            .O(N__48240),
            .I(n14296));
    InMux I__10674 (
            .O(N__48237),
            .I(N__48234));
    LocalMux I__10673 (
            .O(N__48234),
            .I(N__48231));
    Odrv12 I__10672 (
            .O(N__48231),
            .I(n1601));
    CascadeMux I__10671 (
            .O(N__48228),
            .I(n1554_cascade_));
    InMux I__10670 (
            .O(N__48225),
            .I(N__48220));
    InMux I__10669 (
            .O(N__48224),
            .I(N__48217));
    CascadeMux I__10668 (
            .O(N__48223),
            .I(N__48214));
    LocalMux I__10667 (
            .O(N__48220),
            .I(N__48211));
    LocalMux I__10666 (
            .O(N__48217),
            .I(N__48208));
    InMux I__10665 (
            .O(N__48214),
            .I(N__48205));
    Span4Mux_h I__10664 (
            .O(N__48211),
            .I(N__48200));
    Span4Mux_h I__10663 (
            .O(N__48208),
            .I(N__48200));
    LocalMux I__10662 (
            .O(N__48205),
            .I(N__48197));
    Odrv4 I__10661 (
            .O(N__48200),
            .I(n301));
    Odrv4 I__10660 (
            .O(N__48197),
            .I(n301));
    CascadeMux I__10659 (
            .O(N__48192),
            .I(N__48189));
    InMux I__10658 (
            .O(N__48189),
            .I(N__48185));
    CascadeMux I__10657 (
            .O(N__48188),
            .I(N__48182));
    LocalMux I__10656 (
            .O(N__48185),
            .I(N__48178));
    InMux I__10655 (
            .O(N__48182),
            .I(N__48173));
    InMux I__10654 (
            .O(N__48181),
            .I(N__48173));
    Odrv4 I__10653 (
            .O(N__48178),
            .I(n1633_adj_620));
    LocalMux I__10652 (
            .O(N__48173),
            .I(n1633_adj_620));
    CascadeMux I__10651 (
            .O(N__48168),
            .I(N__48164));
    CascadeMux I__10650 (
            .O(N__48167),
            .I(N__48161));
    InMux I__10649 (
            .O(N__48164),
            .I(N__48157));
    InMux I__10648 (
            .O(N__48161),
            .I(N__48154));
    InMux I__10647 (
            .O(N__48160),
            .I(N__48151));
    LocalMux I__10646 (
            .O(N__48157),
            .I(N__48148));
    LocalMux I__10645 (
            .O(N__48154),
            .I(n1532));
    LocalMux I__10644 (
            .O(N__48151),
            .I(n1532));
    Odrv4 I__10643 (
            .O(N__48148),
            .I(n1532));
    CascadeMux I__10642 (
            .O(N__48141),
            .I(N__48138));
    InMux I__10641 (
            .O(N__48138),
            .I(N__48135));
    LocalMux I__10640 (
            .O(N__48135),
            .I(N__48132));
    Odrv4 I__10639 (
            .O(N__48132),
            .I(n11906));
    CascadeMux I__10638 (
            .O(N__48129),
            .I(n14490_cascade_));
    CascadeMux I__10637 (
            .O(N__48126),
            .I(N__48122));
    CascadeMux I__10636 (
            .O(N__48125),
            .I(N__48119));
    InMux I__10635 (
            .O(N__48122),
            .I(N__48116));
    InMux I__10634 (
            .O(N__48119),
            .I(N__48113));
    LocalMux I__10633 (
            .O(N__48116),
            .I(N__48109));
    LocalMux I__10632 (
            .O(N__48113),
            .I(N__48106));
    InMux I__10631 (
            .O(N__48112),
            .I(N__48103));
    Span4Mux_h I__10630 (
            .O(N__48109),
            .I(N__48100));
    Span4Mux_h I__10629 (
            .O(N__48106),
            .I(N__48097));
    LocalMux I__10628 (
            .O(N__48103),
            .I(n1623_adj_610));
    Odrv4 I__10627 (
            .O(N__48100),
            .I(n1623_adj_610));
    Odrv4 I__10626 (
            .O(N__48097),
            .I(n1623_adj_610));
    CascadeMux I__10625 (
            .O(N__48090),
            .I(N__48087));
    InMux I__10624 (
            .O(N__48087),
            .I(N__48084));
    LocalMux I__10623 (
            .O(N__48084),
            .I(N__48081));
    Span4Mux_v I__10622 (
            .O(N__48081),
            .I(N__48078));
    Odrv4 I__10621 (
            .O(N__48078),
            .I(n1690));
    InMux I__10620 (
            .O(N__48075),
            .I(n12573));
    InMux I__10619 (
            .O(N__48072),
            .I(N__48067));
    CascadeMux I__10618 (
            .O(N__48071),
            .I(N__48064));
    InMux I__10617 (
            .O(N__48070),
            .I(N__48061));
    LocalMux I__10616 (
            .O(N__48067),
            .I(N__48058));
    InMux I__10615 (
            .O(N__48064),
            .I(N__48055));
    LocalMux I__10614 (
            .O(N__48061),
            .I(N__48052));
    Odrv4 I__10613 (
            .O(N__48058),
            .I(n1622_adj_609));
    LocalMux I__10612 (
            .O(N__48055),
            .I(n1622_adj_609));
    Odrv4 I__10611 (
            .O(N__48052),
            .I(n1622_adj_609));
    CascadeMux I__10610 (
            .O(N__48045),
            .I(N__48042));
    InMux I__10609 (
            .O(N__48042),
            .I(N__48039));
    LocalMux I__10608 (
            .O(N__48039),
            .I(N__48036));
    Span4Mux_v I__10607 (
            .O(N__48036),
            .I(N__48033));
    Odrv4 I__10606 (
            .O(N__48033),
            .I(n1689));
    InMux I__10605 (
            .O(N__48030),
            .I(n12574));
    InMux I__10604 (
            .O(N__48027),
            .I(N__48023));
    InMux I__10603 (
            .O(N__48026),
            .I(N__48019));
    LocalMux I__10602 (
            .O(N__48023),
            .I(N__48016));
    InMux I__10601 (
            .O(N__48022),
            .I(N__48013));
    LocalMux I__10600 (
            .O(N__48019),
            .I(N__48010));
    Odrv4 I__10599 (
            .O(N__48016),
            .I(n1621_adj_608));
    LocalMux I__10598 (
            .O(N__48013),
            .I(n1621_adj_608));
    Odrv4 I__10597 (
            .O(N__48010),
            .I(n1621_adj_608));
    InMux I__10596 (
            .O(N__48003),
            .I(N__48000));
    LocalMux I__10595 (
            .O(N__48000),
            .I(N__47997));
    Span4Mux_v I__10594 (
            .O(N__47997),
            .I(N__47994));
    Odrv4 I__10593 (
            .O(N__47994),
            .I(n1688));
    InMux I__10592 (
            .O(N__47991),
            .I(n12575));
    InMux I__10591 (
            .O(N__47988),
            .I(N__47985));
    LocalMux I__10590 (
            .O(N__47985),
            .I(N__47982));
    Span12Mux_h I__10589 (
            .O(N__47982),
            .I(N__47978));
    InMux I__10588 (
            .O(N__47981),
            .I(N__47975));
    Odrv12 I__10587 (
            .O(N__47978),
            .I(n15603));
    LocalMux I__10586 (
            .O(N__47975),
            .I(n15603));
    CascadeMux I__10585 (
            .O(N__47970),
            .I(N__47967));
    InMux I__10584 (
            .O(N__47967),
            .I(N__47964));
    LocalMux I__10583 (
            .O(N__47964),
            .I(N__47960));
    InMux I__10582 (
            .O(N__47963),
            .I(N__47957));
    Span4Mux_h I__10581 (
            .O(N__47960),
            .I(N__47954));
    LocalMux I__10580 (
            .O(N__47957),
            .I(N__47951));
    Odrv4 I__10579 (
            .O(N__47954),
            .I(n1620_adj_607));
    Odrv4 I__10578 (
            .O(N__47951),
            .I(n1620_adj_607));
    InMux I__10577 (
            .O(N__47946),
            .I(n12576));
    CascadeMux I__10576 (
            .O(N__47943),
            .I(N__47939));
    InMux I__10575 (
            .O(N__47942),
            .I(N__47936));
    InMux I__10574 (
            .O(N__47939),
            .I(N__47933));
    LocalMux I__10573 (
            .O(N__47936),
            .I(N__47930));
    LocalMux I__10572 (
            .O(N__47933),
            .I(N__47925));
    Span4Mux_v I__10571 (
            .O(N__47930),
            .I(N__47925));
    Odrv4 I__10570 (
            .O(N__47925),
            .I(n1719));
    InMux I__10569 (
            .O(N__47922),
            .I(N__47919));
    LocalMux I__10568 (
            .O(N__47919),
            .I(n1692));
    CascadeMux I__10567 (
            .O(N__47916),
            .I(N__47913));
    InMux I__10566 (
            .O(N__47913),
            .I(N__47910));
    LocalMux I__10565 (
            .O(N__47910),
            .I(N__47906));
    InMux I__10564 (
            .O(N__47909),
            .I(N__47903));
    Span4Mux_h I__10563 (
            .O(N__47906),
            .I(N__47900));
    LocalMux I__10562 (
            .O(N__47903),
            .I(n1523));
    Odrv4 I__10561 (
            .O(N__47900),
            .I(n1523));
    CascadeMux I__10560 (
            .O(N__47895),
            .I(N__47892));
    InMux I__10559 (
            .O(N__47892),
            .I(N__47888));
    CascadeMux I__10558 (
            .O(N__47891),
            .I(N__47885));
    LocalMux I__10557 (
            .O(N__47888),
            .I(N__47881));
    InMux I__10556 (
            .O(N__47885),
            .I(N__47876));
    InMux I__10555 (
            .O(N__47884),
            .I(N__47876));
    Odrv4 I__10554 (
            .O(N__47881),
            .I(n1632_adj_619));
    LocalMux I__10553 (
            .O(N__47876),
            .I(n1632_adj_619));
    InMux I__10552 (
            .O(N__47871),
            .I(N__47868));
    LocalMux I__10551 (
            .O(N__47868),
            .I(n1699));
    InMux I__10550 (
            .O(N__47865),
            .I(n12564));
    CascadeMux I__10549 (
            .O(N__47862),
            .I(N__47858));
    InMux I__10548 (
            .O(N__47861),
            .I(N__47854));
    InMux I__10547 (
            .O(N__47858),
            .I(N__47851));
    InMux I__10546 (
            .O(N__47857),
            .I(N__47848));
    LocalMux I__10545 (
            .O(N__47854),
            .I(n1631_adj_618));
    LocalMux I__10544 (
            .O(N__47851),
            .I(n1631_adj_618));
    LocalMux I__10543 (
            .O(N__47848),
            .I(n1631_adj_618));
    InMux I__10542 (
            .O(N__47841),
            .I(N__47838));
    LocalMux I__10541 (
            .O(N__47838),
            .I(n1698));
    InMux I__10540 (
            .O(N__47835),
            .I(n12565));
    CascadeMux I__10539 (
            .O(N__47832),
            .I(N__47829));
    InMux I__10538 (
            .O(N__47829),
            .I(N__47825));
    InMux I__10537 (
            .O(N__47828),
            .I(N__47822));
    LocalMux I__10536 (
            .O(N__47825),
            .I(n1630_adj_617));
    LocalMux I__10535 (
            .O(N__47822),
            .I(n1630_adj_617));
    InMux I__10534 (
            .O(N__47817),
            .I(N__47814));
    LocalMux I__10533 (
            .O(N__47814),
            .I(n1697));
    InMux I__10532 (
            .O(N__47811),
            .I(n12566));
    InMux I__10531 (
            .O(N__47808),
            .I(n12567));
    InMux I__10530 (
            .O(N__47805),
            .I(n12568));
    InMux I__10529 (
            .O(N__47802),
            .I(N__47799));
    LocalMux I__10528 (
            .O(N__47799),
            .I(n1694));
    InMux I__10527 (
            .O(N__47796),
            .I(n12569));
    InMux I__10526 (
            .O(N__47793),
            .I(bfn_15_18_0_));
    InMux I__10525 (
            .O(N__47790),
            .I(n12571));
    InMux I__10524 (
            .O(N__47787),
            .I(N__47780));
    InMux I__10523 (
            .O(N__47786),
            .I(N__47780));
    InMux I__10522 (
            .O(N__47785),
            .I(N__47777));
    LocalMux I__10521 (
            .O(N__47780),
            .I(N__47774));
    LocalMux I__10520 (
            .O(N__47777),
            .I(n1624_adj_611));
    Odrv4 I__10519 (
            .O(N__47774),
            .I(n1624_adj_611));
    CascadeMux I__10518 (
            .O(N__47769),
            .I(N__47766));
    InMux I__10517 (
            .O(N__47766),
            .I(N__47763));
    LocalMux I__10516 (
            .O(N__47763),
            .I(n1691));
    InMux I__10515 (
            .O(N__47760),
            .I(n12572));
    InMux I__10514 (
            .O(N__47757),
            .I(N__47753));
    InMux I__10513 (
            .O(N__47756),
            .I(N__47750));
    LocalMux I__10512 (
            .O(N__47753),
            .I(n43));
    LocalMux I__10511 (
            .O(N__47750),
            .I(n43));
    InMux I__10510 (
            .O(N__47745),
            .I(N__47740));
    InMux I__10509 (
            .O(N__47744),
            .I(N__47737));
    InMux I__10508 (
            .O(N__47743),
            .I(N__47734));
    LocalMux I__10507 (
            .O(N__47740),
            .I(n23_adj_668));
    LocalMux I__10506 (
            .O(N__47737),
            .I(n23_adj_668));
    LocalMux I__10505 (
            .O(N__47734),
            .I(n23_adj_668));
    CascadeMux I__10504 (
            .O(N__47727),
            .I(n15132_cascade_));
    InMux I__10503 (
            .O(N__47724),
            .I(N__47719));
    InMux I__10502 (
            .O(N__47723),
            .I(N__47716));
    InMux I__10501 (
            .O(N__47722),
            .I(N__47713));
    LocalMux I__10500 (
            .O(N__47719),
            .I(n25_adj_670));
    LocalMux I__10499 (
            .O(N__47716),
            .I(n25_adj_670));
    LocalMux I__10498 (
            .O(N__47713),
            .I(n25_adj_670));
    InMux I__10497 (
            .O(N__47706),
            .I(N__47703));
    LocalMux I__10496 (
            .O(N__47703),
            .I(N__47700));
    Odrv12 I__10495 (
            .O(N__47700),
            .I(n15110));
    SRMux I__10494 (
            .O(N__47697),
            .I(N__47694));
    LocalMux I__10493 (
            .O(N__47694),
            .I(commutation_state_7__N_261));
    InMux I__10492 (
            .O(N__47691),
            .I(N__47686));
    InMux I__10491 (
            .O(N__47690),
            .I(N__47682));
    InMux I__10490 (
            .O(N__47689),
            .I(N__47679));
    LocalMux I__10489 (
            .O(N__47686),
            .I(N__47676));
    InMux I__10488 (
            .O(N__47685),
            .I(N__47673));
    LocalMux I__10487 (
            .O(N__47682),
            .I(N__47663));
    LocalMux I__10486 (
            .O(N__47679),
            .I(N__47663));
    Span4Mux_s1_v I__10485 (
            .O(N__47676),
            .I(N__47663));
    LocalMux I__10484 (
            .O(N__47673),
            .I(N__47663));
    InMux I__10483 (
            .O(N__47672),
            .I(N__47659));
    Span4Mux_v I__10482 (
            .O(N__47663),
            .I(N__47656));
    InMux I__10481 (
            .O(N__47662),
            .I(N__47653));
    LocalMux I__10480 (
            .O(N__47659),
            .I(N__47650));
    Span4Mux_v I__10479 (
            .O(N__47656),
            .I(N__47647));
    LocalMux I__10478 (
            .O(N__47653),
            .I(N__47640));
    Span12Mux_s9_v I__10477 (
            .O(N__47650),
            .I(N__47640));
    Sp12to4 I__10476 (
            .O(N__47647),
            .I(N__47640));
    Odrv12 I__10475 (
            .O(N__47640),
            .I(h3));
    InMux I__10474 (
            .O(N__47637),
            .I(N__47630));
    InMux I__10473 (
            .O(N__47636),
            .I(N__47627));
    InMux I__10472 (
            .O(N__47635),
            .I(N__47622));
    InMux I__10471 (
            .O(N__47634),
            .I(N__47622));
    InMux I__10470 (
            .O(N__47633),
            .I(N__47618));
    LocalMux I__10469 (
            .O(N__47630),
            .I(N__47611));
    LocalMux I__10468 (
            .O(N__47627),
            .I(N__47611));
    LocalMux I__10467 (
            .O(N__47622),
            .I(N__47611));
    InMux I__10466 (
            .O(N__47621),
            .I(N__47608));
    LocalMux I__10465 (
            .O(N__47618),
            .I(N__47603));
    Span4Mux_v I__10464 (
            .O(N__47611),
            .I(N__47603));
    LocalMux I__10463 (
            .O(N__47608),
            .I(h1));
    Odrv4 I__10462 (
            .O(N__47603),
            .I(h1));
    CascadeMux I__10461 (
            .O(N__47598),
            .I(N__47593));
    InMux I__10460 (
            .O(N__47597),
            .I(N__47590));
    InMux I__10459 (
            .O(N__47596),
            .I(N__47587));
    InMux I__10458 (
            .O(N__47593),
            .I(N__47582));
    LocalMux I__10457 (
            .O(N__47590),
            .I(N__47578));
    LocalMux I__10456 (
            .O(N__47587),
            .I(N__47575));
    InMux I__10455 (
            .O(N__47586),
            .I(N__47570));
    InMux I__10454 (
            .O(N__47585),
            .I(N__47570));
    LocalMux I__10453 (
            .O(N__47582),
            .I(N__47567));
    InMux I__10452 (
            .O(N__47581),
            .I(N__47564));
    Span4Mux_v I__10451 (
            .O(N__47578),
            .I(N__47559));
    Span4Mux_s1_v I__10450 (
            .O(N__47575),
            .I(N__47559));
    LocalMux I__10449 (
            .O(N__47570),
            .I(N__47556));
    Span4Mux_s1_v I__10448 (
            .O(N__47567),
            .I(N__47553));
    LocalMux I__10447 (
            .O(N__47564),
            .I(h2));
    Odrv4 I__10446 (
            .O(N__47559),
            .I(h2));
    Odrv12 I__10445 (
            .O(N__47556),
            .I(h2));
    Odrv4 I__10444 (
            .O(N__47553),
            .I(h2));
    InMux I__10443 (
            .O(N__47544),
            .I(N__47539));
    InMux I__10442 (
            .O(N__47543),
            .I(N__47536));
    InMux I__10441 (
            .O(N__47542),
            .I(N__47533));
    LocalMux I__10440 (
            .O(N__47539),
            .I(N__47530));
    LocalMux I__10439 (
            .O(N__47536),
            .I(N__47527));
    LocalMux I__10438 (
            .O(N__47533),
            .I(N__47524));
    Span4Mux_h I__10437 (
            .O(N__47530),
            .I(N__47519));
    Span4Mux_h I__10436 (
            .O(N__47527),
            .I(N__47519));
    Span4Mux_h I__10435 (
            .O(N__47524),
            .I(N__47516));
    Odrv4 I__10434 (
            .O(N__47519),
            .I(n302));
    Odrv4 I__10433 (
            .O(N__47516),
            .I(n302));
    InMux I__10432 (
            .O(N__47511),
            .I(N__47508));
    LocalMux I__10431 (
            .O(N__47508),
            .I(N__47505));
    Odrv4 I__10430 (
            .O(N__47505),
            .I(n1701));
    InMux I__10429 (
            .O(N__47502),
            .I(bfn_15_17_0_));
    InMux I__10428 (
            .O(N__47499),
            .I(N__47496));
    LocalMux I__10427 (
            .O(N__47496),
            .I(n1700));
    InMux I__10426 (
            .O(N__47493),
            .I(n12563));
    InMux I__10425 (
            .O(N__47490),
            .I(N__47486));
    InMux I__10424 (
            .O(N__47489),
            .I(N__47483));
    LocalMux I__10423 (
            .O(N__47486),
            .I(N__47480));
    LocalMux I__10422 (
            .O(N__47483),
            .I(N__47477));
    Span4Mux_h I__10421 (
            .O(N__47480),
            .I(N__47474));
    Odrv4 I__10420 (
            .O(N__47477),
            .I(pwm_setpoint_4));
    Odrv4 I__10419 (
            .O(N__47474),
            .I(pwm_setpoint_4));
    InMux I__10418 (
            .O(N__47469),
            .I(N__47465));
    InMux I__10417 (
            .O(N__47468),
            .I(N__47462));
    LocalMux I__10416 (
            .O(N__47465),
            .I(N__47459));
    LocalMux I__10415 (
            .O(N__47462),
            .I(pwm_counter_4));
    Odrv4 I__10414 (
            .O(N__47459),
            .I(pwm_counter_4));
    InMux I__10413 (
            .O(N__47454),
            .I(N__47451));
    LocalMux I__10412 (
            .O(N__47451),
            .I(N__47448));
    Odrv4 I__10411 (
            .O(N__47448),
            .I(n15150));
    InMux I__10410 (
            .O(N__47445),
            .I(N__47442));
    LocalMux I__10409 (
            .O(N__47442),
            .I(N__47439));
    Span4Mux_h I__10408 (
            .O(N__47439),
            .I(N__47436));
    Span4Mux_h I__10407 (
            .O(N__47436),
            .I(N__47432));
    InMux I__10406 (
            .O(N__47435),
            .I(N__47429));
    Odrv4 I__10405 (
            .O(N__47432),
            .I(n11_adj_660));
    LocalMux I__10404 (
            .O(N__47429),
            .I(n11_adj_660));
    CascadeMux I__10403 (
            .O(N__47424),
            .I(n9_adj_658_cascade_));
    InMux I__10402 (
            .O(N__47421),
            .I(N__47418));
    LocalMux I__10401 (
            .O(N__47418),
            .I(N__47414));
    InMux I__10400 (
            .O(N__47417),
            .I(N__47411));
    Span4Mux_h I__10399 (
            .O(N__47414),
            .I(N__47408));
    LocalMux I__10398 (
            .O(N__47411),
            .I(n13_adj_662));
    Odrv4 I__10397 (
            .O(N__47408),
            .I(n13_adj_662));
    CascadeMux I__10396 (
            .O(N__47403),
            .I(N__47400));
    InMux I__10395 (
            .O(N__47400),
            .I(N__47397));
    LocalMux I__10394 (
            .O(N__47397),
            .I(N__47394));
    Span4Mux_h I__10393 (
            .O(N__47394),
            .I(N__47391));
    Odrv4 I__10392 (
            .O(N__47391),
            .I(n15_adj_663));
    InMux I__10391 (
            .O(N__47388),
            .I(N__47385));
    LocalMux I__10390 (
            .O(N__47385),
            .I(n15205));
    CascadeMux I__10389 (
            .O(N__47382),
            .I(n15201_cascade_));
    InMux I__10388 (
            .O(N__47379),
            .I(N__47376));
    LocalMux I__10387 (
            .O(N__47376),
            .I(N__47373));
    Span4Mux_v I__10386 (
            .O(N__47373),
            .I(N__47370));
    Span4Mux_h I__10385 (
            .O(N__47370),
            .I(N__47367));
    Odrv4 I__10384 (
            .O(N__47367),
            .I(n15261));
    InMux I__10383 (
            .O(N__47364),
            .I(N__47361));
    LocalMux I__10382 (
            .O(N__47361),
            .I(N__47358));
    Span4Mux_h I__10381 (
            .O(N__47358),
            .I(N__47354));
    InMux I__10380 (
            .O(N__47357),
            .I(N__47351));
    Odrv4 I__10379 (
            .O(N__47354),
            .I(pwm_setpoint_8));
    LocalMux I__10378 (
            .O(N__47351),
            .I(pwm_setpoint_8));
    InMux I__10377 (
            .O(N__47346),
            .I(N__47342));
    InMux I__10376 (
            .O(N__47345),
            .I(N__47339));
    LocalMux I__10375 (
            .O(N__47342),
            .I(N__47334));
    LocalMux I__10374 (
            .O(N__47339),
            .I(N__47331));
    InMux I__10373 (
            .O(N__47338),
            .I(N__47328));
    InMux I__10372 (
            .O(N__47337),
            .I(N__47325));
    Span4Mux_s3_v I__10371 (
            .O(N__47334),
            .I(N__47322));
    Span4Mux_s3_v I__10370 (
            .O(N__47331),
            .I(N__47319));
    LocalMux I__10369 (
            .O(N__47328),
            .I(pwm_counter_8));
    LocalMux I__10368 (
            .O(N__47325),
            .I(pwm_counter_8));
    Odrv4 I__10367 (
            .O(N__47322),
            .I(pwm_counter_8));
    Odrv4 I__10366 (
            .O(N__47319),
            .I(pwm_counter_8));
    CascadeMux I__10365 (
            .O(N__47310),
            .I(N__47307));
    InMux I__10364 (
            .O(N__47307),
            .I(N__47302));
    InMux I__10363 (
            .O(N__47306),
            .I(N__47299));
    InMux I__10362 (
            .O(N__47305),
            .I(N__47296));
    LocalMux I__10361 (
            .O(N__47302),
            .I(N__47291));
    LocalMux I__10360 (
            .O(N__47299),
            .I(N__47291));
    LocalMux I__10359 (
            .O(N__47296),
            .I(N__47288));
    Span4Mux_s1_v I__10358 (
            .O(N__47291),
            .I(N__47285));
    Span4Mux_v I__10357 (
            .O(N__47288),
            .I(N__47282));
    Odrv4 I__10356 (
            .O(N__47285),
            .I(pwm_setpoint_9));
    Odrv4 I__10355 (
            .O(N__47282),
            .I(pwm_setpoint_9));
    InMux I__10354 (
            .O(N__47277),
            .I(N__47273));
    InMux I__10353 (
            .O(N__47276),
            .I(N__47270));
    LocalMux I__10352 (
            .O(N__47273),
            .I(N__47263));
    LocalMux I__10351 (
            .O(N__47270),
            .I(N__47263));
    InMux I__10350 (
            .O(N__47269),
            .I(N__47260));
    InMux I__10349 (
            .O(N__47268),
            .I(N__47257));
    Span4Mux_s3_v I__10348 (
            .O(N__47263),
            .I(N__47254));
    LocalMux I__10347 (
            .O(N__47260),
            .I(pwm_counter_9));
    LocalMux I__10346 (
            .O(N__47257),
            .I(pwm_counter_9));
    Odrv4 I__10345 (
            .O(N__47254),
            .I(pwm_counter_9));
    InMux I__10344 (
            .O(N__47247),
            .I(N__47242));
    InMux I__10343 (
            .O(N__47246),
            .I(N__47239));
    InMux I__10342 (
            .O(N__47245),
            .I(N__47236));
    LocalMux I__10341 (
            .O(N__47242),
            .I(n21_adj_667));
    LocalMux I__10340 (
            .O(N__47239),
            .I(n21_adj_667));
    LocalMux I__10339 (
            .O(N__47236),
            .I(n21_adj_667));
    InMux I__10338 (
            .O(N__47229),
            .I(N__47225));
    InMux I__10337 (
            .O(N__47228),
            .I(N__47222));
    LocalMux I__10336 (
            .O(N__47225),
            .I(n19_adj_666));
    LocalMux I__10335 (
            .O(N__47222),
            .I(n19_adj_666));
    CascadeMux I__10334 (
            .O(N__47217),
            .I(N__47214));
    InMux I__10333 (
            .O(N__47214),
            .I(N__47211));
    LocalMux I__10332 (
            .O(N__47211),
            .I(N__47207));
    InMux I__10331 (
            .O(N__47210),
            .I(N__47204));
    Odrv12 I__10330 (
            .O(N__47207),
            .I(n17_adj_665));
    LocalMux I__10329 (
            .O(N__47204),
            .I(n17_adj_665));
    InMux I__10328 (
            .O(N__47199),
            .I(N__47196));
    LocalMux I__10327 (
            .O(N__47196),
            .I(N__47193));
    Odrv4 I__10326 (
            .O(N__47193),
            .I(n9_adj_658));
    InMux I__10325 (
            .O(N__47190),
            .I(N__47183));
    InMux I__10324 (
            .O(N__47189),
            .I(N__47183));
    InMux I__10323 (
            .O(N__47188),
            .I(N__47180));
    LocalMux I__10322 (
            .O(N__47183),
            .I(N__47173));
    LocalMux I__10321 (
            .O(N__47180),
            .I(N__47173));
    InMux I__10320 (
            .O(N__47179),
            .I(N__47170));
    InMux I__10319 (
            .O(N__47178),
            .I(N__47167));
    Span4Mux_s1_v I__10318 (
            .O(N__47173),
            .I(N__47164));
    LocalMux I__10317 (
            .O(N__47170),
            .I(pwm_counter_21));
    LocalMux I__10316 (
            .O(N__47167),
            .I(pwm_counter_21));
    Odrv4 I__10315 (
            .O(N__47164),
            .I(pwm_counter_21));
    InMux I__10314 (
            .O(N__47157),
            .I(N__47152));
    InMux I__10313 (
            .O(N__47156),
            .I(N__47149));
    InMux I__10312 (
            .O(N__47155),
            .I(N__47146));
    LocalMux I__10311 (
            .O(N__47152),
            .I(N__47143));
    LocalMux I__10310 (
            .O(N__47149),
            .I(pwm_counter_12));
    LocalMux I__10309 (
            .O(N__47146),
            .I(pwm_counter_12));
    Odrv4 I__10308 (
            .O(N__47143),
            .I(pwm_counter_12));
    CascadeMux I__10307 (
            .O(N__47136),
            .I(\PWM.n26_cascade_ ));
    InMux I__10306 (
            .O(N__47133),
            .I(N__47130));
    LocalMux I__10305 (
            .O(N__47130),
            .I(\PWM.n28 ));
    CascadeMux I__10304 (
            .O(N__47127),
            .I(\PWM.n29_cascade_ ));
    InMux I__10303 (
            .O(N__47124),
            .I(N__47121));
    LocalMux I__10302 (
            .O(N__47121),
            .I(\PWM.n27 ));
    SRMux I__10301 (
            .O(N__47118),
            .I(N__47115));
    LocalMux I__10300 (
            .O(N__47115),
            .I(N__47112));
    Span4Mux_v I__10299 (
            .O(N__47112),
            .I(N__47106));
    SRMux I__10298 (
            .O(N__47111),
            .I(N__47103));
    SRMux I__10297 (
            .O(N__47110),
            .I(N__47100));
    SRMux I__10296 (
            .O(N__47109),
            .I(N__47097));
    Odrv4 I__10295 (
            .O(N__47106),
            .I(\PWM.pwm_counter_31__N_407 ));
    LocalMux I__10294 (
            .O(N__47103),
            .I(\PWM.pwm_counter_31__N_407 ));
    LocalMux I__10293 (
            .O(N__47100),
            .I(\PWM.pwm_counter_31__N_407 ));
    LocalMux I__10292 (
            .O(N__47097),
            .I(\PWM.pwm_counter_31__N_407 ));
    InMux I__10291 (
            .O(N__47088),
            .I(N__47083));
    InMux I__10290 (
            .O(N__47087),
            .I(N__47080));
    InMux I__10289 (
            .O(N__47086),
            .I(N__47077));
    LocalMux I__10288 (
            .O(N__47083),
            .I(N__47074));
    LocalMux I__10287 (
            .O(N__47080),
            .I(pwm_counter_19));
    LocalMux I__10286 (
            .O(N__47077),
            .I(pwm_counter_19));
    Odrv12 I__10285 (
            .O(N__47074),
            .I(pwm_counter_19));
    CascadeMux I__10284 (
            .O(N__47067),
            .I(N__47064));
    InMux I__10283 (
            .O(N__47064),
            .I(N__47061));
    LocalMux I__10282 (
            .O(N__47061),
            .I(\PWM.n13995 ));
    InMux I__10281 (
            .O(N__47058),
            .I(N__47055));
    LocalMux I__10280 (
            .O(N__47055),
            .I(\PWM.n17 ));
    InMux I__10279 (
            .O(N__47052),
            .I(N__47048));
    InMux I__10278 (
            .O(N__47051),
            .I(N__47045));
    LocalMux I__10277 (
            .O(N__47048),
            .I(pwm_counter_24));
    LocalMux I__10276 (
            .O(N__47045),
            .I(pwm_counter_24));
    InMux I__10275 (
            .O(N__47040),
            .I(N__47036));
    InMux I__10274 (
            .O(N__47039),
            .I(N__47033));
    LocalMux I__10273 (
            .O(N__47036),
            .I(pwm_counter_29));
    LocalMux I__10272 (
            .O(N__47033),
            .I(pwm_counter_29));
    CascadeMux I__10271 (
            .O(N__47028),
            .I(N__47024));
    InMux I__10270 (
            .O(N__47027),
            .I(N__47021));
    InMux I__10269 (
            .O(N__47024),
            .I(N__47018));
    LocalMux I__10268 (
            .O(N__47021),
            .I(pwm_counter_27));
    LocalMux I__10267 (
            .O(N__47018),
            .I(pwm_counter_27));
    InMux I__10266 (
            .O(N__47013),
            .I(N__47009));
    InMux I__10265 (
            .O(N__47012),
            .I(N__47006));
    LocalMux I__10264 (
            .O(N__47009),
            .I(pwm_counter_26));
    LocalMux I__10263 (
            .O(N__47006),
            .I(pwm_counter_26));
    InMux I__10262 (
            .O(N__47001),
            .I(N__46997));
    InMux I__10261 (
            .O(N__47000),
            .I(N__46994));
    LocalMux I__10260 (
            .O(N__46997),
            .I(pwm_counter_30));
    LocalMux I__10259 (
            .O(N__46994),
            .I(pwm_counter_30));
    InMux I__10258 (
            .O(N__46989),
            .I(N__46985));
    InMux I__10257 (
            .O(N__46988),
            .I(N__46982));
    LocalMux I__10256 (
            .O(N__46985),
            .I(pwm_counter_25));
    LocalMux I__10255 (
            .O(N__46982),
            .I(pwm_counter_25));
    CascadeMux I__10254 (
            .O(N__46977),
            .I(n12_adj_566_cascade_));
    InMux I__10253 (
            .O(N__46974),
            .I(N__46970));
    InMux I__10252 (
            .O(N__46973),
            .I(N__46967));
    LocalMux I__10251 (
            .O(N__46970),
            .I(pwm_counter_28));
    LocalMux I__10250 (
            .O(N__46967),
            .I(pwm_counter_28));
    InMux I__10249 (
            .O(N__46962),
            .I(N__46959));
    LocalMux I__10248 (
            .O(N__46959),
            .I(n5162));
    CascadeMux I__10247 (
            .O(N__46956),
            .I(n5162_cascade_));
    InMux I__10246 (
            .O(N__46953),
            .I(N__46948));
    InMux I__10245 (
            .O(N__46952),
            .I(N__46945));
    InMux I__10244 (
            .O(N__46951),
            .I(N__46942));
    LocalMux I__10243 (
            .O(N__46948),
            .I(pwm_counter_31));
    LocalMux I__10242 (
            .O(N__46945),
            .I(pwm_counter_31));
    LocalMux I__10241 (
            .O(N__46942),
            .I(pwm_counter_31));
    SRMux I__10240 (
            .O(N__46935),
            .I(N__46932));
    LocalMux I__10239 (
            .O(N__46932),
            .I(N__46929));
    Span4Mux_s3_v I__10238 (
            .O(N__46929),
            .I(N__46926));
    Odrv4 I__10237 (
            .O(N__46926),
            .I(n5164));
    InMux I__10236 (
            .O(N__46923),
            .I(N__46920));
    LocalMux I__10235 (
            .O(N__46920),
            .I(N__46917));
    Span4Mux_h I__10234 (
            .O(N__46917),
            .I(N__46914));
    Span4Mux_h I__10233 (
            .O(N__46914),
            .I(N__46911));
    Odrv4 I__10232 (
            .O(N__46911),
            .I(pwm_setpoint_23_N_171_8));
    InMux I__10231 (
            .O(N__46908),
            .I(N__46904));
    InMux I__10230 (
            .O(N__46907),
            .I(N__46901));
    LocalMux I__10229 (
            .O(N__46904),
            .I(N__46898));
    LocalMux I__10228 (
            .O(N__46901),
            .I(N__46895));
    Span4Mux_v I__10227 (
            .O(N__46898),
            .I(N__46892));
    Span4Mux_v I__10226 (
            .O(N__46895),
            .I(N__46889));
    Span4Mux_h I__10225 (
            .O(N__46892),
            .I(N__46886));
    Odrv4 I__10224 (
            .O(N__46889),
            .I(duty_8));
    Odrv4 I__10223 (
            .O(N__46886),
            .I(duty_8));
    CascadeMux I__10222 (
            .O(N__46881),
            .I(n14110_cascade_));
    InMux I__10221 (
            .O(N__46878),
            .I(N__46875));
    LocalMux I__10220 (
            .O(N__46875),
            .I(n10_adj_567));
    InMux I__10219 (
            .O(N__46872),
            .I(N__46869));
    LocalMux I__10218 (
            .O(N__46869),
            .I(n15_adj_702));
    InMux I__10217 (
            .O(N__46866),
            .I(N__46863));
    LocalMux I__10216 (
            .O(N__46863),
            .I(N__46860));
    Odrv4 I__10215 (
            .O(N__46860),
            .I(n11853));
    InMux I__10214 (
            .O(N__46857),
            .I(N__46854));
    LocalMux I__10213 (
            .O(N__46854),
            .I(N__46851));
    Odrv4 I__10212 (
            .O(N__46851),
            .I(n23_adj_562));
    InMux I__10211 (
            .O(N__46848),
            .I(N__46845));
    LocalMux I__10210 (
            .O(N__46845),
            .I(N__46842));
    Span4Mux_h I__10209 (
            .O(N__46842),
            .I(N__46838));
    InMux I__10208 (
            .O(N__46841),
            .I(N__46835));
    Span4Mux_h I__10207 (
            .O(N__46838),
            .I(N__46832));
    LocalMux I__10206 (
            .O(N__46835),
            .I(pwm_setpoint_2));
    Odrv4 I__10205 (
            .O(N__46832),
            .I(pwm_setpoint_2));
    InMux I__10204 (
            .O(N__46827),
            .I(N__46823));
    InMux I__10203 (
            .O(N__46826),
            .I(N__46820));
    LocalMux I__10202 (
            .O(N__46823),
            .I(N__46817));
    LocalMux I__10201 (
            .O(N__46820),
            .I(pwm_setpoint_3));
    Odrv4 I__10200 (
            .O(N__46817),
            .I(pwm_setpoint_3));
    CascadeMux I__10199 (
            .O(N__46812),
            .I(N__46808));
    InMux I__10198 (
            .O(N__46811),
            .I(N__46805));
    InMux I__10197 (
            .O(N__46808),
            .I(N__46802));
    LocalMux I__10196 (
            .O(N__46805),
            .I(pwm_counter_2));
    LocalMux I__10195 (
            .O(N__46802),
            .I(pwm_counter_2));
    InMux I__10194 (
            .O(N__46797),
            .I(N__46794));
    LocalMux I__10193 (
            .O(N__46794),
            .I(N__46790));
    InMux I__10192 (
            .O(N__46793),
            .I(N__46786));
    Span4Mux_v I__10191 (
            .O(N__46790),
            .I(N__46783));
    InMux I__10190 (
            .O(N__46789),
            .I(N__46780));
    LocalMux I__10189 (
            .O(N__46786),
            .I(pwm_counter_3));
    Odrv4 I__10188 (
            .O(N__46783),
            .I(pwm_counter_3));
    LocalMux I__10187 (
            .O(N__46780),
            .I(pwm_counter_3));
    InMux I__10186 (
            .O(N__46773),
            .I(N__46768));
    InMux I__10185 (
            .O(N__46772),
            .I(N__46765));
    InMux I__10184 (
            .O(N__46771),
            .I(N__46762));
    LocalMux I__10183 (
            .O(N__46768),
            .I(N__46759));
    LocalMux I__10182 (
            .O(N__46765),
            .I(pwm_counter_5));
    LocalMux I__10181 (
            .O(N__46762),
            .I(pwm_counter_5));
    Odrv12 I__10180 (
            .O(N__46759),
            .I(pwm_counter_5));
    CascadeMux I__10179 (
            .O(N__46752),
            .I(N__46749));
    InMux I__10178 (
            .O(N__46749),
            .I(N__46745));
    InMux I__10177 (
            .O(N__46748),
            .I(N__46742));
    LocalMux I__10176 (
            .O(N__46745),
            .I(N__46737));
    LocalMux I__10175 (
            .O(N__46742),
            .I(N__46734));
    InMux I__10174 (
            .O(N__46741),
            .I(N__46731));
    InMux I__10173 (
            .O(N__46740),
            .I(N__46728));
    Span4Mux_h I__10172 (
            .O(N__46737),
            .I(N__46725));
    Span4Mux_h I__10171 (
            .O(N__46734),
            .I(N__46722));
    LocalMux I__10170 (
            .O(N__46731),
            .I(pwm_counter_7));
    LocalMux I__10169 (
            .O(N__46728),
            .I(pwm_counter_7));
    Odrv4 I__10168 (
            .O(N__46725),
            .I(pwm_counter_7));
    Odrv4 I__10167 (
            .O(N__46722),
            .I(pwm_counter_7));
    InMux I__10166 (
            .O(N__46713),
            .I(N__46710));
    LocalMux I__10165 (
            .O(N__46710),
            .I(N__46704));
    InMux I__10164 (
            .O(N__46709),
            .I(N__46701));
    InMux I__10163 (
            .O(N__46708),
            .I(N__46698));
    InMux I__10162 (
            .O(N__46707),
            .I(N__46695));
    Span4Mux_h I__10161 (
            .O(N__46704),
            .I(N__46692));
    LocalMux I__10160 (
            .O(N__46701),
            .I(N__46689));
    LocalMux I__10159 (
            .O(N__46698),
            .I(pwm_counter_6));
    LocalMux I__10158 (
            .O(N__46695),
            .I(pwm_counter_6));
    Odrv4 I__10157 (
            .O(N__46692),
            .I(pwm_counter_6));
    Odrv12 I__10156 (
            .O(N__46689),
            .I(pwm_counter_6));
    InMux I__10155 (
            .O(N__46680),
            .I(N__46675));
    InMux I__10154 (
            .O(N__46679),
            .I(N__46672));
    InMux I__10153 (
            .O(N__46678),
            .I(N__46669));
    LocalMux I__10152 (
            .O(N__46675),
            .I(N__46666));
    LocalMux I__10151 (
            .O(N__46672),
            .I(pwm_counter_11));
    LocalMux I__10150 (
            .O(N__46669),
            .I(pwm_counter_11));
    Odrv4 I__10149 (
            .O(N__46666),
            .I(pwm_counter_11));
    InMux I__10148 (
            .O(N__46659),
            .I(N__46654));
    InMux I__10147 (
            .O(N__46658),
            .I(N__46651));
    InMux I__10146 (
            .O(N__46657),
            .I(N__46648));
    LocalMux I__10145 (
            .O(N__46654),
            .I(N__46645));
    LocalMux I__10144 (
            .O(N__46651),
            .I(pwm_counter_10));
    LocalMux I__10143 (
            .O(N__46648),
            .I(pwm_counter_10));
    Odrv4 I__10142 (
            .O(N__46645),
            .I(pwm_counter_10));
    CascadeMux I__10141 (
            .O(N__46638),
            .I(N__46634));
    InMux I__10140 (
            .O(N__46637),
            .I(N__46630));
    InMux I__10139 (
            .O(N__46634),
            .I(N__46627));
    InMux I__10138 (
            .O(N__46633),
            .I(N__46624));
    LocalMux I__10137 (
            .O(N__46630),
            .I(N__46621));
    LocalMux I__10136 (
            .O(N__46627),
            .I(pwm_counter_14));
    LocalMux I__10135 (
            .O(N__46624),
            .I(pwm_counter_14));
    Odrv4 I__10134 (
            .O(N__46621),
            .I(pwm_counter_14));
    InMux I__10133 (
            .O(N__46614),
            .I(N__46609));
    InMux I__10132 (
            .O(N__46613),
            .I(N__46606));
    InMux I__10131 (
            .O(N__46612),
            .I(N__46603));
    LocalMux I__10130 (
            .O(N__46609),
            .I(N__46600));
    LocalMux I__10129 (
            .O(N__46606),
            .I(pwm_counter_20));
    LocalMux I__10128 (
            .O(N__46603),
            .I(pwm_counter_20));
    Odrv4 I__10127 (
            .O(N__46600),
            .I(pwm_counter_20));
    InMux I__10126 (
            .O(N__46593),
            .I(N__46586));
    InMux I__10125 (
            .O(N__46592),
            .I(N__46581));
    InMux I__10124 (
            .O(N__46591),
            .I(N__46581));
    InMux I__10123 (
            .O(N__46590),
            .I(N__46578));
    InMux I__10122 (
            .O(N__46589),
            .I(N__46575));
    LocalMux I__10121 (
            .O(N__46586),
            .I(N__46572));
    LocalMux I__10120 (
            .O(N__46581),
            .I(N__46569));
    LocalMux I__10119 (
            .O(N__46578),
            .I(pwm_counter_16));
    LocalMux I__10118 (
            .O(N__46575),
            .I(pwm_counter_16));
    Odrv12 I__10117 (
            .O(N__46572),
            .I(pwm_counter_16));
    Odrv4 I__10116 (
            .O(N__46569),
            .I(pwm_counter_16));
    InMux I__10115 (
            .O(N__46560),
            .I(N__46555));
    InMux I__10114 (
            .O(N__46559),
            .I(N__46552));
    InMux I__10113 (
            .O(N__46558),
            .I(N__46549));
    LocalMux I__10112 (
            .O(N__46555),
            .I(pwm_counter_17));
    LocalMux I__10111 (
            .O(N__46552),
            .I(pwm_counter_17));
    LocalMux I__10110 (
            .O(N__46549),
            .I(pwm_counter_17));
    CascadeMux I__10109 (
            .O(N__46542),
            .I(N__46538));
    InMux I__10108 (
            .O(N__46541),
            .I(N__46534));
    InMux I__10107 (
            .O(N__46538),
            .I(N__46531));
    InMux I__10106 (
            .O(N__46537),
            .I(N__46528));
    LocalMux I__10105 (
            .O(N__46534),
            .I(N__46525));
    LocalMux I__10104 (
            .O(N__46531),
            .I(pwm_counter_13));
    LocalMux I__10103 (
            .O(N__46528),
            .I(pwm_counter_13));
    Odrv4 I__10102 (
            .O(N__46525),
            .I(pwm_counter_13));
    InMux I__10101 (
            .O(N__46518),
            .I(N__46515));
    LocalMux I__10100 (
            .O(N__46515),
            .I(N__46510));
    InMux I__10099 (
            .O(N__46514),
            .I(N__46507));
    InMux I__10098 (
            .O(N__46513),
            .I(N__46504));
    Odrv4 I__10097 (
            .O(N__46510),
            .I(pwm_counter_23));
    LocalMux I__10096 (
            .O(N__46507),
            .I(pwm_counter_23));
    LocalMux I__10095 (
            .O(N__46504),
            .I(pwm_counter_23));
    InMux I__10094 (
            .O(N__46497),
            .I(N__46492));
    InMux I__10093 (
            .O(N__46496),
            .I(N__46489));
    InMux I__10092 (
            .O(N__46495),
            .I(N__46486));
    LocalMux I__10091 (
            .O(N__46492),
            .I(N__46483));
    LocalMux I__10090 (
            .O(N__46489),
            .I(pwm_counter_22));
    LocalMux I__10089 (
            .O(N__46486),
            .I(pwm_counter_22));
    Odrv4 I__10088 (
            .O(N__46483),
            .I(pwm_counter_22));
    InMux I__10087 (
            .O(N__46476),
            .I(N__46471));
    InMux I__10086 (
            .O(N__46475),
            .I(N__46468));
    InMux I__10085 (
            .O(N__46474),
            .I(N__46465));
    LocalMux I__10084 (
            .O(N__46471),
            .I(N__46462));
    LocalMux I__10083 (
            .O(N__46468),
            .I(pwm_counter_18));
    LocalMux I__10082 (
            .O(N__46465),
            .I(pwm_counter_18));
    Odrv4 I__10081 (
            .O(N__46462),
            .I(pwm_counter_18));
    CascadeMux I__10080 (
            .O(N__46455),
            .I(N__46451));
    InMux I__10079 (
            .O(N__46454),
            .I(N__46448));
    InMux I__10078 (
            .O(N__46451),
            .I(N__46445));
    LocalMux I__10077 (
            .O(N__46448),
            .I(N__46441));
    LocalMux I__10076 (
            .O(N__46445),
            .I(N__46438));
    InMux I__10075 (
            .O(N__46444),
            .I(N__46435));
    Span4Mux_v I__10074 (
            .O(N__46441),
            .I(N__46432));
    Odrv4 I__10073 (
            .O(N__46438),
            .I(pwm_counter_15));
    LocalMux I__10072 (
            .O(N__46435),
            .I(pwm_counter_15));
    Odrv4 I__10071 (
            .O(N__46432),
            .I(pwm_counter_15));
    InMux I__10070 (
            .O(N__46425),
            .I(N__46421));
    CascadeMux I__10069 (
            .O(N__46424),
            .I(N__46415));
    LocalMux I__10068 (
            .O(N__46421),
            .I(N__46411));
    CascadeMux I__10067 (
            .O(N__46420),
            .I(N__46405));
    InMux I__10066 (
            .O(N__46419),
            .I(N__46399));
    InMux I__10065 (
            .O(N__46418),
            .I(N__46399));
    InMux I__10064 (
            .O(N__46415),
            .I(N__46394));
    InMux I__10063 (
            .O(N__46414),
            .I(N__46394));
    Span12Mux_h I__10062 (
            .O(N__46411),
            .I(N__46391));
    InMux I__10061 (
            .O(N__46410),
            .I(N__46388));
    InMux I__10060 (
            .O(N__46409),
            .I(N__46385));
    InMux I__10059 (
            .O(N__46408),
            .I(N__46382));
    InMux I__10058 (
            .O(N__46405),
            .I(N__46377));
    InMux I__10057 (
            .O(N__46404),
            .I(N__46377));
    LocalMux I__10056 (
            .O(N__46399),
            .I(N__46374));
    LocalMux I__10055 (
            .O(N__46394),
            .I(N__46371));
    Odrv12 I__10054 (
            .O(N__46391),
            .I(n1059));
    LocalMux I__10053 (
            .O(N__46388),
            .I(n1059));
    LocalMux I__10052 (
            .O(N__46385),
            .I(n1059));
    LocalMux I__10051 (
            .O(N__46382),
            .I(n1059));
    LocalMux I__10050 (
            .O(N__46377),
            .I(n1059));
    Odrv4 I__10049 (
            .O(N__46374),
            .I(n1059));
    Odrv4 I__10048 (
            .O(N__46371),
            .I(n1059));
    InMux I__10047 (
            .O(N__46356),
            .I(N__46353));
    LocalMux I__10046 (
            .O(N__46353),
            .I(N__46350));
    Span4Mux_h I__10045 (
            .O(N__46350),
            .I(N__46347));
    Span4Mux_h I__10044 (
            .O(N__46347),
            .I(N__46344));
    Odrv4 I__10043 (
            .O(N__46344),
            .I(n15499));
    InMux I__10042 (
            .O(N__46341),
            .I(N__46338));
    LocalMux I__10041 (
            .O(N__46338),
            .I(n14470));
    InMux I__10040 (
            .O(N__46335),
            .I(N__46332));
    LocalMux I__10039 (
            .O(N__46332),
            .I(N__46328));
    CascadeMux I__10038 (
            .O(N__46331),
            .I(N__46324));
    Span4Mux_v I__10037 (
            .O(N__46328),
            .I(N__46321));
    InMux I__10036 (
            .O(N__46327),
            .I(N__46318));
    InMux I__10035 (
            .O(N__46324),
            .I(N__46315));
    Sp12to4 I__10034 (
            .O(N__46321),
            .I(N__46310));
    LocalMux I__10033 (
            .O(N__46318),
            .I(N__46310));
    LocalMux I__10032 (
            .O(N__46315),
            .I(encoder0_position_21));
    Odrv12 I__10031 (
            .O(N__46310),
            .I(encoder0_position_21));
    CascadeMux I__10030 (
            .O(N__46305),
            .I(N__46302));
    InMux I__10029 (
            .O(N__46302),
            .I(N__46299));
    LocalMux I__10028 (
            .O(N__46299),
            .I(N__46296));
    Span4Mux_h I__10027 (
            .O(N__46296),
            .I(N__46293));
    Odrv4 I__10026 (
            .O(N__46293),
            .I(n12_adj_633));
    CascadeMux I__10025 (
            .O(N__46290),
            .I(n16_adj_701_cascade_));
    InMux I__10024 (
            .O(N__46287),
            .I(N__46284));
    LocalMux I__10023 (
            .O(N__46284),
            .I(N__46281));
    Odrv12 I__10022 (
            .O(N__46281),
            .I(n24_adj_561));
    InMux I__10021 (
            .O(N__46278),
            .I(N__46275));
    LocalMux I__10020 (
            .O(N__46275),
            .I(N__46272));
    Odrv4 I__10019 (
            .O(N__46272),
            .I(n25));
    CascadeMux I__10018 (
            .O(N__46269),
            .I(n13932_cascade_));
    InMux I__10017 (
            .O(N__46266),
            .I(N__46261));
    InMux I__10016 (
            .O(N__46265),
            .I(N__46258));
    InMux I__10015 (
            .O(N__46264),
            .I(N__46255));
    LocalMux I__10014 (
            .O(N__46261),
            .I(N__46252));
    LocalMux I__10013 (
            .O(N__46258),
            .I(N__46247));
    LocalMux I__10012 (
            .O(N__46255),
            .I(N__46247));
    Span4Mux_h I__10011 (
            .O(N__46252),
            .I(N__46244));
    Odrv4 I__10010 (
            .O(N__46247),
            .I(n296));
    Odrv4 I__10009 (
            .O(N__46244),
            .I(n296));
    CascadeMux I__10008 (
            .O(N__46239),
            .I(N__46236));
    InMux I__10007 (
            .O(N__46236),
            .I(N__46233));
    LocalMux I__10006 (
            .O(N__46233),
            .I(N__46230));
    Odrv4 I__10005 (
            .O(N__46230),
            .I(n1101));
    CascadeMux I__10004 (
            .O(N__46227),
            .I(n1133_cascade_));
    InMux I__10003 (
            .O(N__46224),
            .I(N__46221));
    LocalMux I__10002 (
            .O(N__46221),
            .I(n14428));
    CascadeMux I__10001 (
            .O(N__46218),
            .I(n12000_cascade_));
    CascadeMux I__10000 (
            .O(N__46215),
            .I(n1158_cascade_));
    CascadeMux I__9999 (
            .O(N__46212),
            .I(n1232_cascade_));
    InMux I__9998 (
            .O(N__46209),
            .I(N__46206));
    LocalMux I__9997 (
            .O(N__46206),
            .I(N__46203));
    Odrv12 I__9996 (
            .O(N__46203),
            .I(n12));
    InMux I__9995 (
            .O(N__46200),
            .I(N__46177));
    CascadeMux I__9994 (
            .O(N__46199),
            .I(N__46174));
    InMux I__9993 (
            .O(N__46198),
            .I(N__46166));
    InMux I__9992 (
            .O(N__46197),
            .I(N__46166));
    InMux I__9991 (
            .O(N__46196),
            .I(N__46166));
    CascadeMux I__9990 (
            .O(N__46195),
            .I(N__46161));
    InMux I__9989 (
            .O(N__46194),
            .I(N__46155));
    InMux I__9988 (
            .O(N__46193),
            .I(N__46145));
    InMux I__9987 (
            .O(N__46192),
            .I(N__46145));
    InMux I__9986 (
            .O(N__46191),
            .I(N__46142));
    InMux I__9985 (
            .O(N__46190),
            .I(N__46133));
    InMux I__9984 (
            .O(N__46189),
            .I(N__46133));
    InMux I__9983 (
            .O(N__46188),
            .I(N__46133));
    InMux I__9982 (
            .O(N__46187),
            .I(N__46133));
    InMux I__9981 (
            .O(N__46186),
            .I(N__46124));
    InMux I__9980 (
            .O(N__46185),
            .I(N__46124));
    InMux I__9979 (
            .O(N__46184),
            .I(N__46124));
    InMux I__9978 (
            .O(N__46183),
            .I(N__46124));
    InMux I__9977 (
            .O(N__46182),
            .I(N__46121));
    InMux I__9976 (
            .O(N__46181),
            .I(N__46118));
    InMux I__9975 (
            .O(N__46180),
            .I(N__46115));
    LocalMux I__9974 (
            .O(N__46177),
            .I(N__46112));
    InMux I__9973 (
            .O(N__46174),
            .I(N__46107));
    InMux I__9972 (
            .O(N__46173),
            .I(N__46107));
    LocalMux I__9971 (
            .O(N__46166),
            .I(N__46104));
    CascadeMux I__9970 (
            .O(N__46165),
            .I(N__46099));
    InMux I__9969 (
            .O(N__46164),
            .I(N__46091));
    InMux I__9968 (
            .O(N__46161),
            .I(N__46091));
    InMux I__9967 (
            .O(N__46160),
            .I(N__46091));
    InMux I__9966 (
            .O(N__46159),
            .I(N__46086));
    InMux I__9965 (
            .O(N__46158),
            .I(N__46086));
    LocalMux I__9964 (
            .O(N__46155),
            .I(N__46083));
    InMux I__9963 (
            .O(N__46154),
            .I(N__46076));
    InMux I__9962 (
            .O(N__46153),
            .I(N__46076));
    InMux I__9961 (
            .O(N__46152),
            .I(N__46076));
    InMux I__9960 (
            .O(N__46151),
            .I(N__46071));
    InMux I__9959 (
            .O(N__46150),
            .I(N__46071));
    LocalMux I__9958 (
            .O(N__46145),
            .I(N__46062));
    LocalMux I__9957 (
            .O(N__46142),
            .I(N__46062));
    LocalMux I__9956 (
            .O(N__46133),
            .I(N__46062));
    LocalMux I__9955 (
            .O(N__46124),
            .I(N__46062));
    LocalMux I__9954 (
            .O(N__46121),
            .I(N__46057));
    LocalMux I__9953 (
            .O(N__46118),
            .I(N__46054));
    LocalMux I__9952 (
            .O(N__46115),
            .I(N__46050));
    Span4Mux_v I__9951 (
            .O(N__46112),
            .I(N__46047));
    LocalMux I__9950 (
            .O(N__46107),
            .I(N__46044));
    Span4Mux_v I__9949 (
            .O(N__46104),
            .I(N__46041));
    InMux I__9948 (
            .O(N__46103),
            .I(N__46032));
    InMux I__9947 (
            .O(N__46102),
            .I(N__46032));
    InMux I__9946 (
            .O(N__46099),
            .I(N__46032));
    InMux I__9945 (
            .O(N__46098),
            .I(N__46032));
    LocalMux I__9944 (
            .O(N__46091),
            .I(N__46024));
    LocalMux I__9943 (
            .O(N__46086),
            .I(N__46024));
    Span4Mux_v I__9942 (
            .O(N__46083),
            .I(N__46021));
    LocalMux I__9941 (
            .O(N__46076),
            .I(N__46018));
    LocalMux I__9940 (
            .O(N__46071),
            .I(N__46013));
    Span4Mux_h I__9939 (
            .O(N__46062),
            .I(N__46013));
    InMux I__9938 (
            .O(N__46061),
            .I(N__46010));
    InMux I__9937 (
            .O(N__46060),
            .I(N__46007));
    Span4Mux_h I__9936 (
            .O(N__46057),
            .I(N__46004));
    Span12Mux_v I__9935 (
            .O(N__46054),
            .I(N__46001));
    InMux I__9934 (
            .O(N__46053),
            .I(N__45998));
    Span4Mux_v I__9933 (
            .O(N__46050),
            .I(N__45987));
    Span4Mux_h I__9932 (
            .O(N__46047),
            .I(N__45987));
    Span4Mux_v I__9931 (
            .O(N__46044),
            .I(N__45987));
    Span4Mux_v I__9930 (
            .O(N__46041),
            .I(N__45987));
    LocalMux I__9929 (
            .O(N__46032),
            .I(N__45987));
    InMux I__9928 (
            .O(N__46031),
            .I(N__45980));
    InMux I__9927 (
            .O(N__46030),
            .I(N__45980));
    InMux I__9926 (
            .O(N__46029),
            .I(N__45980));
    Span4Mux_v I__9925 (
            .O(N__46024),
            .I(N__45971));
    Span4Mux_h I__9924 (
            .O(N__46021),
            .I(N__45971));
    Span4Mux_v I__9923 (
            .O(N__46018),
            .I(N__45971));
    Span4Mux_v I__9922 (
            .O(N__46013),
            .I(N__45971));
    LocalMux I__9921 (
            .O(N__46010),
            .I(encoder0_position_31));
    LocalMux I__9920 (
            .O(N__46007),
            .I(encoder0_position_31));
    Odrv4 I__9919 (
            .O(N__46004),
            .I(encoder0_position_31));
    Odrv12 I__9918 (
            .O(N__46001),
            .I(encoder0_position_31));
    LocalMux I__9917 (
            .O(N__45998),
            .I(encoder0_position_31));
    Odrv4 I__9916 (
            .O(N__45987),
            .I(encoder0_position_31));
    LocalMux I__9915 (
            .O(N__45980),
            .I(encoder0_position_31));
    Odrv4 I__9914 (
            .O(N__45971),
            .I(encoder0_position_31));
    InMux I__9913 (
            .O(N__45954),
            .I(N__45951));
    LocalMux I__9912 (
            .O(N__45951),
            .I(n1100));
    CascadeMux I__9911 (
            .O(N__45948),
            .I(N__45945));
    InMux I__9910 (
            .O(N__45945),
            .I(N__45942));
    LocalMux I__9909 (
            .O(N__45942),
            .I(N__45938));
    CascadeMux I__9908 (
            .O(N__45941),
            .I(N__45935));
    Span4Mux_h I__9907 (
            .O(N__45938),
            .I(N__45931));
    InMux I__9906 (
            .O(N__45935),
            .I(N__45928));
    InMux I__9905 (
            .O(N__45934),
            .I(N__45925));
    Odrv4 I__9904 (
            .O(N__45931),
            .I(n1033));
    LocalMux I__9903 (
            .O(N__45928),
            .I(n1033));
    LocalMux I__9902 (
            .O(N__45925),
            .I(n1033));
    CascadeMux I__9901 (
            .O(N__45918),
            .I(n1132_cascade_));
    CascadeMux I__9900 (
            .O(N__45915),
            .I(N__45911));
    InMux I__9899 (
            .O(N__45914),
            .I(N__45908));
    InMux I__9898 (
            .O(N__45911),
            .I(N__45905));
    LocalMux I__9897 (
            .O(N__45908),
            .I(n1032));
    LocalMux I__9896 (
            .O(N__45905),
            .I(n1032));
    CascadeMux I__9895 (
            .O(N__45900),
            .I(N__45897));
    InMux I__9894 (
            .O(N__45897),
            .I(N__45894));
    LocalMux I__9893 (
            .O(N__45894),
            .I(n1099));
    CascadeMux I__9892 (
            .O(N__45891),
            .I(n11908_cascade_));
    CascadeMux I__9891 (
            .O(N__45888),
            .I(n13708_cascade_));
    CascadeMux I__9890 (
            .O(N__45885),
            .I(n1356_cascade_));
    CascadeMux I__9889 (
            .O(N__45882),
            .I(n1433_cascade_));
    InMux I__9888 (
            .O(N__45879),
            .I(N__45876));
    LocalMux I__9887 (
            .O(N__45876),
            .I(N__45871));
    CascadeMux I__9886 (
            .O(N__45875),
            .I(N__45868));
    InMux I__9885 (
            .O(N__45874),
            .I(N__45865));
    Span4Mux_h I__9884 (
            .O(N__45871),
            .I(N__45862));
    InMux I__9883 (
            .O(N__45868),
            .I(N__45859));
    LocalMux I__9882 (
            .O(N__45865),
            .I(N__45856));
    Odrv4 I__9881 (
            .O(N__45862),
            .I(n1031));
    LocalMux I__9880 (
            .O(N__45859),
            .I(n1031));
    Odrv4 I__9879 (
            .O(N__45856),
            .I(n1031));
    InMux I__9878 (
            .O(N__45849),
            .I(N__45846));
    LocalMux I__9877 (
            .O(N__45846),
            .I(n1098));
    CascadeMux I__9876 (
            .O(N__45843),
            .I(n1527_cascade_));
    InMux I__9875 (
            .O(N__45840),
            .I(N__45837));
    LocalMux I__9874 (
            .O(N__45837),
            .I(n14288));
    InMux I__9873 (
            .O(N__45834),
            .I(N__45831));
    LocalMux I__9872 (
            .O(N__45831),
            .I(N__45828));
    Span4Mux_v I__9871 (
            .O(N__45828),
            .I(N__45825));
    Span4Mux_h I__9870 (
            .O(N__45825),
            .I(N__45822));
    Odrv4 I__9869 (
            .O(N__45822),
            .I(n14));
    CascadeMux I__9868 (
            .O(N__45819),
            .I(n1324_cascade_));
    InMux I__9867 (
            .O(N__45816),
            .I(N__45810));
    InMux I__9866 (
            .O(N__45815),
            .I(N__45810));
    LocalMux I__9865 (
            .O(N__45810),
            .I(N__45806));
    CascadeMux I__9864 (
            .O(N__45809),
            .I(N__45803));
    Span4Mux_h I__9863 (
            .O(N__45806),
            .I(N__45800));
    InMux I__9862 (
            .O(N__45803),
            .I(N__45797));
    Span4Mux_h I__9861 (
            .O(N__45800),
            .I(N__45794));
    LocalMux I__9860 (
            .O(N__45797),
            .I(encoder0_position_19));
    Odrv4 I__9859 (
            .O(N__45794),
            .I(encoder0_position_19));
    CascadeMux I__9858 (
            .O(N__45789),
            .I(N__45786));
    InMux I__9857 (
            .O(N__45786),
            .I(N__45783));
    LocalMux I__9856 (
            .O(N__45783),
            .I(N__45780));
    Span4Mux_h I__9855 (
            .O(N__45780),
            .I(N__45777));
    Odrv4 I__9854 (
            .O(N__45777),
            .I(n14_adj_635));
    CascadeMux I__9853 (
            .O(N__45774),
            .I(n1531_cascade_));
    CascadeMux I__9852 (
            .O(N__45771),
            .I(N__45768));
    InMux I__9851 (
            .O(N__45768),
            .I(N__45765));
    LocalMux I__9850 (
            .O(N__45765),
            .I(n1592));
    CascadeMux I__9849 (
            .O(N__45762),
            .I(N__45758));
    InMux I__9848 (
            .O(N__45761),
            .I(N__45755));
    InMux I__9847 (
            .O(N__45758),
            .I(N__45752));
    LocalMux I__9846 (
            .O(N__45755),
            .I(n1533));
    LocalMux I__9845 (
            .O(N__45752),
            .I(n1533));
    InMux I__9844 (
            .O(N__45747),
            .I(N__45744));
    LocalMux I__9843 (
            .O(N__45744),
            .I(n1600));
    CascadeMux I__9842 (
            .O(N__45741),
            .I(n1533_cascade_));
    InMux I__9841 (
            .O(N__45738),
            .I(N__45735));
    LocalMux I__9840 (
            .O(N__45735),
            .I(N__45732));
    Span4Mux_h I__9839 (
            .O(N__45732),
            .I(N__45729));
    Span4Mux_h I__9838 (
            .O(N__45729),
            .I(N__45726));
    Span4Mux_v I__9837 (
            .O(N__45726),
            .I(N__45722));
    InMux I__9836 (
            .O(N__45725),
            .I(N__45719));
    Odrv4 I__9835 (
            .O(N__45722),
            .I(n15582));
    LocalMux I__9834 (
            .O(N__45719),
            .I(n15582));
    CascadeMux I__9833 (
            .O(N__45714),
            .I(n14294_cascade_));
    InMux I__9832 (
            .O(N__45711),
            .I(N__45708));
    LocalMux I__9831 (
            .O(N__45708),
            .I(n11974));
    CascadeMux I__9830 (
            .O(N__45705),
            .I(n11902_cascade_));
    InMux I__9829 (
            .O(N__45702),
            .I(N__45699));
    LocalMux I__9828 (
            .O(N__45699),
            .I(n13736));
    InMux I__9827 (
            .O(N__45696),
            .I(N__45693));
    LocalMux I__9826 (
            .O(N__45693),
            .I(n1599));
    InMux I__9825 (
            .O(N__45690),
            .I(N__45687));
    LocalMux I__9824 (
            .O(N__45687),
            .I(N__45683));
    CascadeMux I__9823 (
            .O(N__45686),
            .I(N__45680));
    Span4Mux_v I__9822 (
            .O(N__45683),
            .I(N__45677));
    InMux I__9821 (
            .O(N__45680),
            .I(N__45674));
    Odrv4 I__9820 (
            .O(N__45677),
            .I(n1731));
    LocalMux I__9819 (
            .O(N__45674),
            .I(n1731));
    InMux I__9818 (
            .O(N__45669),
            .I(N__45666));
    LocalMux I__9817 (
            .O(N__45666),
            .I(N__45662));
    CascadeMux I__9816 (
            .O(N__45665),
            .I(N__45659));
    Span4Mux_h I__9815 (
            .O(N__45662),
            .I(N__45655));
    InMux I__9814 (
            .O(N__45659),
            .I(N__45652));
    InMux I__9813 (
            .O(N__45658),
            .I(N__45649));
    Odrv4 I__9812 (
            .O(N__45655),
            .I(n1733));
    LocalMux I__9811 (
            .O(N__45652),
            .I(n1733));
    LocalMux I__9810 (
            .O(N__45649),
            .I(n1733));
    InMux I__9809 (
            .O(N__45642),
            .I(N__45638));
    InMux I__9808 (
            .O(N__45641),
            .I(N__45635));
    LocalMux I__9807 (
            .O(N__45638),
            .I(N__45631));
    LocalMux I__9806 (
            .O(N__45635),
            .I(N__45628));
    InMux I__9805 (
            .O(N__45634),
            .I(N__45625));
    Span4Mux_h I__9804 (
            .O(N__45631),
            .I(N__45622));
    Span4Mux_v I__9803 (
            .O(N__45628),
            .I(N__45619));
    LocalMux I__9802 (
            .O(N__45625),
            .I(n303));
    Odrv4 I__9801 (
            .O(N__45622),
            .I(n303));
    Odrv4 I__9800 (
            .O(N__45619),
            .I(n303));
    CascadeMux I__9799 (
            .O(N__45612),
            .I(n1731_cascade_));
    InMux I__9798 (
            .O(N__45609),
            .I(N__45606));
    LocalMux I__9797 (
            .O(N__45606),
            .I(N__45603));
    Span4Mux_h I__9796 (
            .O(N__45603),
            .I(N__45600));
    Odrv4 I__9795 (
            .O(N__45600),
            .I(n11970));
    InMux I__9794 (
            .O(N__45597),
            .I(N__45594));
    LocalMux I__9793 (
            .O(N__45594),
            .I(N__45590));
    CascadeMux I__9792 (
            .O(N__45593),
            .I(N__45587));
    Span4Mux_h I__9791 (
            .O(N__45590),
            .I(N__45583));
    InMux I__9790 (
            .O(N__45587),
            .I(N__45580));
    InMux I__9789 (
            .O(N__45586),
            .I(N__45577));
    Odrv4 I__9788 (
            .O(N__45583),
            .I(n1732));
    LocalMux I__9787 (
            .O(N__45580),
            .I(n1732));
    LocalMux I__9786 (
            .O(N__45577),
            .I(n1732));
    InMux I__9785 (
            .O(N__45570),
            .I(N__45567));
    LocalMux I__9784 (
            .O(N__45567),
            .I(n1590));
    InMux I__9783 (
            .O(N__45564),
            .I(N__45561));
    LocalMux I__9782 (
            .O(N__45561),
            .I(n1589));
    CascadeMux I__9781 (
            .O(N__45558),
            .I(N__45554));
    CascadeMux I__9780 (
            .O(N__45557),
            .I(N__45551));
    InMux I__9779 (
            .O(N__45554),
            .I(N__45548));
    InMux I__9778 (
            .O(N__45551),
            .I(N__45545));
    LocalMux I__9777 (
            .O(N__45548),
            .I(n1531));
    LocalMux I__9776 (
            .O(N__45545),
            .I(n1531));
    CascadeMux I__9775 (
            .O(N__45540),
            .I(n14910_cascade_));
    InMux I__9774 (
            .O(N__45537),
            .I(N__45532));
    CascadeMux I__9773 (
            .O(N__45536),
            .I(N__45529));
    InMux I__9772 (
            .O(N__45535),
            .I(N__45526));
    LocalMux I__9771 (
            .O(N__45532),
            .I(N__45523));
    InMux I__9770 (
            .O(N__45529),
            .I(N__45520));
    LocalMux I__9769 (
            .O(N__45526),
            .I(N__45515));
    Span4Mux_v I__9768 (
            .O(N__45523),
            .I(N__45515));
    LocalMux I__9767 (
            .O(N__45520),
            .I(n1730));
    Odrv4 I__9766 (
            .O(N__45515),
            .I(n1730));
    CascadeMux I__9765 (
            .O(N__45510),
            .I(n14514_cascade_));
    CascadeMux I__9764 (
            .O(N__45507),
            .I(n1653_cascade_));
    InMux I__9763 (
            .O(N__45504),
            .I(N__45501));
    LocalMux I__9762 (
            .O(N__45501),
            .I(n1598));
    CascadeMux I__9761 (
            .O(N__45498),
            .I(n1630_adj_617_cascade_));
    CascadeMux I__9760 (
            .O(N__45495),
            .I(N__45490));
    CascadeMux I__9759 (
            .O(N__45494),
            .I(N__45487));
    InMux I__9758 (
            .O(N__45493),
            .I(N__45482));
    InMux I__9757 (
            .O(N__45490),
            .I(N__45482));
    InMux I__9756 (
            .O(N__45487),
            .I(N__45479));
    LocalMux I__9755 (
            .O(N__45482),
            .I(N__45476));
    LocalMux I__9754 (
            .O(N__45479),
            .I(n1729));
    Odrv12 I__9753 (
            .O(N__45476),
            .I(n1729));
    InMux I__9752 (
            .O(N__45471),
            .I(N__45467));
    InMux I__9751 (
            .O(N__45470),
            .I(N__45464));
    LocalMux I__9750 (
            .O(N__45467),
            .I(pwm_setpoint_11));
    LocalMux I__9749 (
            .O(N__45464),
            .I(pwm_setpoint_11));
    InMux I__9748 (
            .O(N__45459),
            .I(N__45455));
    InMux I__9747 (
            .O(N__45458),
            .I(N__45452));
    LocalMux I__9746 (
            .O(N__45455),
            .I(N__45449));
    LocalMux I__9745 (
            .O(N__45452),
            .I(pwm_setpoint_12));
    Odrv4 I__9744 (
            .O(N__45449),
            .I(pwm_setpoint_12));
    InMux I__9743 (
            .O(N__45444),
            .I(N__45440));
    InMux I__9742 (
            .O(N__45443),
            .I(N__45437));
    LocalMux I__9741 (
            .O(N__45440),
            .I(pwm_setpoint_20));
    LocalMux I__9740 (
            .O(N__45437),
            .I(pwm_setpoint_20));
    InMux I__9739 (
            .O(N__45432),
            .I(N__45429));
    LocalMux I__9738 (
            .O(N__45429),
            .I(n41));
    CascadeMux I__9737 (
            .O(N__45426),
            .I(n41_cascade_));
    InMux I__9736 (
            .O(N__45423),
            .I(N__45420));
    LocalMux I__9735 (
            .O(N__45420),
            .I(N__45417));
    Odrv4 I__9734 (
            .O(N__45417),
            .I(n15265));
    InMux I__9733 (
            .O(N__45414),
            .I(N__45411));
    LocalMux I__9732 (
            .O(N__45411),
            .I(n15112));
    InMux I__9731 (
            .O(N__45408),
            .I(N__45405));
    LocalMux I__9730 (
            .O(N__45405),
            .I(N__45402));
    Span4Mux_h I__9729 (
            .O(N__45402),
            .I(N__45399));
    Odrv4 I__9728 (
            .O(N__45399),
            .I(pwm_setpoint_23));
    InMux I__9727 (
            .O(N__45396),
            .I(N__45393));
    LocalMux I__9726 (
            .O(N__45393),
            .I(n15257));
    InMux I__9725 (
            .O(N__45390),
            .I(N__45387));
    LocalMux I__9724 (
            .O(N__45387),
            .I(N__45384));
    Odrv4 I__9723 (
            .O(N__45384),
            .I(n15108));
    InMux I__9722 (
            .O(N__45381),
            .I(N__45374));
    InMux I__9721 (
            .O(N__45380),
            .I(N__45374));
    InMux I__9720 (
            .O(N__45379),
            .I(N__45371));
    LocalMux I__9719 (
            .O(N__45374),
            .I(pwm_setpoint_21));
    LocalMux I__9718 (
            .O(N__45371),
            .I(pwm_setpoint_21));
    InMux I__9717 (
            .O(N__45366),
            .I(N__45362));
    InMux I__9716 (
            .O(N__45365),
            .I(N__45359));
    LocalMux I__9715 (
            .O(N__45362),
            .I(N__45356));
    LocalMux I__9714 (
            .O(N__45359),
            .I(N__45353));
    Odrv4 I__9713 (
            .O(N__45356),
            .I(pwm_setpoint_19));
    Odrv4 I__9712 (
            .O(N__45353),
            .I(pwm_setpoint_19));
    InMux I__9711 (
            .O(N__45348),
            .I(N__45344));
    InMux I__9710 (
            .O(N__45347),
            .I(N__45341));
    LocalMux I__9709 (
            .O(N__45344),
            .I(N__45338));
    LocalMux I__9708 (
            .O(N__45341),
            .I(n39));
    Odrv4 I__9707 (
            .O(N__45338),
            .I(n39));
    InMux I__9706 (
            .O(N__45333),
            .I(\PWM.n13082 ));
    InMux I__9705 (
            .O(N__45330),
            .I(\PWM.n13083 ));
    InMux I__9704 (
            .O(N__45327),
            .I(\PWM.n13084 ));
    InMux I__9703 (
            .O(N__45324),
            .I(\PWM.n13085 ));
    InMux I__9702 (
            .O(N__45321),
            .I(\PWM.n13086 ));
    CEMux I__9701 (
            .O(N__45318),
            .I(N__45315));
    LocalMux I__9700 (
            .O(N__45315),
            .I(N__45312));
    Span4Mux_h I__9699 (
            .O(N__45312),
            .I(N__45309));
    Odrv4 I__9698 (
            .O(N__45309),
            .I(n6_adj_717));
    InMux I__9697 (
            .O(N__45306),
            .I(N__45303));
    LocalMux I__9696 (
            .O(N__45303),
            .I(N__45299));
    InMux I__9695 (
            .O(N__45302),
            .I(N__45296));
    Span4Mux_h I__9694 (
            .O(N__45299),
            .I(N__45293));
    LocalMux I__9693 (
            .O(N__45296),
            .I(N__45290));
    Odrv4 I__9692 (
            .O(N__45293),
            .I(pwm_setpoint_5));
    Odrv4 I__9691 (
            .O(N__45290),
            .I(pwm_setpoint_5));
    InMux I__9690 (
            .O(N__45285),
            .I(N__45281));
    InMux I__9689 (
            .O(N__45284),
            .I(N__45278));
    LocalMux I__9688 (
            .O(N__45281),
            .I(N__45275));
    LocalMux I__9687 (
            .O(N__45278),
            .I(pwm_setpoint_6));
    Odrv12 I__9686 (
            .O(N__45275),
            .I(pwm_setpoint_6));
    InMux I__9685 (
            .O(N__45270),
            .I(N__45266));
    InMux I__9684 (
            .O(N__45269),
            .I(N__45263));
    LocalMux I__9683 (
            .O(N__45266),
            .I(N__45258));
    LocalMux I__9682 (
            .O(N__45263),
            .I(N__45258));
    Odrv12 I__9681 (
            .O(N__45258),
            .I(pwm_setpoint_10));
    InMux I__9680 (
            .O(N__45255),
            .I(\PWM.n13073 ));
    InMux I__9679 (
            .O(N__45252),
            .I(\PWM.n13074 ));
    InMux I__9678 (
            .O(N__45249),
            .I(\PWM.n13075 ));
    InMux I__9677 (
            .O(N__45246),
            .I(\PWM.n13076 ));
    InMux I__9676 (
            .O(N__45243),
            .I(\PWM.n13077 ));
    InMux I__9675 (
            .O(N__45240),
            .I(\PWM.n13078 ));
    InMux I__9674 (
            .O(N__45237),
            .I(bfn_13_29_0_));
    InMux I__9673 (
            .O(N__45234),
            .I(\PWM.n13080 ));
    InMux I__9672 (
            .O(N__45231),
            .I(\PWM.n13081 ));
    InMux I__9671 (
            .O(N__45228),
            .I(\PWM.n13064 ));
    InMux I__9670 (
            .O(N__45225),
            .I(\PWM.n13065 ));
    InMux I__9669 (
            .O(N__45222),
            .I(\PWM.n13066 ));
    InMux I__9668 (
            .O(N__45219),
            .I(\PWM.n13067 ));
    InMux I__9667 (
            .O(N__45216),
            .I(\PWM.n13068 ));
    InMux I__9666 (
            .O(N__45213),
            .I(\PWM.n13069 ));
    InMux I__9665 (
            .O(N__45210),
            .I(\PWM.n13070 ));
    InMux I__9664 (
            .O(N__45207),
            .I(bfn_13_28_0_));
    InMux I__9663 (
            .O(N__45204),
            .I(\PWM.n13072 ));
    CascadeMux I__9662 (
            .O(N__45201),
            .I(N__45198));
    InMux I__9661 (
            .O(N__45198),
            .I(N__45194));
    InMux I__9660 (
            .O(N__45197),
            .I(N__45191));
    LocalMux I__9659 (
            .O(N__45194),
            .I(N__45188));
    LocalMux I__9658 (
            .O(N__45191),
            .I(pwm_counter_0));
    Odrv12 I__9657 (
            .O(N__45188),
            .I(pwm_counter_0));
    InMux I__9656 (
            .O(N__45183),
            .I(bfn_13_26_0_));
    InMux I__9655 (
            .O(N__45180),
            .I(N__45176));
    InMux I__9654 (
            .O(N__45179),
            .I(N__45173));
    LocalMux I__9653 (
            .O(N__45176),
            .I(N__45170));
    LocalMux I__9652 (
            .O(N__45173),
            .I(pwm_counter_1));
    Odrv12 I__9651 (
            .O(N__45170),
            .I(pwm_counter_1));
    InMux I__9650 (
            .O(N__45165),
            .I(\PWM.n13056 ));
    InMux I__9649 (
            .O(N__45162),
            .I(\PWM.n13057 ));
    InMux I__9648 (
            .O(N__45159),
            .I(\PWM.n13058 ));
    InMux I__9647 (
            .O(N__45156),
            .I(\PWM.n13059 ));
    InMux I__9646 (
            .O(N__45153),
            .I(\PWM.n13060 ));
    InMux I__9645 (
            .O(N__45150),
            .I(\PWM.n13061 ));
    InMux I__9644 (
            .O(N__45147),
            .I(\PWM.n13062 ));
    InMux I__9643 (
            .O(N__45144),
            .I(bfn_13_27_0_));
    CascadeMux I__9642 (
            .O(N__45141),
            .I(N__45137));
    CascadeMux I__9641 (
            .O(N__45140),
            .I(N__45134));
    InMux I__9640 (
            .O(N__45137),
            .I(N__45130));
    InMux I__9639 (
            .O(N__45134),
            .I(N__45125));
    InMux I__9638 (
            .O(N__45133),
            .I(N__45125));
    LocalMux I__9637 (
            .O(N__45130),
            .I(n1029));
    LocalMux I__9636 (
            .O(N__45125),
            .I(n1029));
    InMux I__9635 (
            .O(N__45120),
            .I(N__45117));
    LocalMux I__9634 (
            .O(N__45117),
            .I(n1096));
    InMux I__9633 (
            .O(N__45114),
            .I(n12504));
    CascadeMux I__9632 (
            .O(N__45111),
            .I(N__45108));
    InMux I__9631 (
            .O(N__45108),
            .I(N__45104));
    InMux I__9630 (
            .O(N__45107),
            .I(N__45101));
    LocalMux I__9629 (
            .O(N__45104),
            .I(n1028));
    LocalMux I__9628 (
            .O(N__45101),
            .I(n1028));
    InMux I__9627 (
            .O(N__45096),
            .I(N__45093));
    LocalMux I__9626 (
            .O(N__45093),
            .I(n1095));
    InMux I__9625 (
            .O(N__45090),
            .I(n12505));
    CascadeMux I__9624 (
            .O(N__45087),
            .I(N__45084));
    InMux I__9623 (
            .O(N__45084),
            .I(N__45079));
    InMux I__9622 (
            .O(N__45083),
            .I(N__45074));
    InMux I__9621 (
            .O(N__45082),
            .I(N__45074));
    LocalMux I__9620 (
            .O(N__45079),
            .I(n1027));
    LocalMux I__9619 (
            .O(N__45074),
            .I(n1027));
    InMux I__9618 (
            .O(N__45069),
            .I(N__45066));
    LocalMux I__9617 (
            .O(N__45066),
            .I(n1094));
    InMux I__9616 (
            .O(N__45063),
            .I(n12506));
    InMux I__9615 (
            .O(N__45060),
            .I(bfn_13_24_0_));
    CascadeMux I__9614 (
            .O(N__45057),
            .I(N__45053));
    InMux I__9613 (
            .O(N__45056),
            .I(N__45048));
    InMux I__9612 (
            .O(N__45053),
            .I(N__45048));
    LocalMux I__9611 (
            .O(N__45048),
            .I(N__45044));
    InMux I__9610 (
            .O(N__45047),
            .I(N__45041));
    Odrv4 I__9609 (
            .O(N__45044),
            .I(n1026));
    LocalMux I__9608 (
            .O(N__45041),
            .I(n1026));
    InMux I__9607 (
            .O(N__45036),
            .I(N__45033));
    LocalMux I__9606 (
            .O(N__45033),
            .I(n1093));
    CascadeMux I__9605 (
            .O(N__45030),
            .I(N__45026));
    InMux I__9604 (
            .O(N__45029),
            .I(N__45022));
    InMux I__9603 (
            .O(N__45026),
            .I(N__45019));
    InMux I__9602 (
            .O(N__45025),
            .I(N__45016));
    LocalMux I__9601 (
            .O(N__45022),
            .I(n1030));
    LocalMux I__9600 (
            .O(N__45019),
            .I(n1030));
    LocalMux I__9599 (
            .O(N__45016),
            .I(n1030));
    CascadeMux I__9598 (
            .O(N__45009),
            .I(N__45006));
    InMux I__9597 (
            .O(N__45006),
            .I(N__45003));
    LocalMux I__9596 (
            .O(N__45003),
            .I(n1097));
    CascadeMux I__9595 (
            .O(N__45000),
            .I(n13716_cascade_));
    CascadeMux I__9594 (
            .O(N__44997),
            .I(n1059_cascade_));
    CascadeMux I__9593 (
            .O(N__44994),
            .I(n1126_cascade_));
    InMux I__9592 (
            .O(N__44991),
            .I(N__44988));
    LocalMux I__9591 (
            .O(N__44988),
            .I(N__44984));
    CascadeMux I__9590 (
            .O(N__44987),
            .I(N__44981));
    Span4Mux_v I__9589 (
            .O(N__44984),
            .I(N__44977));
    InMux I__9588 (
            .O(N__44981),
            .I(N__44974));
    InMux I__9587 (
            .O(N__44980),
            .I(N__44971));
    Odrv4 I__9586 (
            .O(N__44977),
            .I(n928));
    LocalMux I__9585 (
            .O(N__44974),
            .I(n928));
    LocalMux I__9584 (
            .O(N__44971),
            .I(n928));
    CascadeMux I__9583 (
            .O(N__44964),
            .I(N__44960));
    CascadeMux I__9582 (
            .O(N__44963),
            .I(N__44957));
    InMux I__9581 (
            .O(N__44960),
            .I(N__44949));
    InMux I__9580 (
            .O(N__44957),
            .I(N__44944));
    InMux I__9579 (
            .O(N__44956),
            .I(N__44944));
    InMux I__9578 (
            .O(N__44955),
            .I(N__44941));
    InMux I__9577 (
            .O(N__44954),
            .I(N__44934));
    InMux I__9576 (
            .O(N__44953),
            .I(N__44934));
    InMux I__9575 (
            .O(N__44952),
            .I(N__44934));
    LocalMux I__9574 (
            .O(N__44949),
            .I(n960));
    LocalMux I__9573 (
            .O(N__44944),
            .I(n960));
    LocalMux I__9572 (
            .O(N__44941),
            .I(n960));
    LocalMux I__9571 (
            .O(N__44934),
            .I(n960));
    InMux I__9570 (
            .O(N__44925),
            .I(N__44922));
    LocalMux I__9569 (
            .O(N__44922),
            .I(n995));
    InMux I__9568 (
            .O(N__44919),
            .I(bfn_13_23_0_));
    InMux I__9567 (
            .O(N__44916),
            .I(n12500));
    InMux I__9566 (
            .O(N__44913),
            .I(n12501));
    InMux I__9565 (
            .O(N__44910),
            .I(n12502));
    InMux I__9564 (
            .O(N__44907),
            .I(n12503));
    InMux I__9563 (
            .O(N__44904),
            .I(N__44901));
    LocalMux I__9562 (
            .O(N__44901),
            .I(N__44898));
    Odrv12 I__9561 (
            .O(N__44898),
            .I(n27));
    InMux I__9560 (
            .O(N__44895),
            .I(N__44892));
    LocalMux I__9559 (
            .O(N__44892),
            .I(N__44888));
    InMux I__9558 (
            .O(N__44891),
            .I(N__44884));
    Span4Mux_h I__9557 (
            .O(N__44888),
            .I(N__44881));
    InMux I__9556 (
            .O(N__44887),
            .I(N__44878));
    LocalMux I__9555 (
            .O(N__44884),
            .I(encoder0_position_6));
    Odrv4 I__9554 (
            .O(N__44881),
            .I(encoder0_position_6));
    LocalMux I__9553 (
            .O(N__44878),
            .I(encoder0_position_6));
    InMux I__9552 (
            .O(N__44871),
            .I(N__44867));
    InMux I__9551 (
            .O(N__44870),
            .I(N__44863));
    LocalMux I__9550 (
            .O(N__44867),
            .I(N__44860));
    InMux I__9549 (
            .O(N__44866),
            .I(N__44857));
    LocalMux I__9548 (
            .O(N__44863),
            .I(N__44854));
    Span4Mux_v I__9547 (
            .O(N__44860),
            .I(N__44851));
    LocalMux I__9546 (
            .O(N__44857),
            .I(N__44848));
    Span4Mux_v I__9545 (
            .O(N__44854),
            .I(N__44845));
    Span4Mux_h I__9544 (
            .O(N__44851),
            .I(N__44842));
    Span12Mux_s8_v I__9543 (
            .O(N__44848),
            .I(N__44839));
    Span4Mux_h I__9542 (
            .O(N__44845),
            .I(N__44836));
    Span4Mux_h I__9541 (
            .O(N__44842),
            .I(N__44833));
    Span12Mux_h I__9540 (
            .O(N__44839),
            .I(N__44830));
    Span4Mux_h I__9539 (
            .O(N__44836),
            .I(N__44827));
    Span4Mux_h I__9538 (
            .O(N__44833),
            .I(N__44824));
    Odrv12 I__9537 (
            .O(N__44830),
            .I(n313));
    Odrv4 I__9536 (
            .O(N__44827),
            .I(n313));
    Odrv4 I__9535 (
            .O(N__44824),
            .I(n313));
    InMux I__9534 (
            .O(N__44817),
            .I(N__44814));
    LocalMux I__9533 (
            .O(N__44814),
            .I(N__44811));
    Span4Mux_h I__9532 (
            .O(N__44811),
            .I(N__44808));
    Odrv4 I__9531 (
            .O(N__44808),
            .I(n11));
    InMux I__9530 (
            .O(N__44805),
            .I(N__44799));
    InMux I__9529 (
            .O(N__44804),
            .I(N__44799));
    LocalMux I__9528 (
            .O(N__44799),
            .I(N__44795));
    InMux I__9527 (
            .O(N__44798),
            .I(N__44792));
    Span4Mux_h I__9526 (
            .O(N__44795),
            .I(N__44789));
    LocalMux I__9525 (
            .O(N__44792),
            .I(encoder0_position_22));
    Odrv4 I__9524 (
            .O(N__44789),
            .I(encoder0_position_22));
    CascadeMux I__9523 (
            .O(N__44784),
            .I(N__44781));
    InMux I__9522 (
            .O(N__44781),
            .I(N__44778));
    LocalMux I__9521 (
            .O(N__44778),
            .I(N__44775));
    Span4Mux_h I__9520 (
            .O(N__44775),
            .I(N__44772));
    Odrv4 I__9519 (
            .O(N__44772),
            .I(n11_adj_632));
    InMux I__9518 (
            .O(N__44769),
            .I(N__44766));
    LocalMux I__9517 (
            .O(N__44766),
            .I(N__44763));
    Span4Mux_h I__9516 (
            .O(N__44763),
            .I(N__44760));
    Odrv4 I__9515 (
            .O(N__44760),
            .I(n9));
    InMux I__9514 (
            .O(N__44757),
            .I(N__44753));
    InMux I__9513 (
            .O(N__44756),
            .I(N__44750));
    LocalMux I__9512 (
            .O(N__44753),
            .I(N__44745));
    LocalMux I__9511 (
            .O(N__44750),
            .I(N__44745));
    Span4Mux_v I__9510 (
            .O(N__44745),
            .I(N__44741));
    InMux I__9509 (
            .O(N__44744),
            .I(N__44738));
    Sp12to4 I__9508 (
            .O(N__44741),
            .I(N__44735));
    LocalMux I__9507 (
            .O(N__44738),
            .I(n295));
    Odrv12 I__9506 (
            .O(N__44735),
            .I(n295));
    InMux I__9505 (
            .O(N__44730),
            .I(N__44723));
    InMux I__9504 (
            .O(N__44729),
            .I(N__44723));
    CascadeMux I__9503 (
            .O(N__44728),
            .I(N__44720));
    LocalMux I__9502 (
            .O(N__44723),
            .I(N__44717));
    InMux I__9501 (
            .O(N__44720),
            .I(N__44714));
    Span4Mux_h I__9500 (
            .O(N__44717),
            .I(N__44711));
    LocalMux I__9499 (
            .O(N__44714),
            .I(encoder0_position_24));
    Odrv4 I__9498 (
            .O(N__44711),
            .I(encoder0_position_24));
    CascadeMux I__9497 (
            .O(N__44706),
            .I(N__44703));
    InMux I__9496 (
            .O(N__44703),
            .I(N__44700));
    LocalMux I__9495 (
            .O(N__44700),
            .I(N__44697));
    Span4Mux_h I__9494 (
            .O(N__44697),
            .I(N__44694));
    Odrv4 I__9493 (
            .O(N__44694),
            .I(n9_adj_630));
    InMux I__9492 (
            .O(N__44691),
            .I(N__44688));
    LocalMux I__9491 (
            .O(N__44688),
            .I(N__44684));
    CascadeMux I__9490 (
            .O(N__44687),
            .I(N__44681));
    Span4Mux_v I__9489 (
            .O(N__44684),
            .I(N__44677));
    InMux I__9488 (
            .O(N__44681),
            .I(N__44674));
    InMux I__9487 (
            .O(N__44680),
            .I(N__44671));
    Odrv4 I__9486 (
            .O(N__44677),
            .I(n933));
    LocalMux I__9485 (
            .O(N__44674),
            .I(n933));
    LocalMux I__9484 (
            .O(N__44671),
            .I(n933));
    CascadeMux I__9483 (
            .O(N__44664),
            .I(N__44661));
    InMux I__9482 (
            .O(N__44661),
            .I(N__44658));
    LocalMux I__9481 (
            .O(N__44658),
            .I(n1000));
    CascadeMux I__9480 (
            .O(N__44655),
            .I(n1032_cascade_));
    CascadeMux I__9479 (
            .O(N__44652),
            .I(n11914_cascade_));
    InMux I__9478 (
            .O(N__44649),
            .I(n12556));
    InMux I__9477 (
            .O(N__44646),
            .I(bfn_13_20_0_));
    InMux I__9476 (
            .O(N__44643),
            .I(n12558));
    InMux I__9475 (
            .O(N__44640),
            .I(N__44637));
    LocalMux I__9474 (
            .O(N__44637),
            .I(n1591));
    InMux I__9473 (
            .O(N__44634),
            .I(n12559));
    InMux I__9472 (
            .O(N__44631),
            .I(n12560));
    InMux I__9471 (
            .O(N__44628),
            .I(n12561));
    InMux I__9470 (
            .O(N__44625),
            .I(n12562));
    InMux I__9469 (
            .O(N__44622),
            .I(N__44619));
    LocalMux I__9468 (
            .O(N__44619),
            .I(N__44616));
    Span4Mux_h I__9467 (
            .O(N__44616),
            .I(N__44613));
    Odrv4 I__9466 (
            .O(N__44613),
            .I(n13));
    InMux I__9465 (
            .O(N__44610),
            .I(N__44607));
    LocalMux I__9464 (
            .O(N__44607),
            .I(N__44602));
    InMux I__9463 (
            .O(N__44606),
            .I(N__44599));
    InMux I__9462 (
            .O(N__44605),
            .I(N__44596));
    Span4Mux_v I__9461 (
            .O(N__44602),
            .I(N__44593));
    LocalMux I__9460 (
            .O(N__44599),
            .I(N__44590));
    LocalMux I__9459 (
            .O(N__44596),
            .I(encoder0_position_20));
    Odrv4 I__9458 (
            .O(N__44593),
            .I(encoder0_position_20));
    Odrv4 I__9457 (
            .O(N__44590),
            .I(encoder0_position_20));
    CascadeMux I__9456 (
            .O(N__44583),
            .I(N__44580));
    InMux I__9455 (
            .O(N__44580),
            .I(N__44575));
    InMux I__9454 (
            .O(N__44579),
            .I(N__44572));
    InMux I__9453 (
            .O(N__44578),
            .I(N__44569));
    LocalMux I__9452 (
            .O(N__44575),
            .I(n1720));
    LocalMux I__9451 (
            .O(N__44572),
            .I(n1720));
    LocalMux I__9450 (
            .O(N__44569),
            .I(n1720));
    InMux I__9449 (
            .O(N__44562),
            .I(N__44559));
    LocalMux I__9448 (
            .O(N__44559),
            .I(N__44556));
    Odrv4 I__9447 (
            .O(N__44556),
            .I(n1787));
    InMux I__9446 (
            .O(N__44553),
            .I(n12590));
    InMux I__9445 (
            .O(N__44550),
            .I(N__44547));
    LocalMux I__9444 (
            .O(N__44547),
            .I(N__44544));
    Span4Mux_v I__9443 (
            .O(N__44544),
            .I(N__44540));
    InMux I__9442 (
            .O(N__44543),
            .I(N__44537));
    Span4Mux_h I__9441 (
            .O(N__44540),
            .I(N__44534));
    LocalMux I__9440 (
            .O(N__44537),
            .I(N__44531));
    Odrv4 I__9439 (
            .O(N__44534),
            .I(n15622));
    Odrv4 I__9438 (
            .O(N__44531),
            .I(n15622));
    InMux I__9437 (
            .O(N__44526),
            .I(n12591));
    InMux I__9436 (
            .O(N__44523),
            .I(N__44520));
    LocalMux I__9435 (
            .O(N__44520),
            .I(N__44515));
    InMux I__9434 (
            .O(N__44519),
            .I(N__44512));
    InMux I__9433 (
            .O(N__44518),
            .I(N__44509));
    Span4Mux_v I__9432 (
            .O(N__44515),
            .I(N__44504));
    LocalMux I__9431 (
            .O(N__44512),
            .I(N__44504));
    LocalMux I__9430 (
            .O(N__44509),
            .I(n1818));
    Odrv4 I__9429 (
            .O(N__44504),
            .I(n1818));
    InMux I__9428 (
            .O(N__44499),
            .I(bfn_13_19_0_));
    InMux I__9427 (
            .O(N__44496),
            .I(n12550));
    InMux I__9426 (
            .O(N__44493),
            .I(n12551));
    InMux I__9425 (
            .O(N__44490),
            .I(n12552));
    InMux I__9424 (
            .O(N__44487),
            .I(n12553));
    InMux I__9423 (
            .O(N__44484),
            .I(n12554));
    InMux I__9422 (
            .O(N__44481),
            .I(n12555));
    InMux I__9421 (
            .O(N__44478),
            .I(N__44475));
    LocalMux I__9420 (
            .O(N__44475),
            .I(N__44472));
    Odrv4 I__9419 (
            .O(N__44472),
            .I(n1795));
    InMux I__9418 (
            .O(N__44469),
            .I(n12582));
    CascadeMux I__9417 (
            .O(N__44466),
            .I(N__44463));
    InMux I__9416 (
            .O(N__44463),
            .I(N__44460));
    LocalMux I__9415 (
            .O(N__44460),
            .I(N__44457));
    Odrv4 I__9414 (
            .O(N__44457),
            .I(n1794));
    InMux I__9413 (
            .O(N__44454),
            .I(n12583));
    InMux I__9412 (
            .O(N__44451),
            .I(N__44448));
    LocalMux I__9411 (
            .O(N__44448),
            .I(N__44445));
    Odrv4 I__9410 (
            .O(N__44445),
            .I(n1793));
    InMux I__9409 (
            .O(N__44442),
            .I(bfn_13_18_0_));
    CascadeMux I__9408 (
            .O(N__44439),
            .I(N__44436));
    InMux I__9407 (
            .O(N__44436),
            .I(N__44433));
    LocalMux I__9406 (
            .O(N__44433),
            .I(N__44430));
    Odrv4 I__9405 (
            .O(N__44430),
            .I(n1792));
    InMux I__9404 (
            .O(N__44427),
            .I(n12585));
    InMux I__9403 (
            .O(N__44424),
            .I(N__44421));
    LocalMux I__9402 (
            .O(N__44421),
            .I(N__44418));
    Odrv4 I__9401 (
            .O(N__44418),
            .I(n1791));
    InMux I__9400 (
            .O(N__44415),
            .I(n12586));
    InMux I__9399 (
            .O(N__44412),
            .I(N__44409));
    LocalMux I__9398 (
            .O(N__44409),
            .I(N__44406));
    Span4Mux_v I__9397 (
            .O(N__44406),
            .I(N__44403));
    Odrv4 I__9396 (
            .O(N__44403),
            .I(n1790));
    InMux I__9395 (
            .O(N__44400),
            .I(n12587));
    CascadeMux I__9394 (
            .O(N__44397),
            .I(N__44394));
    InMux I__9393 (
            .O(N__44394),
            .I(N__44390));
    InMux I__9392 (
            .O(N__44393),
            .I(N__44387));
    LocalMux I__9391 (
            .O(N__44390),
            .I(n1722));
    LocalMux I__9390 (
            .O(N__44387),
            .I(n1722));
    InMux I__9389 (
            .O(N__44382),
            .I(N__44379));
    LocalMux I__9388 (
            .O(N__44379),
            .I(n1789));
    InMux I__9387 (
            .O(N__44376),
            .I(n12588));
    InMux I__9386 (
            .O(N__44373),
            .I(N__44368));
    InMux I__9385 (
            .O(N__44372),
            .I(N__44365));
    InMux I__9384 (
            .O(N__44371),
            .I(N__44362));
    LocalMux I__9383 (
            .O(N__44368),
            .I(n1721));
    LocalMux I__9382 (
            .O(N__44365),
            .I(n1721));
    LocalMux I__9381 (
            .O(N__44362),
            .I(n1721));
    InMux I__9380 (
            .O(N__44355),
            .I(N__44352));
    LocalMux I__9379 (
            .O(N__44352),
            .I(N__44349));
    Span4Mux_h I__9378 (
            .O(N__44349),
            .I(N__44346));
    Odrv4 I__9377 (
            .O(N__44346),
            .I(n1788));
    InMux I__9376 (
            .O(N__44343),
            .I(n12589));
    SRMux I__9375 (
            .O(N__44340),
            .I(N__44336));
    InMux I__9374 (
            .O(N__44339),
            .I(N__44333));
    LocalMux I__9373 (
            .O(N__44336),
            .I(N__44330));
    LocalMux I__9372 (
            .O(N__44333),
            .I(N__44327));
    Odrv12 I__9371 (
            .O(N__44330),
            .I(pwm_setpoint_23__N_195));
    Odrv4 I__9370 (
            .O(N__44327),
            .I(pwm_setpoint_23__N_195));
    InMux I__9369 (
            .O(N__44322),
            .I(N__44319));
    LocalMux I__9368 (
            .O(N__44319),
            .I(N__44316));
    Odrv12 I__9367 (
            .O(N__44316),
            .I(pwm_setpoint_23_N_171_21));
    InMux I__9366 (
            .O(N__44313),
            .I(N__44307));
    InMux I__9365 (
            .O(N__44312),
            .I(N__44307));
    LocalMux I__9364 (
            .O(N__44307),
            .I(N__44304));
    Odrv12 I__9363 (
            .O(N__44304),
            .I(duty_21));
    InMux I__9362 (
            .O(N__44301),
            .I(N__44298));
    LocalMux I__9361 (
            .O(N__44298),
            .I(N__44295));
    Span4Mux_v I__9360 (
            .O(N__44295),
            .I(N__44292));
    Span4Mux_h I__9359 (
            .O(N__44292),
            .I(N__44289));
    Odrv4 I__9358 (
            .O(N__44289),
            .I(n1801));
    InMux I__9357 (
            .O(N__44286),
            .I(bfn_13_17_0_));
    CascadeMux I__9356 (
            .O(N__44283),
            .I(N__44280));
    InMux I__9355 (
            .O(N__44280),
            .I(N__44277));
    LocalMux I__9354 (
            .O(N__44277),
            .I(N__44274));
    Span4Mux_v I__9353 (
            .O(N__44274),
            .I(N__44271));
    Odrv4 I__9352 (
            .O(N__44271),
            .I(n1800));
    InMux I__9351 (
            .O(N__44268),
            .I(n12577));
    InMux I__9350 (
            .O(N__44265),
            .I(N__44262));
    LocalMux I__9349 (
            .O(N__44262),
            .I(N__44259));
    Span4Mux_v I__9348 (
            .O(N__44259),
            .I(N__44256));
    Odrv4 I__9347 (
            .O(N__44256),
            .I(n1799));
    InMux I__9346 (
            .O(N__44253),
            .I(n12578));
    InMux I__9345 (
            .O(N__44250),
            .I(N__44247));
    LocalMux I__9344 (
            .O(N__44247),
            .I(N__44244));
    Odrv4 I__9343 (
            .O(N__44244),
            .I(n1798));
    InMux I__9342 (
            .O(N__44241),
            .I(n12579));
    InMux I__9341 (
            .O(N__44238),
            .I(N__44235));
    LocalMux I__9340 (
            .O(N__44235),
            .I(N__44232));
    Odrv4 I__9339 (
            .O(N__44232),
            .I(n1797));
    InMux I__9338 (
            .O(N__44229),
            .I(n12580));
    CascadeMux I__9337 (
            .O(N__44226),
            .I(N__44223));
    InMux I__9336 (
            .O(N__44223),
            .I(N__44220));
    LocalMux I__9335 (
            .O(N__44220),
            .I(N__44217));
    Span4Mux_v I__9334 (
            .O(N__44217),
            .I(N__44214));
    Odrv4 I__9333 (
            .O(N__44214),
            .I(n1796));
    InMux I__9332 (
            .O(N__44211),
            .I(n12581));
    CascadeMux I__9331 (
            .O(N__44208),
            .I(n8_adj_657_cascade_));
    InMux I__9330 (
            .O(N__44205),
            .I(N__44202));
    LocalMux I__9329 (
            .O(N__44202),
            .I(N__44199));
    Odrv12 I__9328 (
            .O(N__44199),
            .I(n15180));
    CascadeMux I__9327 (
            .O(N__44196),
            .I(n15219_cascade_));
    InMux I__9326 (
            .O(N__44193),
            .I(N__44190));
    LocalMux I__9325 (
            .O(N__44190),
            .I(n24_adj_669));
    InMux I__9324 (
            .O(N__44187),
            .I(N__44181));
    InMux I__9323 (
            .O(N__44186),
            .I(N__44181));
    LocalMux I__9322 (
            .O(N__44181),
            .I(N__44178));
    Span4Mux_h I__9321 (
            .O(N__44178),
            .I(N__44175));
    Odrv4 I__9320 (
            .O(N__44175),
            .I(pwm_setpoint_22));
    InMux I__9319 (
            .O(N__44172),
            .I(N__44169));
    LocalMux I__9318 (
            .O(N__44169),
            .I(n15274));
    InMux I__9317 (
            .O(N__44166),
            .I(N__44160));
    InMux I__9316 (
            .O(N__44165),
            .I(N__44153));
    InMux I__9315 (
            .O(N__44164),
            .I(N__44153));
    InMux I__9314 (
            .O(N__44163),
            .I(N__44153));
    LocalMux I__9313 (
            .O(N__44160),
            .I(n45));
    LocalMux I__9312 (
            .O(N__44153),
            .I(n45));
    InMux I__9311 (
            .O(N__44148),
            .I(N__44145));
    LocalMux I__9310 (
            .O(N__44145),
            .I(n15255));
    CascadeMux I__9309 (
            .O(N__44142),
            .I(n40_cascade_));
    InMux I__9308 (
            .O(N__44139),
            .I(N__44135));
    InMux I__9307 (
            .O(N__44138),
            .I(N__44132));
    LocalMux I__9306 (
            .O(N__44135),
            .I(N__44127));
    LocalMux I__9305 (
            .O(N__44132),
            .I(N__44127));
    Span4Mux_s2_v I__9304 (
            .O(N__44127),
            .I(N__44124));
    Odrv4 I__9303 (
            .O(N__44124),
            .I(duty_20));
    InMux I__9302 (
            .O(N__44121),
            .I(N__44118));
    LocalMux I__9301 (
            .O(N__44118),
            .I(N__44115));
    Odrv4 I__9300 (
            .O(N__44115),
            .I(pwm_setpoint_23_N_171_20));
    CascadeMux I__9299 (
            .O(N__44112),
            .I(N__44109));
    InMux I__9298 (
            .O(N__44109),
            .I(N__44106));
    LocalMux I__9297 (
            .O(N__44106),
            .I(N__44103));
    Odrv12 I__9296 (
            .O(N__44103),
            .I(n4_adj_584));
    InMux I__9295 (
            .O(N__44100),
            .I(N__44097));
    LocalMux I__9294 (
            .O(N__44097),
            .I(n16_adj_664));
    InMux I__9293 (
            .O(N__44094),
            .I(N__44090));
    InMux I__9292 (
            .O(N__44093),
            .I(N__44087));
    LocalMux I__9291 (
            .O(N__44090),
            .I(N__44084));
    LocalMux I__9290 (
            .O(N__44087),
            .I(N__44079));
    Span4Mux_h I__9289 (
            .O(N__44084),
            .I(N__44079));
    Odrv4 I__9288 (
            .O(N__44079),
            .I(duty_12));
    InMux I__9287 (
            .O(N__44076),
            .I(N__44073));
    LocalMux I__9286 (
            .O(N__44073),
            .I(N__44070));
    Span4Mux_h I__9285 (
            .O(N__44070),
            .I(N__44067));
    Odrv4 I__9284 (
            .O(N__44067),
            .I(pwm_setpoint_23_N_171_12));
    InMux I__9283 (
            .O(N__44064),
            .I(N__44058));
    InMux I__9282 (
            .O(N__44063),
            .I(N__44058));
    LocalMux I__9281 (
            .O(N__44058),
            .I(n37));
    InMux I__9280 (
            .O(N__44055),
            .I(N__44051));
    InMux I__9279 (
            .O(N__44054),
            .I(N__44048));
    LocalMux I__9278 (
            .O(N__44051),
            .I(N__44045));
    LocalMux I__9277 (
            .O(N__44048),
            .I(N__44042));
    Span4Mux_h I__9276 (
            .O(N__44045),
            .I(N__44039));
    Span4Mux_h I__9275 (
            .O(N__44042),
            .I(N__44036));
    Odrv4 I__9274 (
            .O(N__44039),
            .I(pwm_setpoint_18));
    Odrv4 I__9273 (
            .O(N__44036),
            .I(pwm_setpoint_18));
    InMux I__9272 (
            .O(N__44031),
            .I(N__44028));
    LocalMux I__9271 (
            .O(N__44028),
            .I(N__44025));
    Odrv4 I__9270 (
            .O(N__44025),
            .I(n15277));
    InMux I__9269 (
            .O(N__44022),
            .I(N__44019));
    LocalMux I__9268 (
            .O(N__44019),
            .I(N__44016));
    Odrv4 I__9267 (
            .O(N__44016),
            .I(n6_adj_656));
    CascadeMux I__9266 (
            .O(N__44013),
            .I(n15235_cascade_));
    CascadeMux I__9265 (
            .O(N__44010),
            .I(n15236_cascade_));
    InMux I__9264 (
            .O(N__44007),
            .I(N__44003));
    InMux I__9263 (
            .O(N__44006),
            .I(N__44000));
    LocalMux I__9262 (
            .O(N__44003),
            .I(N__43997));
    LocalMux I__9261 (
            .O(N__44000),
            .I(N__43994));
    Span4Mux_v I__9260 (
            .O(N__43997),
            .I(N__43991));
    Odrv4 I__9259 (
            .O(N__43994),
            .I(duty_11));
    Odrv4 I__9258 (
            .O(N__43991),
            .I(duty_11));
    InMux I__9257 (
            .O(N__43986),
            .I(N__43983));
    LocalMux I__9256 (
            .O(N__43983),
            .I(N__43980));
    Span4Mux_v I__9255 (
            .O(N__43980),
            .I(N__43977));
    Odrv4 I__9254 (
            .O(N__43977),
            .I(pwm_setpoint_23_N_171_11));
    InMux I__9253 (
            .O(N__43974),
            .I(N__43970));
    InMux I__9252 (
            .O(N__43973),
            .I(N__43967));
    LocalMux I__9251 (
            .O(N__43970),
            .I(N__43964));
    LocalMux I__9250 (
            .O(N__43967),
            .I(N__43961));
    Span4Mux_s2_v I__9249 (
            .O(N__43964),
            .I(N__43958));
    Odrv4 I__9248 (
            .O(N__43961),
            .I(duty_17));
    Odrv4 I__9247 (
            .O(N__43958),
            .I(duty_17));
    InMux I__9246 (
            .O(N__43953),
            .I(N__43950));
    LocalMux I__9245 (
            .O(N__43950),
            .I(N__43947));
    Span4Mux_h I__9244 (
            .O(N__43947),
            .I(N__43944));
    Odrv4 I__9243 (
            .O(N__43944),
            .I(pwm_setpoint_23_N_171_17));
    InMux I__9242 (
            .O(N__43941),
            .I(N__43938));
    LocalMux I__9241 (
            .O(N__43938),
            .I(N__43935));
    Span4Mux_h I__9240 (
            .O(N__43935),
            .I(N__43931));
    InMux I__9239 (
            .O(N__43934),
            .I(N__43928));
    Odrv4 I__9238 (
            .O(N__43931),
            .I(pwm_setpoint_17));
    LocalMux I__9237 (
            .O(N__43928),
            .I(pwm_setpoint_17));
    InMux I__9236 (
            .O(N__43923),
            .I(N__43920));
    LocalMux I__9235 (
            .O(N__43920),
            .I(n15278));
    InMux I__9234 (
            .O(N__43917),
            .I(N__43914));
    LocalMux I__9233 (
            .O(N__43914),
            .I(N__43911));
    Odrv12 I__9232 (
            .O(N__43911),
            .I(n6_adj_577));
    InMux I__9231 (
            .O(N__43908),
            .I(N__43904));
    InMux I__9230 (
            .O(N__43907),
            .I(N__43901));
    LocalMux I__9229 (
            .O(N__43904),
            .I(N__43898));
    LocalMux I__9228 (
            .O(N__43901),
            .I(N__43895));
    Span4Mux_s3_v I__9227 (
            .O(N__43898),
            .I(N__43890));
    Span4Mux_h I__9226 (
            .O(N__43895),
            .I(N__43890));
    Odrv4 I__9225 (
            .O(N__43890),
            .I(duty_19));
    InMux I__9224 (
            .O(N__43887),
            .I(n12477));
    CascadeMux I__9223 (
            .O(N__43884),
            .I(N__43881));
    InMux I__9222 (
            .O(N__43881),
            .I(N__43878));
    LocalMux I__9221 (
            .O(N__43878),
            .I(n5_adj_578));
    InMux I__9220 (
            .O(N__43875),
            .I(n12478));
    InMux I__9219 (
            .O(N__43872),
            .I(N__43869));
    LocalMux I__9218 (
            .O(N__43869),
            .I(N__43866));
    Odrv12 I__9217 (
            .O(N__43866),
            .I(n4_adj_579));
    InMux I__9216 (
            .O(N__43863),
            .I(n12479));
    InMux I__9215 (
            .O(N__43860),
            .I(N__43857));
    LocalMux I__9214 (
            .O(N__43857),
            .I(N__43854));
    Span4Mux_v I__9213 (
            .O(N__43854),
            .I(N__43851));
    Odrv4 I__9212 (
            .O(N__43851),
            .I(n3_adj_580));
    InMux I__9211 (
            .O(N__43848),
            .I(N__43842));
    InMux I__9210 (
            .O(N__43847),
            .I(N__43842));
    LocalMux I__9209 (
            .O(N__43842),
            .I(N__43839));
    Span12Mux_s4_v I__9208 (
            .O(N__43839),
            .I(N__43836));
    Odrv12 I__9207 (
            .O(N__43836),
            .I(duty_22));
    InMux I__9206 (
            .O(N__43833),
            .I(n12480));
    InMux I__9205 (
            .O(N__43830),
            .I(N__43827));
    LocalMux I__9204 (
            .O(N__43827),
            .I(n2_adj_581));
    InMux I__9203 (
            .O(N__43824),
            .I(n12481));
    InMux I__9202 (
            .O(N__43821),
            .I(N__43812));
    InMux I__9201 (
            .O(N__43820),
            .I(N__43812));
    InMux I__9200 (
            .O(N__43819),
            .I(N__43812));
    LocalMux I__9199 (
            .O(N__43812),
            .I(N__43809));
    Odrv4 I__9198 (
            .O(N__43809),
            .I(n35));
    InMux I__9197 (
            .O(N__43806),
            .I(N__43803));
    LocalMux I__9196 (
            .O(N__43803),
            .I(N__43800));
    Span4Mux_h I__9195 (
            .O(N__43800),
            .I(N__43797));
    Odrv4 I__9194 (
            .O(N__43797),
            .I(n33_adj_675));
    CascadeMux I__9193 (
            .O(N__43794),
            .I(n35_cascade_));
    InMux I__9192 (
            .O(N__43791),
            .I(N__43788));
    LocalMux I__9191 (
            .O(N__43788),
            .I(N__43785));
    Odrv12 I__9190 (
            .O(N__43785),
            .I(n15225));
    InMux I__9189 (
            .O(N__43782),
            .I(N__43778));
    InMux I__9188 (
            .O(N__43781),
            .I(N__43775));
    LocalMux I__9187 (
            .O(N__43778),
            .I(N__43772));
    LocalMux I__9186 (
            .O(N__43775),
            .I(pwm_setpoint_13));
    Odrv4 I__9185 (
            .O(N__43772),
            .I(pwm_setpoint_13));
    CascadeMux I__9184 (
            .O(N__43767),
            .I(N__43764));
    InMux I__9183 (
            .O(N__43764),
            .I(N__43759));
    InMux I__9182 (
            .O(N__43763),
            .I(N__43756));
    InMux I__9181 (
            .O(N__43762),
            .I(N__43753));
    LocalMux I__9180 (
            .O(N__43759),
            .I(N__43750));
    LocalMux I__9179 (
            .O(N__43756),
            .I(N__43745));
    LocalMux I__9178 (
            .O(N__43753),
            .I(N__43745));
    Sp12to4 I__9177 (
            .O(N__43750),
            .I(N__43742));
    Span4Mux_h I__9176 (
            .O(N__43745),
            .I(N__43739));
    Odrv12 I__9175 (
            .O(N__43742),
            .I(n27_adj_671));
    Odrv4 I__9174 (
            .O(N__43739),
            .I(n27_adj_671));
    InMux I__9173 (
            .O(N__43734),
            .I(N__43731));
    LocalMux I__9172 (
            .O(N__43731),
            .I(n14_adj_569));
    InMux I__9171 (
            .O(N__43728),
            .I(n12469));
    InMux I__9170 (
            .O(N__43725),
            .I(N__43722));
    LocalMux I__9169 (
            .O(N__43722),
            .I(N__43719));
    Odrv12 I__9168 (
            .O(N__43719),
            .I(n13_adj_570));
    InMux I__9167 (
            .O(N__43716),
            .I(n12470));
    InMux I__9166 (
            .O(N__43713),
            .I(N__43710));
    LocalMux I__9165 (
            .O(N__43710),
            .I(N__43707));
    Span4Mux_v I__9164 (
            .O(N__43707),
            .I(N__43704));
    Odrv4 I__9163 (
            .O(N__43704),
            .I(n12_adj_571));
    InMux I__9162 (
            .O(N__43701),
            .I(N__43698));
    LocalMux I__9161 (
            .O(N__43698),
            .I(N__43694));
    InMux I__9160 (
            .O(N__43697),
            .I(N__43691));
    Span4Mux_v I__9159 (
            .O(N__43694),
            .I(N__43688));
    LocalMux I__9158 (
            .O(N__43691),
            .I(duty_13));
    Odrv4 I__9157 (
            .O(N__43688),
            .I(duty_13));
    InMux I__9156 (
            .O(N__43683),
            .I(n12471));
    InMux I__9155 (
            .O(N__43680),
            .I(N__43677));
    LocalMux I__9154 (
            .O(N__43677),
            .I(n11_adj_572));
    InMux I__9153 (
            .O(N__43674),
            .I(N__43670));
    InMux I__9152 (
            .O(N__43673),
            .I(N__43667));
    LocalMux I__9151 (
            .O(N__43670),
            .I(N__43662));
    LocalMux I__9150 (
            .O(N__43667),
            .I(N__43662));
    Span4Mux_v I__9149 (
            .O(N__43662),
            .I(N__43659));
    Odrv4 I__9148 (
            .O(N__43659),
            .I(duty_14));
    InMux I__9147 (
            .O(N__43656),
            .I(n12472));
    CascadeMux I__9146 (
            .O(N__43653),
            .I(N__43650));
    InMux I__9145 (
            .O(N__43650),
            .I(N__43647));
    LocalMux I__9144 (
            .O(N__43647),
            .I(N__43644));
    Span4Mux_v I__9143 (
            .O(N__43644),
            .I(N__43641));
    Sp12to4 I__9142 (
            .O(N__43641),
            .I(N__43638));
    Odrv12 I__9141 (
            .O(N__43638),
            .I(n10_adj_573));
    InMux I__9140 (
            .O(N__43635),
            .I(N__43631));
    InMux I__9139 (
            .O(N__43634),
            .I(N__43628));
    LocalMux I__9138 (
            .O(N__43631),
            .I(N__43625));
    LocalMux I__9137 (
            .O(N__43628),
            .I(N__43622));
    Span4Mux_v I__9136 (
            .O(N__43625),
            .I(N__43619));
    Span4Mux_h I__9135 (
            .O(N__43622),
            .I(N__43616));
    Odrv4 I__9134 (
            .O(N__43619),
            .I(duty_15));
    Odrv4 I__9133 (
            .O(N__43616),
            .I(duty_15));
    InMux I__9132 (
            .O(N__43611),
            .I(n12473));
    InMux I__9131 (
            .O(N__43608),
            .I(N__43605));
    LocalMux I__9130 (
            .O(N__43605),
            .I(N__43602));
    Odrv4 I__9129 (
            .O(N__43602),
            .I(n9_adj_574));
    InMux I__9128 (
            .O(N__43599),
            .I(N__43595));
    InMux I__9127 (
            .O(N__43598),
            .I(N__43592));
    LocalMux I__9126 (
            .O(N__43595),
            .I(N__43589));
    LocalMux I__9125 (
            .O(N__43592),
            .I(N__43586));
    Span4Mux_h I__9124 (
            .O(N__43589),
            .I(N__43581));
    Span4Mux_v I__9123 (
            .O(N__43586),
            .I(N__43581));
    Odrv4 I__9122 (
            .O(N__43581),
            .I(duty_16));
    InMux I__9121 (
            .O(N__43578),
            .I(bfn_12_28_0_));
    InMux I__9120 (
            .O(N__43575),
            .I(N__43572));
    LocalMux I__9119 (
            .O(N__43572),
            .I(N__43569));
    Span4Mux_h I__9118 (
            .O(N__43569),
            .I(N__43566));
    Odrv4 I__9117 (
            .O(N__43566),
            .I(n8_adj_575));
    InMux I__9116 (
            .O(N__43563),
            .I(n12475));
    InMux I__9115 (
            .O(N__43560),
            .I(N__43557));
    LocalMux I__9114 (
            .O(N__43557),
            .I(n7_adj_576));
    InMux I__9113 (
            .O(N__43554),
            .I(N__43550));
    InMux I__9112 (
            .O(N__43553),
            .I(N__43547));
    LocalMux I__9111 (
            .O(N__43550),
            .I(N__43544));
    LocalMux I__9110 (
            .O(N__43547),
            .I(N__43541));
    Span4Mux_v I__9109 (
            .O(N__43544),
            .I(N__43538));
    Span4Mux_h I__9108 (
            .O(N__43541),
            .I(N__43535));
    Odrv4 I__9107 (
            .O(N__43538),
            .I(duty_18));
    Odrv4 I__9106 (
            .O(N__43535),
            .I(duty_18));
    InMux I__9105 (
            .O(N__43530),
            .I(n12476));
    InMux I__9104 (
            .O(N__43527),
            .I(N__43524));
    LocalMux I__9103 (
            .O(N__43524),
            .I(N__43521));
    Odrv4 I__9102 (
            .O(N__43521),
            .I(n22_adj_555));
    InMux I__9101 (
            .O(N__43518),
            .I(N__43515));
    LocalMux I__9100 (
            .O(N__43515),
            .I(N__43511));
    InMux I__9099 (
            .O(N__43514),
            .I(N__43508));
    Span4Mux_h I__9098 (
            .O(N__43511),
            .I(N__43505));
    LocalMux I__9097 (
            .O(N__43508),
            .I(duty_3));
    Odrv4 I__9096 (
            .O(N__43505),
            .I(duty_3));
    InMux I__9095 (
            .O(N__43500),
            .I(n12461));
    CascadeMux I__9094 (
            .O(N__43497),
            .I(N__43494));
    InMux I__9093 (
            .O(N__43494),
            .I(N__43491));
    LocalMux I__9092 (
            .O(N__43491),
            .I(N__43488));
    Odrv4 I__9091 (
            .O(N__43488),
            .I(n21_adj_556));
    InMux I__9090 (
            .O(N__43485),
            .I(N__43482));
    LocalMux I__9089 (
            .O(N__43482),
            .I(N__43479));
    Span4Mux_s2_v I__9088 (
            .O(N__43479),
            .I(N__43475));
    InMux I__9087 (
            .O(N__43478),
            .I(N__43472));
    Sp12to4 I__9086 (
            .O(N__43475),
            .I(N__43467));
    LocalMux I__9085 (
            .O(N__43472),
            .I(N__43467));
    Span12Mux_s11_h I__9084 (
            .O(N__43467),
            .I(N__43464));
    Odrv12 I__9083 (
            .O(N__43464),
            .I(duty_4));
    InMux I__9082 (
            .O(N__43461),
            .I(n12462));
    InMux I__9081 (
            .O(N__43458),
            .I(N__43455));
    LocalMux I__9080 (
            .O(N__43455),
            .I(N__43452));
    Odrv12 I__9079 (
            .O(N__43452),
            .I(n20_adj_557));
    InMux I__9078 (
            .O(N__43449),
            .I(N__43443));
    InMux I__9077 (
            .O(N__43448),
            .I(N__43443));
    LocalMux I__9076 (
            .O(N__43443),
            .I(N__43440));
    Span4Mux_v I__9075 (
            .O(N__43440),
            .I(N__43437));
    Odrv4 I__9074 (
            .O(N__43437),
            .I(duty_5));
    InMux I__9073 (
            .O(N__43434),
            .I(n12463));
    InMux I__9072 (
            .O(N__43431),
            .I(N__43428));
    LocalMux I__9071 (
            .O(N__43428),
            .I(n19_adj_558));
    CascadeMux I__9070 (
            .O(N__43425),
            .I(N__43422));
    InMux I__9069 (
            .O(N__43422),
            .I(N__43416));
    InMux I__9068 (
            .O(N__43421),
            .I(N__43416));
    LocalMux I__9067 (
            .O(N__43416),
            .I(N__43413));
    Span4Mux_v I__9066 (
            .O(N__43413),
            .I(N__43410));
    Odrv4 I__9065 (
            .O(N__43410),
            .I(duty_6));
    InMux I__9064 (
            .O(N__43407),
            .I(n12464));
    CascadeMux I__9063 (
            .O(N__43404),
            .I(N__43401));
    InMux I__9062 (
            .O(N__43401),
            .I(N__43398));
    LocalMux I__9061 (
            .O(N__43398),
            .I(N__43395));
    Odrv12 I__9060 (
            .O(N__43395),
            .I(n18_adj_559));
    InMux I__9059 (
            .O(N__43392),
            .I(N__43388));
    InMux I__9058 (
            .O(N__43391),
            .I(N__43385));
    LocalMux I__9057 (
            .O(N__43388),
            .I(N__43382));
    LocalMux I__9056 (
            .O(N__43385),
            .I(N__43377));
    Span4Mux_h I__9055 (
            .O(N__43382),
            .I(N__43377));
    Odrv4 I__9054 (
            .O(N__43377),
            .I(duty_7));
    InMux I__9053 (
            .O(N__43374),
            .I(n12465));
    InMux I__9052 (
            .O(N__43371),
            .I(N__43368));
    LocalMux I__9051 (
            .O(N__43368),
            .I(N__43365));
    Odrv12 I__9050 (
            .O(N__43365),
            .I(n17_adj_560));
    InMux I__9049 (
            .O(N__43362),
            .I(bfn_12_27_0_));
    InMux I__9048 (
            .O(N__43359),
            .I(N__43356));
    LocalMux I__9047 (
            .O(N__43356),
            .I(n16_adj_563));
    InMux I__9046 (
            .O(N__43353),
            .I(N__43349));
    InMux I__9045 (
            .O(N__43352),
            .I(N__43346));
    LocalMux I__9044 (
            .O(N__43349),
            .I(N__43341));
    LocalMux I__9043 (
            .O(N__43346),
            .I(N__43341));
    Span4Mux_v I__9042 (
            .O(N__43341),
            .I(N__43338));
    Odrv4 I__9041 (
            .O(N__43338),
            .I(duty_9));
    InMux I__9040 (
            .O(N__43335),
            .I(n12467));
    InMux I__9039 (
            .O(N__43332),
            .I(N__43329));
    LocalMux I__9038 (
            .O(N__43329),
            .I(n15_adj_568));
    InMux I__9037 (
            .O(N__43326),
            .I(N__43320));
    InMux I__9036 (
            .O(N__43325),
            .I(N__43320));
    LocalMux I__9035 (
            .O(N__43320),
            .I(N__43317));
    Span4Mux_h I__9034 (
            .O(N__43317),
            .I(N__43314));
    Odrv4 I__9033 (
            .O(N__43314),
            .I(duty_10));
    InMux I__9032 (
            .O(N__43311),
            .I(n12468));
    CascadeMux I__9031 (
            .O(N__43308),
            .I(N__43305));
    InMux I__9030 (
            .O(N__43305),
            .I(N__43302));
    LocalMux I__9029 (
            .O(N__43302),
            .I(n404));
    InMux I__9028 (
            .O(N__43299),
            .I(N__43296));
    LocalMux I__9027 (
            .O(N__43296),
            .I(n2539));
    InMux I__9026 (
            .O(N__43293),
            .I(n12484));
    CascadeMux I__9025 (
            .O(N__43290),
            .I(N__43287));
    InMux I__9024 (
            .O(N__43287),
            .I(N__43284));
    LocalMux I__9023 (
            .O(N__43284),
            .I(N__43281));
    Odrv4 I__9022 (
            .O(N__43281),
            .I(n403));
    InMux I__9021 (
            .O(N__43278),
            .I(N__43275));
    LocalMux I__9020 (
            .O(N__43275),
            .I(n2538));
    InMux I__9019 (
            .O(N__43272),
            .I(n12485));
    CascadeMux I__9018 (
            .O(N__43269),
            .I(N__43266));
    InMux I__9017 (
            .O(N__43266),
            .I(N__43263));
    LocalMux I__9016 (
            .O(N__43263),
            .I(N__43260));
    Odrv12 I__9015 (
            .O(N__43260),
            .I(n402));
    InMux I__9014 (
            .O(N__43257),
            .I(n12486));
    InMux I__9013 (
            .O(N__43254),
            .I(N__43251));
    LocalMux I__9012 (
            .O(N__43251),
            .I(n2537));
    InMux I__9011 (
            .O(N__43248),
            .I(N__43245));
    LocalMux I__9010 (
            .O(N__43245),
            .I(N__43242));
    Span4Mux_h I__9009 (
            .O(N__43242),
            .I(N__43239));
    Span4Mux_h I__9008 (
            .O(N__43239),
            .I(N__43236));
    Odrv4 I__9007 (
            .O(N__43236),
            .I(encoder0_position_scaled_6));
    InMux I__9006 (
            .O(N__43233),
            .I(N__43230));
    LocalMux I__9005 (
            .O(N__43230),
            .I(N__43227));
    Span4Mux_h I__9004 (
            .O(N__43227),
            .I(N__43222));
    InMux I__9003 (
            .O(N__43226),
            .I(N__43219));
    InMux I__9002 (
            .O(N__43225),
            .I(N__43216));
    Span4Mux_v I__9001 (
            .O(N__43222),
            .I(N__43213));
    LocalMux I__9000 (
            .O(N__43219),
            .I(N__43208));
    LocalMux I__8999 (
            .O(N__43216),
            .I(N__43208));
    Span4Mux_h I__8998 (
            .O(N__43213),
            .I(N__43205));
    Span4Mux_v I__8997 (
            .O(N__43208),
            .I(N__43202));
    Odrv4 I__8996 (
            .O(N__43205),
            .I(n3109));
    Odrv4 I__8995 (
            .O(N__43202),
            .I(n3109));
    CascadeMux I__8994 (
            .O(N__43197),
            .I(N__43194));
    InMux I__8993 (
            .O(N__43194),
            .I(N__43191));
    LocalMux I__8992 (
            .O(N__43191),
            .I(N__43188));
    Span4Mux_v I__8991 (
            .O(N__43188),
            .I(N__43185));
    Span4Mux_h I__8990 (
            .O(N__43185),
            .I(N__43182));
    Odrv4 I__8989 (
            .O(N__43182),
            .I(n3176));
    InMux I__8988 (
            .O(N__43179),
            .I(N__43175));
    InMux I__8987 (
            .O(N__43178),
            .I(N__43163));
    LocalMux I__8986 (
            .O(N__43175),
            .I(N__43160));
    CascadeMux I__8985 (
            .O(N__43174),
            .I(N__43157));
    CascadeMux I__8984 (
            .O(N__43173),
            .I(N__43153));
    CascadeMux I__8983 (
            .O(N__43172),
            .I(N__43143));
    CascadeMux I__8982 (
            .O(N__43171),
            .I(N__43140));
    CascadeMux I__8981 (
            .O(N__43170),
            .I(N__43135));
    CascadeMux I__8980 (
            .O(N__43169),
            .I(N__43130));
    CascadeMux I__8979 (
            .O(N__43168),
            .I(N__43126));
    CascadeMux I__8978 (
            .O(N__43167),
            .I(N__43121));
    CascadeMux I__8977 (
            .O(N__43166),
            .I(N__43118));
    LocalMux I__8976 (
            .O(N__43163),
            .I(N__43114));
    Span4Mux_h I__8975 (
            .O(N__43160),
            .I(N__43111));
    InMux I__8974 (
            .O(N__43157),
            .I(N__43106));
    InMux I__8973 (
            .O(N__43156),
            .I(N__43106));
    InMux I__8972 (
            .O(N__43153),
            .I(N__43097));
    InMux I__8971 (
            .O(N__43152),
            .I(N__43097));
    InMux I__8970 (
            .O(N__43151),
            .I(N__43097));
    InMux I__8969 (
            .O(N__43150),
            .I(N__43097));
    CascadeMux I__8968 (
            .O(N__43149),
            .I(N__43094));
    CascadeMux I__8967 (
            .O(N__43148),
            .I(N__43090));
    CascadeMux I__8966 (
            .O(N__43147),
            .I(N__43087));
    InMux I__8965 (
            .O(N__43146),
            .I(N__43082));
    InMux I__8964 (
            .O(N__43143),
            .I(N__43073));
    InMux I__8963 (
            .O(N__43140),
            .I(N__43073));
    InMux I__8962 (
            .O(N__43139),
            .I(N__43073));
    InMux I__8961 (
            .O(N__43138),
            .I(N__43073));
    InMux I__8960 (
            .O(N__43135),
            .I(N__43066));
    InMux I__8959 (
            .O(N__43134),
            .I(N__43066));
    InMux I__8958 (
            .O(N__43133),
            .I(N__43066));
    InMux I__8957 (
            .O(N__43130),
            .I(N__43057));
    InMux I__8956 (
            .O(N__43129),
            .I(N__43057));
    InMux I__8955 (
            .O(N__43126),
            .I(N__43057));
    InMux I__8954 (
            .O(N__43125),
            .I(N__43057));
    InMux I__8953 (
            .O(N__43124),
            .I(N__43048));
    InMux I__8952 (
            .O(N__43121),
            .I(N__43048));
    InMux I__8951 (
            .O(N__43118),
            .I(N__43048));
    InMux I__8950 (
            .O(N__43117),
            .I(N__43048));
    Span4Mux_v I__8949 (
            .O(N__43114),
            .I(N__43039));
    Span4Mux_h I__8948 (
            .O(N__43111),
            .I(N__43039));
    LocalMux I__8947 (
            .O(N__43106),
            .I(N__43039));
    LocalMux I__8946 (
            .O(N__43097),
            .I(N__43039));
    InMux I__8945 (
            .O(N__43094),
            .I(N__43026));
    InMux I__8944 (
            .O(N__43093),
            .I(N__43026));
    InMux I__8943 (
            .O(N__43090),
            .I(N__43026));
    InMux I__8942 (
            .O(N__43087),
            .I(N__43026));
    InMux I__8941 (
            .O(N__43086),
            .I(N__43026));
    InMux I__8940 (
            .O(N__43085),
            .I(N__43026));
    LocalMux I__8939 (
            .O(N__43082),
            .I(n3138));
    LocalMux I__8938 (
            .O(N__43073),
            .I(n3138));
    LocalMux I__8937 (
            .O(N__43066),
            .I(n3138));
    LocalMux I__8936 (
            .O(N__43057),
            .I(n3138));
    LocalMux I__8935 (
            .O(N__43048),
            .I(n3138));
    Odrv4 I__8934 (
            .O(N__43039),
            .I(n3138));
    LocalMux I__8933 (
            .O(N__43026),
            .I(n3138));
    InMux I__8932 (
            .O(N__43011),
            .I(N__43007));
    CascadeMux I__8931 (
            .O(N__43010),
            .I(N__43003));
    LocalMux I__8930 (
            .O(N__43007),
            .I(N__43000));
    InMux I__8929 (
            .O(N__43006),
            .I(N__42995));
    InMux I__8928 (
            .O(N__43003),
            .I(N__42995));
    Span4Mux_v I__8927 (
            .O(N__43000),
            .I(N__42992));
    LocalMux I__8926 (
            .O(N__42995),
            .I(N__42989));
    Span4Mux_h I__8925 (
            .O(N__42992),
            .I(N__42986));
    Span4Mux_h I__8924 (
            .O(N__42989),
            .I(N__42983));
    Odrv4 I__8923 (
            .O(N__42986),
            .I(n3208));
    Odrv4 I__8922 (
            .O(N__42983),
            .I(n3208));
    InMux I__8921 (
            .O(N__42978),
            .I(N__42975));
    LocalMux I__8920 (
            .O(N__42975),
            .I(N__42972));
    Odrv4 I__8919 (
            .O(N__42972),
            .I(n25_adj_552));
    InMux I__8918 (
            .O(N__42969),
            .I(N__42965));
    InMux I__8917 (
            .O(N__42968),
            .I(N__42962));
    LocalMux I__8916 (
            .O(N__42965),
            .I(N__42959));
    LocalMux I__8915 (
            .O(N__42962),
            .I(N__42956));
    Span4Mux_h I__8914 (
            .O(N__42959),
            .I(N__42953));
    Odrv12 I__8913 (
            .O(N__42956),
            .I(duty_0));
    Odrv4 I__8912 (
            .O(N__42953),
            .I(duty_0));
    InMux I__8911 (
            .O(N__42948),
            .I(bfn_12_26_0_));
    InMux I__8910 (
            .O(N__42945),
            .I(N__42942));
    LocalMux I__8909 (
            .O(N__42942),
            .I(N__42939));
    Span4Mux_v I__8908 (
            .O(N__42939),
            .I(N__42936));
    Odrv4 I__8907 (
            .O(N__42936),
            .I(n24_adj_553));
    InMux I__8906 (
            .O(N__42933),
            .I(N__42929));
    InMux I__8905 (
            .O(N__42932),
            .I(N__42926));
    LocalMux I__8904 (
            .O(N__42929),
            .I(N__42923));
    LocalMux I__8903 (
            .O(N__42926),
            .I(N__42920));
    Span4Mux_h I__8902 (
            .O(N__42923),
            .I(N__42917));
    Odrv12 I__8901 (
            .O(N__42920),
            .I(duty_1));
    Odrv4 I__8900 (
            .O(N__42917),
            .I(duty_1));
    InMux I__8899 (
            .O(N__42912),
            .I(n12459));
    CascadeMux I__8898 (
            .O(N__42909),
            .I(N__42906));
    InMux I__8897 (
            .O(N__42906),
            .I(N__42903));
    LocalMux I__8896 (
            .O(N__42903),
            .I(N__42900));
    Odrv4 I__8895 (
            .O(N__42900),
            .I(n23_adj_554));
    InMux I__8894 (
            .O(N__42897),
            .I(N__42893));
    InMux I__8893 (
            .O(N__42896),
            .I(N__42890));
    LocalMux I__8892 (
            .O(N__42893),
            .I(N__42887));
    LocalMux I__8891 (
            .O(N__42890),
            .I(N__42884));
    Span4Mux_v I__8890 (
            .O(N__42887),
            .I(N__42881));
    Span4Mux_v I__8889 (
            .O(N__42884),
            .I(N__42878));
    Odrv4 I__8888 (
            .O(N__42881),
            .I(duty_2));
    Odrv4 I__8887 (
            .O(N__42878),
            .I(duty_2));
    InMux I__8886 (
            .O(N__42873),
            .I(n12460));
    InMux I__8885 (
            .O(N__42870),
            .I(N__42867));
    LocalMux I__8884 (
            .O(N__42867),
            .I(N__42862));
    InMux I__8883 (
            .O(N__42866),
            .I(N__42859));
    InMux I__8882 (
            .O(N__42865),
            .I(N__42856));
    Odrv4 I__8881 (
            .O(N__42862),
            .I(n6));
    LocalMux I__8880 (
            .O(N__42859),
            .I(n6));
    LocalMux I__8879 (
            .O(N__42856),
            .I(n6));
    CascadeMux I__8878 (
            .O(N__42849),
            .I(N__42843));
    CascadeMux I__8877 (
            .O(N__42848),
            .I(N__42840));
    InMux I__8876 (
            .O(N__42847),
            .I(N__42837));
    InMux I__8875 (
            .O(N__42846),
            .I(N__42834));
    InMux I__8874 (
            .O(N__42843),
            .I(N__42829));
    InMux I__8873 (
            .O(N__42840),
            .I(N__42829));
    LocalMux I__8872 (
            .O(N__42837),
            .I(n13641));
    LocalMux I__8871 (
            .O(N__42834),
            .I(n13641));
    LocalMux I__8870 (
            .O(N__42829),
            .I(n13641));
    CascadeMux I__8869 (
            .O(N__42822),
            .I(n13648_cascade_));
    InMux I__8868 (
            .O(N__42819),
            .I(N__42816));
    LocalMux I__8867 (
            .O(N__42816),
            .I(N__42810));
    CascadeMux I__8866 (
            .O(N__42815),
            .I(N__42807));
    CascadeMux I__8865 (
            .O(N__42814),
            .I(N__42804));
    InMux I__8864 (
            .O(N__42813),
            .I(N__42801));
    Span4Mux_h I__8863 (
            .O(N__42810),
            .I(N__42798));
    InMux I__8862 (
            .O(N__42807),
            .I(N__42793));
    InMux I__8861 (
            .O(N__42804),
            .I(N__42793));
    LocalMux I__8860 (
            .O(N__42801),
            .I(encoder0_position_27));
    Odrv4 I__8859 (
            .O(N__42798),
            .I(encoder0_position_27));
    LocalMux I__8858 (
            .O(N__42793),
            .I(encoder0_position_27));
    CascadeMux I__8857 (
            .O(N__42786),
            .I(N__42783));
    InMux I__8856 (
            .O(N__42783),
            .I(N__42779));
    InMux I__8855 (
            .O(N__42782),
            .I(N__42775));
    LocalMux I__8854 (
            .O(N__42779),
            .I(N__42772));
    InMux I__8853 (
            .O(N__42778),
            .I(N__42769));
    LocalMux I__8852 (
            .O(N__42775),
            .I(n832));
    Odrv4 I__8851 (
            .O(N__42772),
            .I(n832));
    LocalMux I__8850 (
            .O(N__42769),
            .I(n832));
    InMux I__8849 (
            .O(N__42762),
            .I(N__42759));
    LocalMux I__8848 (
            .O(N__42759),
            .I(N__42756));
    Odrv4 I__8847 (
            .O(N__42756),
            .I(n999));
    CascadeMux I__8846 (
            .O(N__42753),
            .I(N__42749));
    CascadeMux I__8845 (
            .O(N__42752),
            .I(N__42746));
    InMux I__8844 (
            .O(N__42749),
            .I(N__42742));
    InMux I__8843 (
            .O(N__42746),
            .I(N__42739));
    InMux I__8842 (
            .O(N__42745),
            .I(N__42736));
    LocalMux I__8841 (
            .O(N__42742),
            .I(n932));
    LocalMux I__8840 (
            .O(N__42739),
            .I(n932));
    LocalMux I__8839 (
            .O(N__42736),
            .I(n932));
    CascadeMux I__8838 (
            .O(N__42729),
            .I(N__42725));
    InMux I__8837 (
            .O(N__42728),
            .I(N__42721));
    InMux I__8836 (
            .O(N__42725),
            .I(N__42718));
    CascadeMux I__8835 (
            .O(N__42724),
            .I(N__42715));
    LocalMux I__8834 (
            .O(N__42721),
            .I(N__42710));
    LocalMux I__8833 (
            .O(N__42718),
            .I(N__42710));
    InMux I__8832 (
            .O(N__42715),
            .I(N__42706));
    Span4Mux_h I__8831 (
            .O(N__42710),
            .I(N__42703));
    InMux I__8830 (
            .O(N__42709),
            .I(N__42700));
    LocalMux I__8829 (
            .O(N__42706),
            .I(encoder0_position_26));
    Odrv4 I__8828 (
            .O(N__42703),
            .I(encoder0_position_26));
    LocalMux I__8827 (
            .O(N__42700),
            .I(encoder0_position_26));
    InMux I__8826 (
            .O(N__42693),
            .I(N__42690));
    LocalMux I__8825 (
            .O(N__42690),
            .I(n13650));
    CascadeMux I__8824 (
            .O(N__42687),
            .I(N__42684));
    InMux I__8823 (
            .O(N__42684),
            .I(N__42679));
    CascadeMux I__8822 (
            .O(N__42683),
            .I(N__42676));
    InMux I__8821 (
            .O(N__42682),
            .I(N__42673));
    LocalMux I__8820 (
            .O(N__42679),
            .I(N__42670));
    InMux I__8819 (
            .O(N__42676),
            .I(N__42667));
    LocalMux I__8818 (
            .O(N__42673),
            .I(n833));
    Odrv4 I__8817 (
            .O(N__42670),
            .I(n833));
    LocalMux I__8816 (
            .O(N__42667),
            .I(n833));
    InMux I__8815 (
            .O(N__42660),
            .I(N__42657));
    LocalMux I__8814 (
            .O(N__42657),
            .I(N__42654));
    Span4Mux_h I__8813 (
            .O(N__42654),
            .I(N__42651));
    Span4Mux_h I__8812 (
            .O(N__42651),
            .I(N__42648));
    Odrv4 I__8811 (
            .O(N__42648),
            .I(encoder0_position_scaled_3));
    CascadeMux I__8810 (
            .O(N__42645),
            .I(N__42642));
    InMux I__8809 (
            .O(N__42642),
            .I(N__42638));
    InMux I__8808 (
            .O(N__42641),
            .I(N__42635));
    LocalMux I__8807 (
            .O(N__42638),
            .I(n293));
    LocalMux I__8806 (
            .O(N__42635),
            .I(n293));
    InMux I__8805 (
            .O(N__42630),
            .I(N__42627));
    LocalMux I__8804 (
            .O(N__42627),
            .I(n2542));
    InMux I__8803 (
            .O(N__42624),
            .I(bfn_12_25_0_));
    CascadeMux I__8802 (
            .O(N__42621),
            .I(N__42618));
    InMux I__8801 (
            .O(N__42618),
            .I(N__42615));
    LocalMux I__8800 (
            .O(N__42615),
            .I(N__42612));
    Odrv4 I__8799 (
            .O(N__42612),
            .I(n292));
    CascadeMux I__8798 (
            .O(N__42609),
            .I(N__42606));
    InMux I__8797 (
            .O(N__42606),
            .I(N__42603));
    LocalMux I__8796 (
            .O(N__42603),
            .I(n2541));
    InMux I__8795 (
            .O(N__42600),
            .I(n12482));
    CascadeMux I__8794 (
            .O(N__42597),
            .I(N__42594));
    InMux I__8793 (
            .O(N__42594),
            .I(N__42591));
    LocalMux I__8792 (
            .O(N__42591),
            .I(n174));
    InMux I__8791 (
            .O(N__42588),
            .I(N__42585));
    LocalMux I__8790 (
            .O(N__42585),
            .I(n2540));
    InMux I__8789 (
            .O(N__42582),
            .I(n12483));
    InMux I__8788 (
            .O(N__42579),
            .I(n12499));
    CascadeMux I__8787 (
            .O(N__42576),
            .I(N__42573));
    InMux I__8786 (
            .O(N__42573),
            .I(N__42570));
    LocalMux I__8785 (
            .O(N__42570),
            .I(n1001));
    InMux I__8784 (
            .O(N__42567),
            .I(N__42563));
    InMux I__8783 (
            .O(N__42566),
            .I(N__42560));
    LocalMux I__8782 (
            .O(N__42563),
            .I(n927));
    LocalMux I__8781 (
            .O(N__42560),
            .I(n927));
    CascadeMux I__8780 (
            .O(N__42555),
            .I(n14466_cascade_));
    InMux I__8779 (
            .O(N__42552),
            .I(N__42549));
    LocalMux I__8778 (
            .O(N__42549),
            .I(n11940));
    CascadeMux I__8777 (
            .O(N__42546),
            .I(N__42543));
    InMux I__8776 (
            .O(N__42543),
            .I(N__42540));
    LocalMux I__8775 (
            .O(N__42540),
            .I(N__42535));
    InMux I__8774 (
            .O(N__42539),
            .I(N__42530));
    InMux I__8773 (
            .O(N__42538),
            .I(N__42530));
    Odrv4 I__8772 (
            .O(N__42535),
            .I(n930));
    LocalMux I__8771 (
            .O(N__42530),
            .I(n930));
    CascadeMux I__8770 (
            .O(N__42525),
            .I(n960_cascade_));
    InMux I__8769 (
            .O(N__42522),
            .I(N__42519));
    LocalMux I__8768 (
            .O(N__42519),
            .I(n997));
    CascadeMux I__8767 (
            .O(N__42516),
            .I(N__42512));
    CascadeMux I__8766 (
            .O(N__42515),
            .I(N__42508));
    InMux I__8765 (
            .O(N__42512),
            .I(N__42505));
    InMux I__8764 (
            .O(N__42511),
            .I(N__42500));
    InMux I__8763 (
            .O(N__42508),
            .I(N__42500));
    LocalMux I__8762 (
            .O(N__42505),
            .I(n929));
    LocalMux I__8761 (
            .O(N__42500),
            .I(n929));
    CascadeMux I__8760 (
            .O(N__42495),
            .I(N__42492));
    InMux I__8759 (
            .O(N__42492),
            .I(N__42489));
    LocalMux I__8758 (
            .O(N__42489),
            .I(n996));
    CascadeMux I__8757 (
            .O(N__42486),
            .I(n1028_cascade_));
    InMux I__8756 (
            .O(N__42483),
            .I(N__42480));
    LocalMux I__8755 (
            .O(N__42480),
            .I(n998));
    CascadeMux I__8754 (
            .O(N__42477),
            .I(N__42474));
    InMux I__8753 (
            .O(N__42474),
            .I(N__42470));
    CascadeMux I__8752 (
            .O(N__42473),
            .I(N__42467));
    LocalMux I__8751 (
            .O(N__42470),
            .I(N__42464));
    InMux I__8750 (
            .O(N__42467),
            .I(N__42461));
    Odrv4 I__8749 (
            .O(N__42464),
            .I(n931));
    LocalMux I__8748 (
            .O(N__42461),
            .I(n931));
    InMux I__8747 (
            .O(N__42456),
            .I(N__42453));
    LocalMux I__8746 (
            .O(N__42453),
            .I(N__42450));
    Span4Mux_h I__8745 (
            .O(N__42450),
            .I(N__42447));
    Odrv4 I__8744 (
            .O(N__42447),
            .I(encoder0_position_scaled_8));
    InMux I__8743 (
            .O(N__42444),
            .I(N__42438));
    InMux I__8742 (
            .O(N__42443),
            .I(N__42438));
    LocalMux I__8741 (
            .O(N__42438),
            .I(N__42434));
    InMux I__8740 (
            .O(N__42437),
            .I(N__42431));
    Span4Mux_h I__8739 (
            .O(N__42434),
            .I(N__42428));
    LocalMux I__8738 (
            .O(N__42431),
            .I(encoder0_position_15));
    Odrv4 I__8737 (
            .O(N__42428),
            .I(encoder0_position_15));
    InMux I__8736 (
            .O(N__42423),
            .I(N__42420));
    LocalMux I__8735 (
            .O(N__42420),
            .I(N__42416));
    InMux I__8734 (
            .O(N__42419),
            .I(N__42413));
    Span4Mux_h I__8733 (
            .O(N__42416),
            .I(N__42410));
    LocalMux I__8732 (
            .O(N__42413),
            .I(N__42407));
    Sp12to4 I__8731 (
            .O(N__42410),
            .I(N__42403));
    Span4Mux_v I__8730 (
            .O(N__42407),
            .I(N__42400));
    InMux I__8729 (
            .O(N__42406),
            .I(N__42397));
    Odrv12 I__8728 (
            .O(N__42403),
            .I(n304));
    Odrv4 I__8727 (
            .O(N__42400),
            .I(n304));
    LocalMux I__8726 (
            .O(N__42397),
            .I(n304));
    InMux I__8725 (
            .O(N__42390),
            .I(N__42387));
    LocalMux I__8724 (
            .O(N__42387),
            .I(N__42384));
    Span12Mux_h I__8723 (
            .O(N__42384),
            .I(N__42381));
    Odrv12 I__8722 (
            .O(N__42381),
            .I(n15));
    InMux I__8721 (
            .O(N__42378),
            .I(N__42375));
    LocalMux I__8720 (
            .O(N__42375),
            .I(N__42370));
    InMux I__8719 (
            .O(N__42374),
            .I(N__42367));
    InMux I__8718 (
            .O(N__42373),
            .I(N__42364));
    Span4Mux_h I__8717 (
            .O(N__42370),
            .I(N__42361));
    LocalMux I__8716 (
            .O(N__42367),
            .I(N__42358));
    LocalMux I__8715 (
            .O(N__42364),
            .I(encoder0_position_18));
    Odrv4 I__8714 (
            .O(N__42361),
            .I(encoder0_position_18));
    Odrv4 I__8713 (
            .O(N__42358),
            .I(encoder0_position_18));
    InMux I__8712 (
            .O(N__42351),
            .I(bfn_12_22_0_));
    InMux I__8711 (
            .O(N__42348),
            .I(n12493));
    InMux I__8710 (
            .O(N__42345),
            .I(n12494));
    InMux I__8709 (
            .O(N__42342),
            .I(n12495));
    InMux I__8708 (
            .O(N__42339),
            .I(n12496));
    InMux I__8707 (
            .O(N__42336),
            .I(n12497));
    InMux I__8706 (
            .O(N__42333),
            .I(n12498));
    InMux I__8705 (
            .O(N__42330),
            .I(N__42327));
    LocalMux I__8704 (
            .O(N__42327),
            .I(N__42323));
    InMux I__8703 (
            .O(N__42326),
            .I(N__42320));
    Span4Mux_h I__8702 (
            .O(N__42323),
            .I(N__42317));
    LocalMux I__8701 (
            .O(N__42320),
            .I(N__42311));
    Span4Mux_v I__8700 (
            .O(N__42317),
            .I(N__42311));
    InMux I__8699 (
            .O(N__42316),
            .I(N__42308));
    Odrv4 I__8698 (
            .O(N__42311),
            .I(n2));
    LocalMux I__8697 (
            .O(N__42308),
            .I(n2));
    InMux I__8696 (
            .O(N__42303),
            .I(N__42300));
    LocalMux I__8695 (
            .O(N__42300),
            .I(N__42297));
    Span4Mux_h I__8694 (
            .O(N__42297),
            .I(N__42294));
    Odrv4 I__8693 (
            .O(N__42294),
            .I(n16));
    InMux I__8692 (
            .O(N__42291),
            .I(N__42284));
    InMux I__8691 (
            .O(N__42290),
            .I(N__42284));
    CascadeMux I__8690 (
            .O(N__42289),
            .I(N__42281));
    LocalMux I__8689 (
            .O(N__42284),
            .I(N__42278));
    InMux I__8688 (
            .O(N__42281),
            .I(N__42275));
    Span4Mux_h I__8687 (
            .O(N__42278),
            .I(N__42272));
    LocalMux I__8686 (
            .O(N__42275),
            .I(encoder0_position_17));
    Odrv4 I__8685 (
            .O(N__42272),
            .I(encoder0_position_17));
    InMux I__8684 (
            .O(N__42267),
            .I(N__42264));
    LocalMux I__8683 (
            .O(N__42264),
            .I(N__42261));
    Span4Mux_h I__8682 (
            .O(N__42261),
            .I(N__42258));
    Odrv4 I__8681 (
            .O(N__42258),
            .I(n30));
    InMux I__8680 (
            .O(N__42255),
            .I(N__42252));
    LocalMux I__8679 (
            .O(N__42252),
            .I(N__42247));
    InMux I__8678 (
            .O(N__42251),
            .I(N__42244));
    CascadeMux I__8677 (
            .O(N__42250),
            .I(N__42241));
    Span4Mux_v I__8676 (
            .O(N__42247),
            .I(N__42236));
    LocalMux I__8675 (
            .O(N__42244),
            .I(N__42236));
    InMux I__8674 (
            .O(N__42241),
            .I(N__42233));
    Span4Mux_h I__8673 (
            .O(N__42236),
            .I(N__42230));
    LocalMux I__8672 (
            .O(N__42233),
            .I(encoder0_position_3));
    Odrv4 I__8671 (
            .O(N__42230),
            .I(encoder0_position_3));
    InMux I__8670 (
            .O(N__42225),
            .I(N__42221));
    InMux I__8669 (
            .O(N__42224),
            .I(N__42217));
    LocalMux I__8668 (
            .O(N__42221),
            .I(N__42214));
    InMux I__8667 (
            .O(N__42220),
            .I(N__42211));
    LocalMux I__8666 (
            .O(N__42217),
            .I(N__42204));
    Span4Mux_h I__8665 (
            .O(N__42214),
            .I(N__42204));
    LocalMux I__8664 (
            .O(N__42211),
            .I(N__42204));
    Span4Mux_h I__8663 (
            .O(N__42204),
            .I(N__42201));
    Sp12to4 I__8662 (
            .O(N__42201),
            .I(N__42198));
    Span12Mux_v I__8661 (
            .O(N__42198),
            .I(N__42195));
    Odrv12 I__8660 (
            .O(N__42195),
            .I(n316));
    CascadeMux I__8659 (
            .O(N__42192),
            .I(N__42168));
    CascadeMux I__8658 (
            .O(N__42191),
            .I(N__42165));
    CascadeMux I__8657 (
            .O(N__42190),
            .I(N__42162));
    CascadeMux I__8656 (
            .O(N__42189),
            .I(N__42159));
    CascadeMux I__8655 (
            .O(N__42188),
            .I(N__42156));
    CascadeMux I__8654 (
            .O(N__42187),
            .I(N__42153));
    CascadeMux I__8653 (
            .O(N__42186),
            .I(N__42150));
    CascadeMux I__8652 (
            .O(N__42185),
            .I(N__42147));
    CascadeMux I__8651 (
            .O(N__42184),
            .I(N__42144));
    CascadeMux I__8650 (
            .O(N__42183),
            .I(N__42141));
    CascadeMux I__8649 (
            .O(N__42182),
            .I(N__42138));
    CascadeMux I__8648 (
            .O(N__42181),
            .I(N__42135));
    CascadeMux I__8647 (
            .O(N__42180),
            .I(N__42132));
    CascadeMux I__8646 (
            .O(N__42179),
            .I(N__42129));
    CascadeMux I__8645 (
            .O(N__42178),
            .I(N__42125));
    CascadeMux I__8644 (
            .O(N__42177),
            .I(N__42122));
    CascadeMux I__8643 (
            .O(N__42176),
            .I(N__42119));
    CascadeMux I__8642 (
            .O(N__42175),
            .I(N__42116));
    CascadeMux I__8641 (
            .O(N__42174),
            .I(N__42112));
    CascadeMux I__8640 (
            .O(N__42173),
            .I(N__42109));
    CascadeMux I__8639 (
            .O(N__42172),
            .I(N__42106));
    CascadeMux I__8638 (
            .O(N__42171),
            .I(N__42103));
    InMux I__8637 (
            .O(N__42168),
            .I(N__42093));
    InMux I__8636 (
            .O(N__42165),
            .I(N__42093));
    InMux I__8635 (
            .O(N__42162),
            .I(N__42093));
    InMux I__8634 (
            .O(N__42159),
            .I(N__42093));
    InMux I__8633 (
            .O(N__42156),
            .I(N__42084));
    InMux I__8632 (
            .O(N__42153),
            .I(N__42084));
    InMux I__8631 (
            .O(N__42150),
            .I(N__42084));
    InMux I__8630 (
            .O(N__42147),
            .I(N__42084));
    InMux I__8629 (
            .O(N__42144),
            .I(N__42075));
    InMux I__8628 (
            .O(N__42141),
            .I(N__42075));
    InMux I__8627 (
            .O(N__42138),
            .I(N__42075));
    InMux I__8626 (
            .O(N__42135),
            .I(N__42075));
    InMux I__8625 (
            .O(N__42132),
            .I(N__42066));
    InMux I__8624 (
            .O(N__42129),
            .I(N__42066));
    InMux I__8623 (
            .O(N__42128),
            .I(N__42066));
    InMux I__8622 (
            .O(N__42125),
            .I(N__42066));
    InMux I__8621 (
            .O(N__42122),
            .I(N__42057));
    InMux I__8620 (
            .O(N__42119),
            .I(N__42057));
    InMux I__8619 (
            .O(N__42116),
            .I(N__42057));
    InMux I__8618 (
            .O(N__42115),
            .I(N__42057));
    InMux I__8617 (
            .O(N__42112),
            .I(N__42048));
    InMux I__8616 (
            .O(N__42109),
            .I(N__42048));
    InMux I__8615 (
            .O(N__42106),
            .I(N__42048));
    InMux I__8614 (
            .O(N__42103),
            .I(N__42048));
    CascadeMux I__8613 (
            .O(N__42102),
            .I(N__42045));
    LocalMux I__8612 (
            .O(N__42093),
            .I(N__42040));
    LocalMux I__8611 (
            .O(N__42084),
            .I(N__42040));
    LocalMux I__8610 (
            .O(N__42075),
            .I(N__42033));
    LocalMux I__8609 (
            .O(N__42066),
            .I(N__42033));
    LocalMux I__8608 (
            .O(N__42057),
            .I(N__42033));
    LocalMux I__8607 (
            .O(N__42048),
            .I(N__42030));
    InMux I__8606 (
            .O(N__42045),
            .I(N__42027));
    Span4Mux_v I__8605 (
            .O(N__42040),
            .I(N__42022));
    Span4Mux_v I__8604 (
            .O(N__42033),
            .I(N__42022));
    Span4Mux_h I__8603 (
            .O(N__42030),
            .I(N__42017));
    LocalMux I__8602 (
            .O(N__42027),
            .I(N__42017));
    Span4Mux_h I__8601 (
            .O(N__42022),
            .I(N__42012));
    Span4Mux_v I__8600 (
            .O(N__42017),
            .I(N__42012));
    Odrv4 I__8599 (
            .O(N__42012),
            .I(n2_adj_623));
    InMux I__8598 (
            .O(N__42009),
            .I(N__42006));
    LocalMux I__8597 (
            .O(N__42006),
            .I(N__42003));
    Span4Mux_v I__8596 (
            .O(N__42003),
            .I(N__42000));
    Span4Mux_h I__8595 (
            .O(N__42000),
            .I(N__41997));
    Odrv4 I__8594 (
            .O(N__41997),
            .I(encoder0_position_scaled_7));
    InMux I__8593 (
            .O(N__41994),
            .I(N__41989));
    InMux I__8592 (
            .O(N__41993),
            .I(N__41986));
    CascadeMux I__8591 (
            .O(N__41992),
            .I(N__41983));
    LocalMux I__8590 (
            .O(N__41989),
            .I(N__41980));
    LocalMux I__8589 (
            .O(N__41986),
            .I(N__41977));
    InMux I__8588 (
            .O(N__41983),
            .I(N__41974));
    Span4Mux_h I__8587 (
            .O(N__41980),
            .I(N__41971));
    Span4Mux_h I__8586 (
            .O(N__41977),
            .I(N__41968));
    LocalMux I__8585 (
            .O(N__41974),
            .I(encoder0_position_23));
    Odrv4 I__8584 (
            .O(N__41971),
            .I(encoder0_position_23));
    Odrv4 I__8583 (
            .O(N__41968),
            .I(encoder0_position_23));
    CascadeMux I__8582 (
            .O(N__41961),
            .I(N__41958));
    InMux I__8581 (
            .O(N__41958),
            .I(N__41955));
    LocalMux I__8580 (
            .O(N__41955),
            .I(N__41952));
    Span4Mux_v I__8579 (
            .O(N__41952),
            .I(N__41949));
    Odrv4 I__8578 (
            .O(N__41949),
            .I(n10_adj_631));
    CascadeMux I__8577 (
            .O(N__41946),
            .I(N__41943));
    InMux I__8576 (
            .O(N__41943),
            .I(N__41940));
    LocalMux I__8575 (
            .O(N__41940),
            .I(N__41937));
    Span4Mux_v I__8574 (
            .O(N__41937),
            .I(N__41934));
    Odrv4 I__8573 (
            .O(N__41934),
            .I(n18_adj_639));
    InMux I__8572 (
            .O(N__41931),
            .I(N__41928));
    LocalMux I__8571 (
            .O(N__41928),
            .I(N__41925));
    Span4Mux_v I__8570 (
            .O(N__41925),
            .I(N__41922));
    Odrv4 I__8569 (
            .O(N__41922),
            .I(n17));
    CascadeMux I__8568 (
            .O(N__41919),
            .I(N__41915));
    InMux I__8567 (
            .O(N__41918),
            .I(N__41912));
    InMux I__8566 (
            .O(N__41915),
            .I(N__41909));
    LocalMux I__8565 (
            .O(N__41912),
            .I(N__41905));
    LocalMux I__8564 (
            .O(N__41909),
            .I(N__41902));
    InMux I__8563 (
            .O(N__41908),
            .I(N__41899));
    Span4Mux_h I__8562 (
            .O(N__41905),
            .I(N__41896));
    Span4Mux_v I__8561 (
            .O(N__41902),
            .I(N__41893));
    LocalMux I__8560 (
            .O(N__41899),
            .I(encoder0_position_16));
    Odrv4 I__8559 (
            .O(N__41896),
            .I(encoder0_position_16));
    Odrv4 I__8558 (
            .O(N__41893),
            .I(encoder0_position_16));
    InMux I__8557 (
            .O(N__41886),
            .I(N__41883));
    LocalMux I__8556 (
            .O(N__41883),
            .I(N__41880));
    Span4Mux_h I__8555 (
            .O(N__41880),
            .I(N__41877));
    Odrv4 I__8554 (
            .O(N__41877),
            .I(n18));
    InMux I__8553 (
            .O(N__41874),
            .I(bfn_12_19_0_));
    CascadeMux I__8552 (
            .O(N__41871),
            .I(N__41868));
    InMux I__8551 (
            .O(N__41868),
            .I(N__41865));
    LocalMux I__8550 (
            .O(N__41865),
            .I(N__41862));
    Odrv4 I__8549 (
            .O(N__41862),
            .I(n1885));
    CascadeMux I__8548 (
            .O(N__41859),
            .I(n1722_cascade_));
    InMux I__8547 (
            .O(N__41856),
            .I(N__41851));
    InMux I__8546 (
            .O(N__41855),
            .I(N__41848));
    InMux I__8545 (
            .O(N__41854),
            .I(N__41845));
    LocalMux I__8544 (
            .O(N__41851),
            .I(n1821));
    LocalMux I__8543 (
            .O(N__41848),
            .I(n1821));
    LocalMux I__8542 (
            .O(N__41845),
            .I(n1821));
    CascadeMux I__8541 (
            .O(N__41838),
            .I(N__41835));
    InMux I__8540 (
            .O(N__41835),
            .I(N__41831));
    CascadeMux I__8539 (
            .O(N__41834),
            .I(N__41828));
    LocalMux I__8538 (
            .O(N__41831),
            .I(N__41824));
    InMux I__8537 (
            .O(N__41828),
            .I(N__41821));
    InMux I__8536 (
            .O(N__41827),
            .I(N__41818));
    Span4Mux_h I__8535 (
            .O(N__41824),
            .I(N__41815));
    LocalMux I__8534 (
            .O(N__41821),
            .I(N__41810));
    LocalMux I__8533 (
            .O(N__41818),
            .I(N__41810));
    Odrv4 I__8532 (
            .O(N__41815),
            .I(n1827));
    Odrv4 I__8531 (
            .O(N__41810),
            .I(n1827));
    InMux I__8530 (
            .O(N__41805),
            .I(N__41800));
    CascadeMux I__8529 (
            .O(N__41804),
            .I(N__41797));
    CascadeMux I__8528 (
            .O(N__41803),
            .I(N__41793));
    LocalMux I__8527 (
            .O(N__41800),
            .I(N__41786));
    InMux I__8526 (
            .O(N__41797),
            .I(N__41780));
    InMux I__8525 (
            .O(N__41796),
            .I(N__41780));
    InMux I__8524 (
            .O(N__41793),
            .I(N__41777));
    CascadeMux I__8523 (
            .O(N__41792),
            .I(N__41774));
    CascadeMux I__8522 (
            .O(N__41791),
            .I(N__41771));
    CascadeMux I__8521 (
            .O(N__41790),
            .I(N__41764));
    CascadeMux I__8520 (
            .O(N__41789),
            .I(N__41761));
    Span12Mux_s10_h I__8519 (
            .O(N__41786),
            .I(N__41755));
    InMux I__8518 (
            .O(N__41785),
            .I(N__41752));
    LocalMux I__8517 (
            .O(N__41780),
            .I(N__41747));
    LocalMux I__8516 (
            .O(N__41777),
            .I(N__41747));
    InMux I__8515 (
            .O(N__41774),
            .I(N__41738));
    InMux I__8514 (
            .O(N__41771),
            .I(N__41738));
    InMux I__8513 (
            .O(N__41770),
            .I(N__41738));
    InMux I__8512 (
            .O(N__41769),
            .I(N__41738));
    InMux I__8511 (
            .O(N__41768),
            .I(N__41727));
    InMux I__8510 (
            .O(N__41767),
            .I(N__41727));
    InMux I__8509 (
            .O(N__41764),
            .I(N__41727));
    InMux I__8508 (
            .O(N__41761),
            .I(N__41727));
    InMux I__8507 (
            .O(N__41760),
            .I(N__41727));
    InMux I__8506 (
            .O(N__41759),
            .I(N__41722));
    InMux I__8505 (
            .O(N__41758),
            .I(N__41722));
    Odrv12 I__8504 (
            .O(N__41755),
            .I(n1752));
    LocalMux I__8503 (
            .O(N__41752),
            .I(n1752));
    Odrv4 I__8502 (
            .O(N__41747),
            .I(n1752));
    LocalMux I__8501 (
            .O(N__41738),
            .I(n1752));
    LocalMux I__8500 (
            .O(N__41727),
            .I(n1752));
    LocalMux I__8499 (
            .O(N__41722),
            .I(n1752));
    CascadeMux I__8498 (
            .O(N__41709),
            .I(N__41706));
    InMux I__8497 (
            .O(N__41706),
            .I(N__41703));
    LocalMux I__8496 (
            .O(N__41703),
            .I(N__41700));
    Span4Mux_h I__8495 (
            .O(N__41700),
            .I(N__41697));
    Odrv4 I__8494 (
            .O(N__41697),
            .I(n16_adj_637));
    CascadeMux I__8493 (
            .O(N__41694),
            .I(N__41690));
    CascadeMux I__8492 (
            .O(N__41693),
            .I(N__41687));
    InMux I__8491 (
            .O(N__41690),
            .I(N__41684));
    InMux I__8490 (
            .O(N__41687),
            .I(N__41681));
    LocalMux I__8489 (
            .O(N__41684),
            .I(n1826));
    LocalMux I__8488 (
            .O(N__41681),
            .I(n1826));
    InMux I__8487 (
            .O(N__41676),
            .I(N__41673));
    LocalMux I__8486 (
            .O(N__41673),
            .I(N__41670));
    Span4Mux_h I__8485 (
            .O(N__41670),
            .I(N__41667));
    Odrv4 I__8484 (
            .O(N__41667),
            .I(n1893));
    InMux I__8483 (
            .O(N__41664),
            .I(bfn_12_18_0_));
    CascadeMux I__8482 (
            .O(N__41661),
            .I(N__41657));
    InMux I__8481 (
            .O(N__41660),
            .I(N__41653));
    InMux I__8480 (
            .O(N__41657),
            .I(N__41650));
    InMux I__8479 (
            .O(N__41656),
            .I(N__41647));
    LocalMux I__8478 (
            .O(N__41653),
            .I(n1825));
    LocalMux I__8477 (
            .O(N__41650),
            .I(n1825));
    LocalMux I__8476 (
            .O(N__41647),
            .I(n1825));
    InMux I__8475 (
            .O(N__41640),
            .I(N__41637));
    LocalMux I__8474 (
            .O(N__41637),
            .I(N__41634));
    Odrv4 I__8473 (
            .O(N__41634),
            .I(n1892));
    InMux I__8472 (
            .O(N__41631),
            .I(n12600));
    CascadeMux I__8471 (
            .O(N__41628),
            .I(N__41623));
    CascadeMux I__8470 (
            .O(N__41627),
            .I(N__41620));
    InMux I__8469 (
            .O(N__41626),
            .I(N__41617));
    InMux I__8468 (
            .O(N__41623),
            .I(N__41614));
    InMux I__8467 (
            .O(N__41620),
            .I(N__41611));
    LocalMux I__8466 (
            .O(N__41617),
            .I(n1824));
    LocalMux I__8465 (
            .O(N__41614),
            .I(n1824));
    LocalMux I__8464 (
            .O(N__41611),
            .I(n1824));
    InMux I__8463 (
            .O(N__41604),
            .I(N__41601));
    LocalMux I__8462 (
            .O(N__41601),
            .I(N__41598));
    Odrv4 I__8461 (
            .O(N__41598),
            .I(n1891));
    InMux I__8460 (
            .O(N__41595),
            .I(n12601));
    CascadeMux I__8459 (
            .O(N__41592),
            .I(N__41588));
    InMux I__8458 (
            .O(N__41591),
            .I(N__41584));
    InMux I__8457 (
            .O(N__41588),
            .I(N__41581));
    InMux I__8456 (
            .O(N__41587),
            .I(N__41578));
    LocalMux I__8455 (
            .O(N__41584),
            .I(n1823));
    LocalMux I__8454 (
            .O(N__41581),
            .I(n1823));
    LocalMux I__8453 (
            .O(N__41578),
            .I(n1823));
    CascadeMux I__8452 (
            .O(N__41571),
            .I(N__41568));
    InMux I__8451 (
            .O(N__41568),
            .I(N__41565));
    LocalMux I__8450 (
            .O(N__41565),
            .I(N__41562));
    Span4Mux_h I__8449 (
            .O(N__41562),
            .I(N__41559));
    Odrv4 I__8448 (
            .O(N__41559),
            .I(n1890));
    InMux I__8447 (
            .O(N__41556),
            .I(n12602));
    InMux I__8446 (
            .O(N__41553),
            .I(N__41549));
    CascadeMux I__8445 (
            .O(N__41552),
            .I(N__41546));
    LocalMux I__8444 (
            .O(N__41549),
            .I(N__41543));
    InMux I__8443 (
            .O(N__41546),
            .I(N__41540));
    Span4Mux_h I__8442 (
            .O(N__41543),
            .I(N__41536));
    LocalMux I__8441 (
            .O(N__41540),
            .I(N__41533));
    InMux I__8440 (
            .O(N__41539),
            .I(N__41530));
    Odrv4 I__8439 (
            .O(N__41536),
            .I(n1822));
    Odrv4 I__8438 (
            .O(N__41533),
            .I(n1822));
    LocalMux I__8437 (
            .O(N__41530),
            .I(n1822));
    CascadeMux I__8436 (
            .O(N__41523),
            .I(N__41520));
    InMux I__8435 (
            .O(N__41520),
            .I(N__41517));
    LocalMux I__8434 (
            .O(N__41517),
            .I(N__41514));
    Odrv12 I__8433 (
            .O(N__41514),
            .I(n1889));
    InMux I__8432 (
            .O(N__41511),
            .I(n12603));
    InMux I__8431 (
            .O(N__41508),
            .I(N__41505));
    LocalMux I__8430 (
            .O(N__41505),
            .I(n1888));
    InMux I__8429 (
            .O(N__41502),
            .I(n12604));
    CascadeMux I__8428 (
            .O(N__41499),
            .I(N__41496));
    InMux I__8427 (
            .O(N__41496),
            .I(N__41492));
    InMux I__8426 (
            .O(N__41495),
            .I(N__41489));
    LocalMux I__8425 (
            .O(N__41492),
            .I(N__41486));
    LocalMux I__8424 (
            .O(N__41489),
            .I(n1820));
    Odrv4 I__8423 (
            .O(N__41486),
            .I(n1820));
    InMux I__8422 (
            .O(N__41481),
            .I(N__41478));
    LocalMux I__8421 (
            .O(N__41478),
            .I(n1887));
    InMux I__8420 (
            .O(N__41475),
            .I(n12605));
    CascadeMux I__8419 (
            .O(N__41472),
            .I(N__41468));
    InMux I__8418 (
            .O(N__41471),
            .I(N__41465));
    InMux I__8417 (
            .O(N__41468),
            .I(N__41462));
    LocalMux I__8416 (
            .O(N__41465),
            .I(n1819));
    LocalMux I__8415 (
            .O(N__41462),
            .I(n1819));
    InMux I__8414 (
            .O(N__41457),
            .I(N__41454));
    LocalMux I__8413 (
            .O(N__41454),
            .I(n1886));
    InMux I__8412 (
            .O(N__41451),
            .I(n12606));
    InMux I__8411 (
            .O(N__41448),
            .I(N__41445));
    LocalMux I__8410 (
            .O(N__41445),
            .I(N__41442));
    Odrv4 I__8409 (
            .O(N__41442),
            .I(n1901));
    InMux I__8408 (
            .O(N__41439),
            .I(bfn_12_17_0_));
    CascadeMux I__8407 (
            .O(N__41436),
            .I(N__41433));
    InMux I__8406 (
            .O(N__41433),
            .I(N__41428));
    InMux I__8405 (
            .O(N__41432),
            .I(N__41425));
    InMux I__8404 (
            .O(N__41431),
            .I(N__41422));
    LocalMux I__8403 (
            .O(N__41428),
            .I(N__41419));
    LocalMux I__8402 (
            .O(N__41425),
            .I(n1833));
    LocalMux I__8401 (
            .O(N__41422),
            .I(n1833));
    Odrv4 I__8400 (
            .O(N__41419),
            .I(n1833));
    InMux I__8399 (
            .O(N__41412),
            .I(N__41409));
    LocalMux I__8398 (
            .O(N__41409),
            .I(N__41406));
    Span4Mux_v I__8397 (
            .O(N__41406),
            .I(N__41403));
    Odrv4 I__8396 (
            .O(N__41403),
            .I(n1900));
    InMux I__8395 (
            .O(N__41400),
            .I(n12592));
    CascadeMux I__8394 (
            .O(N__41397),
            .I(N__41393));
    CascadeMux I__8393 (
            .O(N__41396),
            .I(N__41390));
    InMux I__8392 (
            .O(N__41393),
            .I(N__41387));
    InMux I__8391 (
            .O(N__41390),
            .I(N__41384));
    LocalMux I__8390 (
            .O(N__41387),
            .I(N__41381));
    LocalMux I__8389 (
            .O(N__41384),
            .I(n1832));
    Odrv4 I__8388 (
            .O(N__41381),
            .I(n1832));
    InMux I__8387 (
            .O(N__41376),
            .I(N__41373));
    LocalMux I__8386 (
            .O(N__41373),
            .I(N__41370));
    Odrv4 I__8385 (
            .O(N__41370),
            .I(n1899));
    InMux I__8384 (
            .O(N__41367),
            .I(n12593));
    CascadeMux I__8383 (
            .O(N__41364),
            .I(N__41360));
    CascadeMux I__8382 (
            .O(N__41363),
            .I(N__41357));
    InMux I__8381 (
            .O(N__41360),
            .I(N__41354));
    InMux I__8380 (
            .O(N__41357),
            .I(N__41350));
    LocalMux I__8379 (
            .O(N__41354),
            .I(N__41347));
    InMux I__8378 (
            .O(N__41353),
            .I(N__41344));
    LocalMux I__8377 (
            .O(N__41350),
            .I(n1831));
    Odrv4 I__8376 (
            .O(N__41347),
            .I(n1831));
    LocalMux I__8375 (
            .O(N__41344),
            .I(n1831));
    InMux I__8374 (
            .O(N__41337),
            .I(N__41334));
    LocalMux I__8373 (
            .O(N__41334),
            .I(N__41331));
    Span4Mux_v I__8372 (
            .O(N__41331),
            .I(N__41328));
    Odrv4 I__8371 (
            .O(N__41328),
            .I(n1898));
    InMux I__8370 (
            .O(N__41325),
            .I(n12594));
    CascadeMux I__8369 (
            .O(N__41322),
            .I(N__41317));
    InMux I__8368 (
            .O(N__41321),
            .I(N__41312));
    InMux I__8367 (
            .O(N__41320),
            .I(N__41312));
    InMux I__8366 (
            .O(N__41317),
            .I(N__41309));
    LocalMux I__8365 (
            .O(N__41312),
            .I(N__41304));
    LocalMux I__8364 (
            .O(N__41309),
            .I(N__41304));
    Odrv4 I__8363 (
            .O(N__41304),
            .I(n1830));
    InMux I__8362 (
            .O(N__41301),
            .I(N__41298));
    LocalMux I__8361 (
            .O(N__41298),
            .I(n1897));
    InMux I__8360 (
            .O(N__41295),
            .I(n12595));
    CascadeMux I__8359 (
            .O(N__41292),
            .I(N__41287));
    InMux I__8358 (
            .O(N__41291),
            .I(N__41282));
    InMux I__8357 (
            .O(N__41290),
            .I(N__41282));
    InMux I__8356 (
            .O(N__41287),
            .I(N__41279));
    LocalMux I__8355 (
            .O(N__41282),
            .I(n1829));
    LocalMux I__8354 (
            .O(N__41279),
            .I(n1829));
    CascadeMux I__8353 (
            .O(N__41274),
            .I(N__41271));
    InMux I__8352 (
            .O(N__41271),
            .I(N__41268));
    LocalMux I__8351 (
            .O(N__41268),
            .I(n1896));
    InMux I__8350 (
            .O(N__41265),
            .I(n12596));
    CascadeMux I__8349 (
            .O(N__41262),
            .I(N__41258));
    InMux I__8348 (
            .O(N__41261),
            .I(N__41254));
    InMux I__8347 (
            .O(N__41258),
            .I(N__41251));
    InMux I__8346 (
            .O(N__41257),
            .I(N__41248));
    LocalMux I__8345 (
            .O(N__41254),
            .I(n1828));
    LocalMux I__8344 (
            .O(N__41251),
            .I(n1828));
    LocalMux I__8343 (
            .O(N__41248),
            .I(n1828));
    CascadeMux I__8342 (
            .O(N__41241),
            .I(N__41238));
    InMux I__8341 (
            .O(N__41238),
            .I(N__41235));
    LocalMux I__8340 (
            .O(N__41235),
            .I(N__41232));
    Odrv4 I__8339 (
            .O(N__41232),
            .I(n1895));
    InMux I__8338 (
            .O(N__41229),
            .I(n12597));
    InMux I__8337 (
            .O(N__41226),
            .I(N__41223));
    LocalMux I__8336 (
            .O(N__41223),
            .I(N__41220));
    Odrv4 I__8335 (
            .O(N__41220),
            .I(n1894));
    InMux I__8334 (
            .O(N__41217),
            .I(n12598));
    InMux I__8333 (
            .O(N__41214),
            .I(N__41211));
    LocalMux I__8332 (
            .O(N__41211),
            .I(n6_adj_677));
    InMux I__8331 (
            .O(N__41208),
            .I(n13106));
    CascadeMux I__8330 (
            .O(N__41205),
            .I(N__41201));
    CascadeMux I__8329 (
            .O(N__41204),
            .I(N__41198));
    InMux I__8328 (
            .O(N__41201),
            .I(N__41192));
    InMux I__8327 (
            .O(N__41198),
            .I(N__41192));
    InMux I__8326 (
            .O(N__41197),
            .I(N__41189));
    LocalMux I__8325 (
            .O(N__41192),
            .I(blink_counter_21));
    LocalMux I__8324 (
            .O(N__41189),
            .I(blink_counter_21));
    InMux I__8323 (
            .O(N__41184),
            .I(n13107));
    InMux I__8322 (
            .O(N__41181),
            .I(N__41174));
    InMux I__8321 (
            .O(N__41180),
            .I(N__41174));
    InMux I__8320 (
            .O(N__41179),
            .I(N__41171));
    LocalMux I__8319 (
            .O(N__41174),
            .I(blink_counter_22));
    LocalMux I__8318 (
            .O(N__41171),
            .I(blink_counter_22));
    InMux I__8317 (
            .O(N__41166),
            .I(n13108));
    InMux I__8316 (
            .O(N__41163),
            .I(N__41156));
    InMux I__8315 (
            .O(N__41162),
            .I(N__41156));
    InMux I__8314 (
            .O(N__41161),
            .I(N__41153));
    LocalMux I__8313 (
            .O(N__41156),
            .I(blink_counter_23));
    LocalMux I__8312 (
            .O(N__41153),
            .I(blink_counter_23));
    InMux I__8311 (
            .O(N__41148),
            .I(n13109));
    InMux I__8310 (
            .O(N__41145),
            .I(N__41138));
    InMux I__8309 (
            .O(N__41144),
            .I(N__41138));
    InMux I__8308 (
            .O(N__41143),
            .I(N__41135));
    LocalMux I__8307 (
            .O(N__41138),
            .I(blink_counter_24));
    LocalMux I__8306 (
            .O(N__41135),
            .I(blink_counter_24));
    InMux I__8305 (
            .O(N__41130),
            .I(bfn_11_32_0_));
    InMux I__8304 (
            .O(N__41127),
            .I(n13111));
    InMux I__8303 (
            .O(N__41124),
            .I(N__41121));
    LocalMux I__8302 (
            .O(N__41121),
            .I(N__41117));
    InMux I__8301 (
            .O(N__41120),
            .I(N__41114));
    Odrv4 I__8300 (
            .O(N__41117),
            .I(blink_counter_25));
    LocalMux I__8299 (
            .O(N__41114),
            .I(blink_counter_25));
    InMux I__8298 (
            .O(N__41109),
            .I(N__41106));
    LocalMux I__8297 (
            .O(N__41106),
            .I(N__41103));
    Odrv4 I__8296 (
            .O(N__41103),
            .I(pwm_setpoint_23_N_171_19));
    InMux I__8295 (
            .O(N__41100),
            .I(N__41097));
    LocalMux I__8294 (
            .O(N__41097),
            .I(N__41094));
    Odrv4 I__8293 (
            .O(N__41094),
            .I(n8_adj_588));
    InMux I__8292 (
            .O(N__41091),
            .I(N__41088));
    LocalMux I__8291 (
            .O(N__41088),
            .I(N__41085));
    Odrv4 I__8290 (
            .O(N__41085),
            .I(n5_adj_585));
    InMux I__8289 (
            .O(N__41082),
            .I(N__41079));
    LocalMux I__8288 (
            .O(N__41079),
            .I(n14_adj_685));
    InMux I__8287 (
            .O(N__41076),
            .I(n13098));
    InMux I__8286 (
            .O(N__41073),
            .I(N__41070));
    LocalMux I__8285 (
            .O(N__41070),
            .I(n13_adj_684));
    InMux I__8284 (
            .O(N__41067),
            .I(n13099));
    InMux I__8283 (
            .O(N__41064),
            .I(N__41061));
    LocalMux I__8282 (
            .O(N__41061),
            .I(n12_adj_683));
    InMux I__8281 (
            .O(N__41058),
            .I(n13100));
    InMux I__8280 (
            .O(N__41055),
            .I(N__41052));
    LocalMux I__8279 (
            .O(N__41052),
            .I(n11_adj_682));
    InMux I__8278 (
            .O(N__41049),
            .I(n13101));
    InMux I__8277 (
            .O(N__41046),
            .I(N__41043));
    LocalMux I__8276 (
            .O(N__41043),
            .I(n10_adj_681));
    InMux I__8275 (
            .O(N__41040),
            .I(bfn_11_31_0_));
    InMux I__8274 (
            .O(N__41037),
            .I(N__41034));
    LocalMux I__8273 (
            .O(N__41034),
            .I(n9_adj_680));
    InMux I__8272 (
            .O(N__41031),
            .I(n13103));
    InMux I__8271 (
            .O(N__41028),
            .I(N__41025));
    LocalMux I__8270 (
            .O(N__41025),
            .I(n8_adj_679));
    InMux I__8269 (
            .O(N__41022),
            .I(n13104));
    InMux I__8268 (
            .O(N__41019),
            .I(N__41016));
    LocalMux I__8267 (
            .O(N__41016),
            .I(n7_adj_678));
    InMux I__8266 (
            .O(N__41013),
            .I(n13105));
    InMux I__8265 (
            .O(N__41010),
            .I(N__41007));
    LocalMux I__8264 (
            .O(N__41007),
            .I(n23_adj_694));
    InMux I__8263 (
            .O(N__41004),
            .I(n13089));
    InMux I__8262 (
            .O(N__41001),
            .I(N__40998));
    LocalMux I__8261 (
            .O(N__40998),
            .I(n22_adj_693));
    InMux I__8260 (
            .O(N__40995),
            .I(n13090));
    InMux I__8259 (
            .O(N__40992),
            .I(N__40989));
    LocalMux I__8258 (
            .O(N__40989),
            .I(n21_adj_692));
    InMux I__8257 (
            .O(N__40986),
            .I(n13091));
    InMux I__8256 (
            .O(N__40983),
            .I(N__40980));
    LocalMux I__8255 (
            .O(N__40980),
            .I(n20_adj_691));
    InMux I__8254 (
            .O(N__40977),
            .I(n13092));
    InMux I__8253 (
            .O(N__40974),
            .I(N__40971));
    LocalMux I__8252 (
            .O(N__40971),
            .I(n19_adj_690));
    InMux I__8251 (
            .O(N__40968),
            .I(n13093));
    InMux I__8250 (
            .O(N__40965),
            .I(N__40962));
    LocalMux I__8249 (
            .O(N__40962),
            .I(n18_adj_689));
    InMux I__8248 (
            .O(N__40959),
            .I(bfn_11_30_0_));
    InMux I__8247 (
            .O(N__40956),
            .I(N__40953));
    LocalMux I__8246 (
            .O(N__40953),
            .I(n17_adj_688));
    InMux I__8245 (
            .O(N__40950),
            .I(n13095));
    InMux I__8244 (
            .O(N__40947),
            .I(N__40944));
    LocalMux I__8243 (
            .O(N__40944),
            .I(n16_adj_687));
    InMux I__8242 (
            .O(N__40941),
            .I(n13096));
    InMux I__8241 (
            .O(N__40938),
            .I(N__40935));
    LocalMux I__8240 (
            .O(N__40935),
            .I(n15_adj_686));
    InMux I__8239 (
            .O(N__40932),
            .I(n13097));
    InMux I__8238 (
            .O(N__40929),
            .I(N__40926));
    LocalMux I__8237 (
            .O(N__40926),
            .I(n12_adj_661));
    InMux I__8236 (
            .O(N__40923),
            .I(N__40920));
    LocalMux I__8235 (
            .O(N__40920),
            .I(N__40917));
    Span4Mux_h I__8234 (
            .O(N__40917),
            .I(N__40914));
    Odrv4 I__8233 (
            .O(N__40914),
            .I(pwm_setpoint_23_N_171_7));
    InMux I__8232 (
            .O(N__40911),
            .I(N__40906));
    InMux I__8231 (
            .O(N__40910),
            .I(N__40901));
    InMux I__8230 (
            .O(N__40909),
            .I(N__40901));
    LocalMux I__8229 (
            .O(N__40906),
            .I(pwm_setpoint_16));
    LocalMux I__8228 (
            .O(N__40901),
            .I(pwm_setpoint_16));
    InMux I__8227 (
            .O(N__40896),
            .I(N__40891));
    InMux I__8226 (
            .O(N__40895),
            .I(N__40886));
    InMux I__8225 (
            .O(N__40894),
            .I(N__40886));
    LocalMux I__8224 (
            .O(N__40891),
            .I(pwm_setpoint_7));
    LocalMux I__8223 (
            .O(N__40886),
            .I(pwm_setpoint_7));
    InMux I__8222 (
            .O(N__40881),
            .I(N__40878));
    LocalMux I__8221 (
            .O(N__40878),
            .I(n15119));
    InMux I__8220 (
            .O(N__40875),
            .I(N__40872));
    LocalMux I__8219 (
            .O(N__40872),
            .I(N__40869));
    Span4Mux_h I__8218 (
            .O(N__40869),
            .I(N__40866));
    Span4Mux_v I__8217 (
            .O(N__40866),
            .I(N__40863));
    Odrv4 I__8216 (
            .O(N__40863),
            .I(encoder0_position_scaled_9));
    InMux I__8215 (
            .O(N__40860),
            .I(N__40857));
    LocalMux I__8214 (
            .O(N__40857),
            .I(n26_adj_697));
    InMux I__8213 (
            .O(N__40854),
            .I(bfn_11_29_0_));
    InMux I__8212 (
            .O(N__40851),
            .I(N__40848));
    LocalMux I__8211 (
            .O(N__40848),
            .I(n25_adj_696));
    InMux I__8210 (
            .O(N__40845),
            .I(n13087));
    InMux I__8209 (
            .O(N__40842),
            .I(N__40839));
    LocalMux I__8208 (
            .O(N__40839),
            .I(n24_adj_695));
    InMux I__8207 (
            .O(N__40836),
            .I(n13088));
    InMux I__8206 (
            .O(N__40833),
            .I(N__40830));
    LocalMux I__8205 (
            .O(N__40830),
            .I(N__40827));
    Span4Mux_v I__8204 (
            .O(N__40827),
            .I(N__40824));
    Odrv4 I__8203 (
            .O(N__40824),
            .I(encoder0_position_scaled_10));
    InMux I__8202 (
            .O(N__40821),
            .I(N__40818));
    LocalMux I__8201 (
            .O(N__40818),
            .I(N__40815));
    Span4Mux_v I__8200 (
            .O(N__40815),
            .I(N__40812));
    Odrv4 I__8199 (
            .O(N__40812),
            .I(pwm_setpoint_23_N_171_3));
    InMux I__8198 (
            .O(N__40809),
            .I(N__40806));
    LocalMux I__8197 (
            .O(N__40806),
            .I(N__40803));
    Span4Mux_h I__8196 (
            .O(N__40803),
            .I(N__40800));
    Odrv4 I__8195 (
            .O(N__40800),
            .I(encoder0_position_scaled_11));
    InMux I__8194 (
            .O(N__40797),
            .I(N__40794));
    LocalMux I__8193 (
            .O(N__40794),
            .I(N__40791));
    Span4Mux_h I__8192 (
            .O(N__40791),
            .I(N__40788));
    Odrv4 I__8191 (
            .O(N__40788),
            .I(pwm_setpoint_23_N_171_13));
    CascadeMux I__8190 (
            .O(N__40785),
            .I(n15_adj_663_cascade_));
    InMux I__8189 (
            .O(N__40782),
            .I(N__40779));
    LocalMux I__8188 (
            .O(N__40779),
            .I(n15125));
    InMux I__8187 (
            .O(N__40776),
            .I(N__40773));
    LocalMux I__8186 (
            .O(N__40773),
            .I(N__40770));
    Span4Mux_v I__8185 (
            .O(N__40770),
            .I(N__40767));
    Odrv4 I__8184 (
            .O(N__40767),
            .I(encoder0_position_scaled_18));
    InMux I__8183 (
            .O(N__40764),
            .I(N__40761));
    LocalMux I__8182 (
            .O(N__40761),
            .I(N__40758));
    Span4Mux_h I__8181 (
            .O(N__40758),
            .I(N__40755));
    Odrv4 I__8180 (
            .O(N__40755),
            .I(encoder0_position_scaled_20));
    InMux I__8179 (
            .O(N__40752),
            .I(N__40749));
    LocalMux I__8178 (
            .O(N__40749),
            .I(N__40746));
    Span4Mux_h I__8177 (
            .O(N__40746),
            .I(N__40743));
    Odrv4 I__8176 (
            .O(N__40743),
            .I(encoder0_position_scaled_23));
    InMux I__8175 (
            .O(N__40740),
            .I(N__40737));
    LocalMux I__8174 (
            .O(N__40737),
            .I(N__40732));
    InMux I__8173 (
            .O(N__40736),
            .I(N__40729));
    InMux I__8172 (
            .O(N__40735),
            .I(N__40725));
    Span4Mux_h I__8171 (
            .O(N__40732),
            .I(N__40722));
    LocalMux I__8170 (
            .O(N__40729),
            .I(N__40719));
    InMux I__8169 (
            .O(N__40728),
            .I(N__40716));
    LocalMux I__8168 (
            .O(N__40725),
            .I(encoder0_position_29));
    Odrv4 I__8167 (
            .O(N__40722),
            .I(encoder0_position_29));
    Odrv4 I__8166 (
            .O(N__40719),
            .I(encoder0_position_29));
    LocalMux I__8165 (
            .O(N__40716),
            .I(encoder0_position_29));
    CascadeMux I__8164 (
            .O(N__40707),
            .I(N__40702));
    InMux I__8163 (
            .O(N__40706),
            .I(N__40699));
    InMux I__8162 (
            .O(N__40705),
            .I(N__40694));
    InMux I__8161 (
            .O(N__40702),
            .I(N__40694));
    LocalMux I__8160 (
            .O(N__40699),
            .I(n4));
    LocalMux I__8159 (
            .O(N__40694),
            .I(n4));
    CascadeMux I__8158 (
            .O(N__40689),
            .I(N__40685));
    CascadeMux I__8157 (
            .O(N__40688),
            .I(N__40681));
    InMux I__8156 (
            .O(N__40685),
            .I(N__40675));
    InMux I__8155 (
            .O(N__40684),
            .I(N__40675));
    InMux I__8154 (
            .O(N__40681),
            .I(N__40670));
    InMux I__8153 (
            .O(N__40680),
            .I(N__40670));
    LocalMux I__8152 (
            .O(N__40675),
            .I(n3));
    LocalMux I__8151 (
            .O(N__40670),
            .I(n3));
    CascadeMux I__8150 (
            .O(N__40665),
            .I(N__40660));
    InMux I__8149 (
            .O(N__40664),
            .I(N__40657));
    CascadeMux I__8148 (
            .O(N__40663),
            .I(N__40654));
    InMux I__8147 (
            .O(N__40660),
            .I(N__40650));
    LocalMux I__8146 (
            .O(N__40657),
            .I(N__40647));
    InMux I__8145 (
            .O(N__40654),
            .I(N__40644));
    InMux I__8144 (
            .O(N__40653),
            .I(N__40641));
    LocalMux I__8143 (
            .O(N__40650),
            .I(encoder0_position_30));
    Odrv12 I__8142 (
            .O(N__40647),
            .I(encoder0_position_30));
    LocalMux I__8141 (
            .O(N__40644),
            .I(encoder0_position_30));
    LocalMux I__8140 (
            .O(N__40641),
            .I(encoder0_position_30));
    CascadeMux I__8139 (
            .O(N__40632),
            .I(n13642_cascade_));
    CascadeMux I__8138 (
            .O(N__40629),
            .I(N__40625));
    InMux I__8137 (
            .O(N__40628),
            .I(N__40622));
    InMux I__8136 (
            .O(N__40625),
            .I(N__40619));
    LocalMux I__8135 (
            .O(N__40622),
            .I(N__40615));
    LocalMux I__8134 (
            .O(N__40619),
            .I(N__40612));
    InMux I__8133 (
            .O(N__40618),
            .I(N__40609));
    Odrv4 I__8132 (
            .O(N__40615),
            .I(n829));
    Odrv12 I__8131 (
            .O(N__40612),
            .I(n829));
    LocalMux I__8130 (
            .O(N__40609),
            .I(n829));
    InMux I__8129 (
            .O(N__40602),
            .I(N__40599));
    LocalMux I__8128 (
            .O(N__40599),
            .I(N__40596));
    Span4Mux_v I__8127 (
            .O(N__40596),
            .I(N__40593));
    Odrv4 I__8126 (
            .O(N__40593),
            .I(n32));
    InMux I__8125 (
            .O(N__40590),
            .I(N__40586));
    CascadeMux I__8124 (
            .O(N__40589),
            .I(N__40583));
    LocalMux I__8123 (
            .O(N__40586),
            .I(N__40580));
    InMux I__8122 (
            .O(N__40583),
            .I(N__40576));
    Span4Mux_v I__8121 (
            .O(N__40580),
            .I(N__40573));
    InMux I__8120 (
            .O(N__40579),
            .I(N__40570));
    LocalMux I__8119 (
            .O(N__40576),
            .I(encoder0_position_1));
    Odrv4 I__8118 (
            .O(N__40573),
            .I(encoder0_position_1));
    LocalMux I__8117 (
            .O(N__40570),
            .I(encoder0_position_1));
    CascadeMux I__8116 (
            .O(N__40563),
            .I(N__40560));
    InMux I__8115 (
            .O(N__40560),
            .I(N__40555));
    InMux I__8114 (
            .O(N__40559),
            .I(N__40552));
    InMux I__8113 (
            .O(N__40558),
            .I(N__40549));
    LocalMux I__8112 (
            .O(N__40555),
            .I(N__40546));
    LocalMux I__8111 (
            .O(N__40552),
            .I(N__40541));
    LocalMux I__8110 (
            .O(N__40549),
            .I(N__40541));
    Span4Mux_v I__8109 (
            .O(N__40546),
            .I(N__40538));
    Span4Mux_v I__8108 (
            .O(N__40541),
            .I(N__40535));
    Span4Mux_h I__8107 (
            .O(N__40538),
            .I(N__40532));
    Span4Mux_h I__8106 (
            .O(N__40535),
            .I(N__40529));
    Odrv4 I__8105 (
            .O(N__40532),
            .I(n318));
    Odrv4 I__8104 (
            .O(N__40529),
            .I(n318));
    InMux I__8103 (
            .O(N__40524),
            .I(N__40521));
    LocalMux I__8102 (
            .O(N__40521),
            .I(N__40518));
    Span4Mux_h I__8101 (
            .O(N__40518),
            .I(N__40515));
    Odrv4 I__8100 (
            .O(N__40515),
            .I(encoder0_position_scaled_14));
    CascadeMux I__8099 (
            .O(N__40512),
            .I(n10_adj_606_cascade_));
    CascadeMux I__8098 (
            .O(N__40509),
            .I(n15_adj_565_cascade_));
    InMux I__8097 (
            .O(N__40506),
            .I(N__40503));
    LocalMux I__8096 (
            .O(N__40503),
            .I(n16_adj_564));
    CascadeMux I__8095 (
            .O(N__40500),
            .I(n13644_cascade_));
    CascadeMux I__8094 (
            .O(N__40497),
            .I(N__40494));
    InMux I__8093 (
            .O(N__40494),
            .I(N__40490));
    InMux I__8092 (
            .O(N__40493),
            .I(N__40486));
    LocalMux I__8091 (
            .O(N__40490),
            .I(N__40483));
    InMux I__8090 (
            .O(N__40489),
            .I(N__40480));
    LocalMux I__8089 (
            .O(N__40486),
            .I(n830));
    Odrv4 I__8088 (
            .O(N__40483),
            .I(n830));
    LocalMux I__8087 (
            .O(N__40480),
            .I(n830));
    InMux I__8086 (
            .O(N__40473),
            .I(N__40467));
    InMux I__8085 (
            .O(N__40472),
            .I(N__40467));
    LocalMux I__8084 (
            .O(N__40467),
            .I(n7));
    InMux I__8083 (
            .O(N__40464),
            .I(N__40461));
    LocalMux I__8082 (
            .O(N__40461),
            .I(n5_adj_676));
    CascadeMux I__8081 (
            .O(N__40458),
            .I(n5_adj_676_cascade_));
    CascadeMux I__8080 (
            .O(N__40455),
            .I(n13641_cascade_));
    CascadeMux I__8079 (
            .O(N__40452),
            .I(n13646_cascade_));
    CascadeMux I__8078 (
            .O(N__40449),
            .I(N__40446));
    InMux I__8077 (
            .O(N__40446),
            .I(N__40443));
    LocalMux I__8076 (
            .O(N__40443),
            .I(N__40438));
    InMux I__8075 (
            .O(N__40442),
            .I(N__40433));
    InMux I__8074 (
            .O(N__40441),
            .I(N__40433));
    Odrv4 I__8073 (
            .O(N__40438),
            .I(n831));
    LocalMux I__8072 (
            .O(N__40433),
            .I(n831));
    CascadeMux I__8071 (
            .O(N__40428),
            .I(N__40423));
    InMux I__8070 (
            .O(N__40427),
            .I(N__40420));
    InMux I__8069 (
            .O(N__40426),
            .I(N__40417));
    InMux I__8068 (
            .O(N__40423),
            .I(N__40413));
    LocalMux I__8067 (
            .O(N__40420),
            .I(N__40408));
    LocalMux I__8066 (
            .O(N__40417),
            .I(N__40408));
    InMux I__8065 (
            .O(N__40416),
            .I(N__40405));
    LocalMux I__8064 (
            .O(N__40413),
            .I(encoder0_position_28));
    Odrv4 I__8063 (
            .O(N__40408),
            .I(encoder0_position_28));
    LocalMux I__8062 (
            .O(N__40405),
            .I(encoder0_position_28));
    CascadeMux I__8061 (
            .O(N__40398),
            .I(N__40394));
    InMux I__8060 (
            .O(N__40397),
            .I(N__40386));
    InMux I__8059 (
            .O(N__40394),
            .I(N__40386));
    InMux I__8058 (
            .O(N__40393),
            .I(N__40386));
    LocalMux I__8057 (
            .O(N__40386),
            .I(n5));
    CascadeMux I__8056 (
            .O(N__40383),
            .I(n931_cascade_));
    CascadeMux I__8055 (
            .O(N__40380),
            .I(N__40377));
    InMux I__8054 (
            .O(N__40377),
            .I(N__40374));
    LocalMux I__8053 (
            .O(N__40374),
            .I(n10));
    CascadeMux I__8052 (
            .O(N__40371),
            .I(N__40368));
    InMux I__8051 (
            .O(N__40368),
            .I(N__40365));
    LocalMux I__8050 (
            .O(N__40365),
            .I(n897));
    CascadeMux I__8049 (
            .O(N__40362),
            .I(N__40359));
    InMux I__8048 (
            .O(N__40359),
            .I(N__40356));
    LocalMux I__8047 (
            .O(N__40356),
            .I(N__40352));
    InMux I__8046 (
            .O(N__40355),
            .I(N__40348));
    Span4Mux_h I__8045 (
            .O(N__40352),
            .I(N__40345));
    InMux I__8044 (
            .O(N__40351),
            .I(N__40342));
    LocalMux I__8043 (
            .O(N__40348),
            .I(encoder0_position_25));
    Odrv4 I__8042 (
            .O(N__40345),
            .I(encoder0_position_25));
    LocalMux I__8041 (
            .O(N__40342),
            .I(encoder0_position_25));
    InMux I__8040 (
            .O(N__40335),
            .I(N__40332));
    LocalMux I__8039 (
            .O(N__40332),
            .I(n8));
    CascadeMux I__8038 (
            .O(N__40329),
            .I(N__40324));
    InMux I__8037 (
            .O(N__40328),
            .I(N__40321));
    InMux I__8036 (
            .O(N__40327),
            .I(N__40318));
    InMux I__8035 (
            .O(N__40324),
            .I(N__40315));
    LocalMux I__8034 (
            .O(N__40321),
            .I(N__40312));
    LocalMux I__8033 (
            .O(N__40318),
            .I(n294));
    LocalMux I__8032 (
            .O(N__40315),
            .I(n294));
    Odrv4 I__8031 (
            .O(N__40312),
            .I(n294));
    CascadeMux I__8030 (
            .O(N__40305),
            .I(N__40302));
    InMux I__8029 (
            .O(N__40302),
            .I(N__40299));
    LocalMux I__8028 (
            .O(N__40299),
            .I(n14574));
    CascadeMux I__8027 (
            .O(N__40296),
            .I(N__40293));
    InMux I__8026 (
            .O(N__40293),
            .I(N__40290));
    LocalMux I__8025 (
            .O(N__40290),
            .I(N__40287));
    Odrv4 I__8024 (
            .O(N__40287),
            .I(n828));
    CascadeMux I__8023 (
            .O(N__40284),
            .I(n828_cascade_));
    InMux I__8022 (
            .O(N__40281),
            .I(N__40278));
    LocalMux I__8021 (
            .O(N__40278),
            .I(n12012));
    InMux I__8020 (
            .O(N__40275),
            .I(N__40270));
    CascadeMux I__8019 (
            .O(N__40274),
            .I(N__40267));
    CascadeMux I__8018 (
            .O(N__40273),
            .I(N__40264));
    LocalMux I__8017 (
            .O(N__40270),
            .I(N__40258));
    InMux I__8016 (
            .O(N__40267),
            .I(N__40247));
    InMux I__8015 (
            .O(N__40264),
            .I(N__40247));
    InMux I__8014 (
            .O(N__40263),
            .I(N__40247));
    InMux I__8013 (
            .O(N__40262),
            .I(N__40247));
    InMux I__8012 (
            .O(N__40261),
            .I(N__40247));
    Odrv4 I__8011 (
            .O(N__40258),
            .I(n861));
    LocalMux I__8010 (
            .O(N__40247),
            .I(n861));
    CascadeMux I__8009 (
            .O(N__40242),
            .I(n861_cascade_));
    InMux I__8008 (
            .O(N__40239),
            .I(N__40236));
    LocalMux I__8007 (
            .O(N__40236),
            .I(N__40233));
    Odrv4 I__8006 (
            .O(N__40233),
            .I(n898));
    InMux I__8005 (
            .O(N__40230),
            .I(n12487));
    InMux I__8004 (
            .O(N__40227),
            .I(n12488));
    InMux I__8003 (
            .O(N__40224),
            .I(n12489));
    InMux I__8002 (
            .O(N__40221),
            .I(n12490));
    InMux I__8001 (
            .O(N__40218),
            .I(n12491));
    InMux I__8000 (
            .O(N__40215),
            .I(n12492));
    CascadeMux I__7999 (
            .O(N__40212),
            .I(N__40209));
    InMux I__7998 (
            .O(N__40209),
            .I(N__40206));
    LocalMux I__7997 (
            .O(N__40206),
            .I(N__40203));
    Odrv12 I__7996 (
            .O(N__40203),
            .I(n901));
    InMux I__7995 (
            .O(N__40200),
            .I(N__40197));
    LocalMux I__7994 (
            .O(N__40197),
            .I(n896));
    CascadeMux I__7993 (
            .O(N__40194),
            .I(N__40191));
    InMux I__7992 (
            .O(N__40191),
            .I(N__40188));
    LocalMux I__7991 (
            .O(N__40188),
            .I(n900));
    InMux I__7990 (
            .O(N__40185),
            .I(N__40182));
    LocalMux I__7989 (
            .O(N__40182),
            .I(n899));
    CascadeMux I__7988 (
            .O(N__40179),
            .I(n1820_cascade_));
    InMux I__7987 (
            .O(N__40176),
            .I(N__40173));
    LocalMux I__7986 (
            .O(N__40173),
            .I(N__40170));
    Odrv4 I__7985 (
            .O(N__40170),
            .I(n14538));
    CascadeMux I__7984 (
            .O(N__40167),
            .I(N__40164));
    InMux I__7983 (
            .O(N__40164),
            .I(N__40161));
    LocalMux I__7982 (
            .O(N__40161),
            .I(n30_adj_651));
    InMux I__7981 (
            .O(N__40158),
            .I(N__40155));
    LocalMux I__7980 (
            .O(N__40155),
            .I(n26));
    InMux I__7979 (
            .O(N__40152),
            .I(N__40148));
    CascadeMux I__7978 (
            .O(N__40151),
            .I(N__40145));
    LocalMux I__7977 (
            .O(N__40148),
            .I(N__40142));
    InMux I__7976 (
            .O(N__40145),
            .I(N__40138));
    Span4Mux_h I__7975 (
            .O(N__40142),
            .I(N__40135));
    InMux I__7974 (
            .O(N__40141),
            .I(N__40132));
    LocalMux I__7973 (
            .O(N__40138),
            .I(encoder0_position_7));
    Odrv4 I__7972 (
            .O(N__40135),
            .I(encoder0_position_7));
    LocalMux I__7971 (
            .O(N__40132),
            .I(encoder0_position_7));
    InMux I__7970 (
            .O(N__40125),
            .I(N__40122));
    LocalMux I__7969 (
            .O(N__40122),
            .I(N__40118));
    InMux I__7968 (
            .O(N__40121),
            .I(N__40114));
    Span4Mux_v I__7967 (
            .O(N__40118),
            .I(N__40111));
    InMux I__7966 (
            .O(N__40117),
            .I(N__40108));
    LocalMux I__7965 (
            .O(N__40114),
            .I(N__40105));
    Span4Mux_v I__7964 (
            .O(N__40111),
            .I(N__40100));
    LocalMux I__7963 (
            .O(N__40108),
            .I(N__40100));
    Span4Mux_h I__7962 (
            .O(N__40105),
            .I(N__40097));
    Span4Mux_h I__7961 (
            .O(N__40100),
            .I(N__40094));
    Span4Mux_h I__7960 (
            .O(N__40097),
            .I(N__40091));
    Odrv4 I__7959 (
            .O(N__40094),
            .I(n312));
    Odrv4 I__7958 (
            .O(N__40091),
            .I(n312));
    InMux I__7957 (
            .O(N__40086),
            .I(N__40083));
    LocalMux I__7956 (
            .O(N__40083),
            .I(n31));
    InMux I__7955 (
            .O(N__40080),
            .I(N__40077));
    LocalMux I__7954 (
            .O(N__40077),
            .I(N__40073));
    InMux I__7953 (
            .O(N__40076),
            .I(N__40069));
    Span4Mux_h I__7952 (
            .O(N__40073),
            .I(N__40066));
    InMux I__7951 (
            .O(N__40072),
            .I(N__40063));
    LocalMux I__7950 (
            .O(N__40069),
            .I(encoder0_position_2));
    Odrv4 I__7949 (
            .O(N__40066),
            .I(encoder0_position_2));
    LocalMux I__7948 (
            .O(N__40063),
            .I(encoder0_position_2));
    InMux I__7947 (
            .O(N__40056),
            .I(N__40051));
    InMux I__7946 (
            .O(N__40055),
            .I(N__40048));
    InMux I__7945 (
            .O(N__40054),
            .I(N__40045));
    LocalMux I__7944 (
            .O(N__40051),
            .I(N__40042));
    LocalMux I__7943 (
            .O(N__40048),
            .I(N__40039));
    LocalMux I__7942 (
            .O(N__40045),
            .I(N__40036));
    Span4Mux_h I__7941 (
            .O(N__40042),
            .I(N__40033));
    Span4Mux_v I__7940 (
            .O(N__40039),
            .I(N__40030));
    Span4Mux_h I__7939 (
            .O(N__40036),
            .I(N__40027));
    Span4Mux_v I__7938 (
            .O(N__40033),
            .I(N__40024));
    Span4Mux_h I__7937 (
            .O(N__40030),
            .I(N__40021));
    Span4Mux_v I__7936 (
            .O(N__40027),
            .I(N__40018));
    Sp12to4 I__7935 (
            .O(N__40024),
            .I(N__40015));
    Odrv4 I__7934 (
            .O(N__40021),
            .I(n317));
    Odrv4 I__7933 (
            .O(N__40018),
            .I(n317));
    Odrv12 I__7932 (
            .O(N__40015),
            .I(n317));
    CascadeMux I__7931 (
            .O(N__40008),
            .I(N__40003));
    InMux I__7930 (
            .O(N__40007),
            .I(N__40000));
    InMux I__7929 (
            .O(N__40006),
            .I(N__39997));
    InMux I__7928 (
            .O(N__40003),
            .I(N__39994));
    LocalMux I__7927 (
            .O(N__40000),
            .I(N__39991));
    LocalMux I__7926 (
            .O(N__39997),
            .I(N__39988));
    LocalMux I__7925 (
            .O(N__39994),
            .I(N__39981));
    Span4Mux_h I__7924 (
            .O(N__39991),
            .I(N__39981));
    Span4Mux_v I__7923 (
            .O(N__39988),
            .I(N__39981));
    Odrv4 I__7922 (
            .O(N__39981),
            .I(encoder0_position_10));
    CascadeMux I__7921 (
            .O(N__39978),
            .I(N__39975));
    InMux I__7920 (
            .O(N__39975),
            .I(N__39972));
    LocalMux I__7919 (
            .O(N__39972),
            .I(n23_adj_644));
    InMux I__7918 (
            .O(N__39969),
            .I(N__39966));
    LocalMux I__7917 (
            .O(N__39966),
            .I(N__39963));
    Span4Mux_h I__7916 (
            .O(N__39963),
            .I(N__39960));
    Odrv4 I__7915 (
            .O(N__39960),
            .I(encoder0_position_scaled_1));
    InMux I__7914 (
            .O(N__39957),
            .I(bfn_11_22_0_));
    CascadeMux I__7913 (
            .O(N__39954),
            .I(N__39951));
    InMux I__7912 (
            .O(N__39951),
            .I(N__39947));
    InMux I__7911 (
            .O(N__39950),
            .I(N__39943));
    LocalMux I__7910 (
            .O(N__39947),
            .I(N__39940));
    InMux I__7909 (
            .O(N__39946),
            .I(N__39937));
    LocalMux I__7908 (
            .O(N__39943),
            .I(N__39932));
    Span4Mux_v I__7907 (
            .O(N__39940),
            .I(N__39932));
    LocalMux I__7906 (
            .O(N__39937),
            .I(n1931));
    Odrv4 I__7905 (
            .O(N__39932),
            .I(n1931));
    CascadeMux I__7904 (
            .O(N__39927),
            .I(N__39923));
    CascadeMux I__7903 (
            .O(N__39926),
            .I(N__39920));
    InMux I__7902 (
            .O(N__39923),
            .I(N__39915));
    InMux I__7901 (
            .O(N__39920),
            .I(N__39915));
    LocalMux I__7900 (
            .O(N__39915),
            .I(N__39911));
    InMux I__7899 (
            .O(N__39914),
            .I(N__39908));
    Odrv4 I__7898 (
            .O(N__39911),
            .I(n1918));
    LocalMux I__7897 (
            .O(N__39908),
            .I(n1918));
    CascadeMux I__7896 (
            .O(N__39903),
            .I(N__39900));
    InMux I__7895 (
            .O(N__39900),
            .I(N__39897));
    LocalMux I__7894 (
            .O(N__39897),
            .I(n14520));
    CascadeMux I__7893 (
            .O(N__39894),
            .I(n14176_cascade_));
    CascadeMux I__7892 (
            .O(N__39891),
            .I(n1752_cascade_));
    InMux I__7891 (
            .O(N__39888),
            .I(N__39885));
    LocalMux I__7890 (
            .O(N__39885),
            .I(N__39878));
    CascadeMux I__7889 (
            .O(N__39884),
            .I(N__39875));
    InMux I__7888 (
            .O(N__39883),
            .I(N__39869));
    CascadeMux I__7887 (
            .O(N__39882),
            .I(N__39864));
    CascadeMux I__7886 (
            .O(N__39881),
            .I(N__39861));
    Span4Mux_v I__7885 (
            .O(N__39878),
            .I(N__39856));
    InMux I__7884 (
            .O(N__39875),
            .I(N__39853));
    CascadeMux I__7883 (
            .O(N__39874),
            .I(N__39849));
    CascadeMux I__7882 (
            .O(N__39873),
            .I(N__39846));
    CascadeMux I__7881 (
            .O(N__39872),
            .I(N__39842));
    LocalMux I__7880 (
            .O(N__39869),
            .I(N__39835));
    InMux I__7879 (
            .O(N__39868),
            .I(N__39830));
    InMux I__7878 (
            .O(N__39867),
            .I(N__39830));
    InMux I__7877 (
            .O(N__39864),
            .I(N__39821));
    InMux I__7876 (
            .O(N__39861),
            .I(N__39821));
    InMux I__7875 (
            .O(N__39860),
            .I(N__39821));
    InMux I__7874 (
            .O(N__39859),
            .I(N__39821));
    Span4Mux_h I__7873 (
            .O(N__39856),
            .I(N__39816));
    LocalMux I__7872 (
            .O(N__39853),
            .I(N__39816));
    InMux I__7871 (
            .O(N__39852),
            .I(N__39807));
    InMux I__7870 (
            .O(N__39849),
            .I(N__39807));
    InMux I__7869 (
            .O(N__39846),
            .I(N__39807));
    InMux I__7868 (
            .O(N__39845),
            .I(N__39807));
    InMux I__7867 (
            .O(N__39842),
            .I(N__39802));
    InMux I__7866 (
            .O(N__39841),
            .I(N__39802));
    InMux I__7865 (
            .O(N__39840),
            .I(N__39795));
    InMux I__7864 (
            .O(N__39839),
            .I(N__39795));
    InMux I__7863 (
            .O(N__39838),
            .I(N__39795));
    Odrv12 I__7862 (
            .O(N__39835),
            .I(n1851));
    LocalMux I__7861 (
            .O(N__39830),
            .I(n1851));
    LocalMux I__7860 (
            .O(N__39821),
            .I(n1851));
    Odrv4 I__7859 (
            .O(N__39816),
            .I(n1851));
    LocalMux I__7858 (
            .O(N__39807),
            .I(n1851));
    LocalMux I__7857 (
            .O(N__39802),
            .I(n1851));
    LocalMux I__7856 (
            .O(N__39795),
            .I(n1851));
    InMux I__7855 (
            .O(N__39780),
            .I(N__39777));
    LocalMux I__7854 (
            .O(N__39777),
            .I(N__39774));
    Span4Mux_h I__7853 (
            .O(N__39774),
            .I(N__39771));
    Span4Mux_v I__7852 (
            .O(N__39771),
            .I(N__39768));
    Odrv4 I__7851 (
            .O(N__39768),
            .I(n15644));
    CascadeMux I__7850 (
            .O(N__39765),
            .I(n1832_cascade_));
    InMux I__7849 (
            .O(N__39762),
            .I(N__39759));
    LocalMux I__7848 (
            .O(N__39759),
            .I(N__39756));
    Odrv4 I__7847 (
            .O(N__39756),
            .I(n11968));
    CascadeMux I__7846 (
            .O(N__39753),
            .I(n1819_cascade_));
    InMux I__7845 (
            .O(N__39750),
            .I(N__39747));
    LocalMux I__7844 (
            .O(N__39747),
            .I(n14532));
    CascadeMux I__7843 (
            .O(N__39744),
            .I(n1851_cascade_));
    InMux I__7842 (
            .O(N__39741),
            .I(N__39738));
    LocalMux I__7841 (
            .O(N__39738),
            .I(N__39734));
    InMux I__7840 (
            .O(N__39737),
            .I(N__39731));
    Span4Mux_v I__7839 (
            .O(N__39734),
            .I(N__39725));
    LocalMux I__7838 (
            .O(N__39731),
            .I(N__39725));
    InMux I__7837 (
            .O(N__39730),
            .I(N__39722));
    Odrv4 I__7836 (
            .O(N__39725),
            .I(n1920));
    LocalMux I__7835 (
            .O(N__39722),
            .I(n1920));
    InMux I__7834 (
            .O(N__39717),
            .I(N__39713));
    InMux I__7833 (
            .O(N__39716),
            .I(N__39710));
    LocalMux I__7832 (
            .O(N__39713),
            .I(N__39707));
    LocalMux I__7831 (
            .O(N__39710),
            .I(N__39704));
    Span4Mux_h I__7830 (
            .O(N__39707),
            .I(N__39698));
    Span4Mux_v I__7829 (
            .O(N__39704),
            .I(N__39698));
    InMux I__7828 (
            .O(N__39703),
            .I(N__39695));
    Odrv4 I__7827 (
            .O(N__39698),
            .I(n1919));
    LocalMux I__7826 (
            .O(N__39695),
            .I(n1919));
    CascadeMux I__7825 (
            .O(N__39690),
            .I(N__39687));
    InMux I__7824 (
            .O(N__39687),
            .I(N__39683));
    InMux I__7823 (
            .O(N__39686),
            .I(N__39680));
    LocalMux I__7822 (
            .O(N__39683),
            .I(N__39677));
    LocalMux I__7821 (
            .O(N__39680),
            .I(N__39674));
    Span4Mux_h I__7820 (
            .O(N__39677),
            .I(N__39671));
    Odrv4 I__7819 (
            .O(N__39674),
            .I(n1930));
    Odrv4 I__7818 (
            .O(N__39671),
            .I(n1930));
    CascadeMux I__7817 (
            .O(N__39666),
            .I(n1930_cascade_));
    CascadeMux I__7816 (
            .O(N__39663),
            .I(N__39659));
    CascadeMux I__7815 (
            .O(N__39662),
            .I(N__39656));
    InMux I__7814 (
            .O(N__39659),
            .I(N__39653));
    InMux I__7813 (
            .O(N__39656),
            .I(N__39649));
    LocalMux I__7812 (
            .O(N__39653),
            .I(N__39646));
    InMux I__7811 (
            .O(N__39652),
            .I(N__39643));
    LocalMux I__7810 (
            .O(N__39649),
            .I(N__39640));
    Span4Mux_h I__7809 (
            .O(N__39646),
            .I(N__39635));
    LocalMux I__7808 (
            .O(N__39643),
            .I(N__39635));
    Odrv4 I__7807 (
            .O(N__39640),
            .I(n1929));
    Odrv4 I__7806 (
            .O(N__39635),
            .I(n1929));
    CascadeMux I__7805 (
            .O(N__39630),
            .I(N__39627));
    InMux I__7804 (
            .O(N__39627),
            .I(N__39624));
    LocalMux I__7803 (
            .O(N__39624),
            .I(n14540));
    CascadeMux I__7802 (
            .O(N__39621),
            .I(n1826_cascade_));
    CascadeMux I__7801 (
            .O(N__39618),
            .I(N__39614));
    CascadeMux I__7800 (
            .O(N__39617),
            .I(N__39611));
    InMux I__7799 (
            .O(N__39614),
            .I(N__39608));
    InMux I__7798 (
            .O(N__39611),
            .I(N__39604));
    LocalMux I__7797 (
            .O(N__39608),
            .I(N__39601));
    InMux I__7796 (
            .O(N__39607),
            .I(N__39598));
    LocalMux I__7795 (
            .O(N__39604),
            .I(n1928));
    Odrv4 I__7794 (
            .O(N__39601),
            .I(n1928));
    LocalMux I__7793 (
            .O(N__39598),
            .I(n1928));
    InMux I__7792 (
            .O(N__39591),
            .I(N__39588));
    LocalMux I__7791 (
            .O(N__39588),
            .I(n14526));
    CascadeMux I__7790 (
            .O(N__39585),
            .I(n14530_cascade_));
    InMux I__7789 (
            .O(N__39582),
            .I(N__39579));
    LocalMux I__7788 (
            .O(N__39579),
            .I(n11_adj_591));
    InMux I__7787 (
            .O(N__39576),
            .I(N__39573));
    LocalMux I__7786 (
            .O(N__39573),
            .I(pwm_setpoint_23_N_171_18));
    InMux I__7785 (
            .O(N__39570),
            .I(N__39567));
    LocalMux I__7784 (
            .O(N__39567),
            .I(n3_adj_583));
    InMux I__7783 (
            .O(N__39564),
            .I(N__39561));
    LocalMux I__7782 (
            .O(N__39561),
            .I(n9_adj_589));
    InMux I__7781 (
            .O(N__39558),
            .I(N__39555));
    LocalMux I__7780 (
            .O(N__39555),
            .I(N__39551));
    InMux I__7779 (
            .O(N__39554),
            .I(N__39548));
    Odrv12 I__7778 (
            .O(N__39551),
            .I(reg_B_2));
    LocalMux I__7777 (
            .O(N__39548),
            .I(reg_B_2));
    InMux I__7776 (
            .O(N__39543),
            .I(N__39540));
    LocalMux I__7775 (
            .O(N__39540),
            .I(N__39536));
    InMux I__7774 (
            .O(N__39539),
            .I(N__39533));
    Span4Mux_s2_h I__7773 (
            .O(N__39536),
            .I(N__39530));
    LocalMux I__7772 (
            .O(N__39533),
            .I(N__39527));
    Span4Mux_v I__7771 (
            .O(N__39530),
            .I(N__39523));
    Span4Mux_v I__7770 (
            .O(N__39527),
            .I(N__39520));
    InMux I__7769 (
            .O(N__39526),
            .I(N__39517));
    Span4Mux_v I__7768 (
            .O(N__39523),
            .I(N__39513));
    Sp12to4 I__7767 (
            .O(N__39520),
            .I(N__39508));
    LocalMux I__7766 (
            .O(N__39517),
            .I(N__39508));
    InMux I__7765 (
            .O(N__39516),
            .I(N__39505));
    Odrv4 I__7764 (
            .O(N__39513),
            .I(n14125));
    Odrv12 I__7763 (
            .O(N__39508),
            .I(n14125));
    LocalMux I__7762 (
            .O(N__39505),
            .I(n14125));
    InMux I__7761 (
            .O(N__39498),
            .I(N__39495));
    LocalMux I__7760 (
            .O(N__39495),
            .I(n14937));
    CascadeMux I__7759 (
            .O(N__39492),
            .I(n14936_cascade_));
    IoInMux I__7758 (
            .O(N__39489),
            .I(N__39486));
    LocalMux I__7757 (
            .O(N__39486),
            .I(N__39483));
    Span4Mux_s0_v I__7756 (
            .O(N__39483),
            .I(N__39480));
    Span4Mux_h I__7755 (
            .O(N__39480),
            .I(N__39477));
    Odrv4 I__7754 (
            .O(N__39477),
            .I(LED_c));
    InMux I__7753 (
            .O(N__39474),
            .I(N__39471));
    LocalMux I__7752 (
            .O(N__39471),
            .I(pwm_setpoint_23_N_171_22));
    InMux I__7751 (
            .O(N__39468),
            .I(N__39465));
    LocalMux I__7750 (
            .O(N__39465),
            .I(n19_adj_599));
    InMux I__7749 (
            .O(N__39462),
            .I(N__39459));
    LocalMux I__7748 (
            .O(N__39459),
            .I(pwm_setpoint_23_N_171_6));
    InMux I__7747 (
            .O(N__39456),
            .I(N__39453));
    LocalMux I__7746 (
            .O(N__39453),
            .I(pwm_setpoint_23_N_171_10));
    InMux I__7745 (
            .O(N__39450),
            .I(N__39447));
    LocalMux I__7744 (
            .O(N__39447),
            .I(pwm_setpoint_23_N_171_9));
    InMux I__7743 (
            .O(N__39444),
            .I(N__39441));
    LocalMux I__7742 (
            .O(N__39441),
            .I(pwm_setpoint_23_N_171_4));
    InMux I__7741 (
            .O(N__39438),
            .I(N__39435));
    LocalMux I__7740 (
            .O(N__39435),
            .I(n7_adj_587));
    InMux I__7739 (
            .O(N__39432),
            .I(N__39429));
    LocalMux I__7738 (
            .O(N__39429),
            .I(pwm_setpoint_23_N_171_15));
    InMux I__7737 (
            .O(N__39426),
            .I(N__39422));
    InMux I__7736 (
            .O(N__39425),
            .I(N__39419));
    LocalMux I__7735 (
            .O(N__39422),
            .I(N__39416));
    LocalMux I__7734 (
            .O(N__39419),
            .I(N__39413));
    Span4Mux_v I__7733 (
            .O(N__39416),
            .I(N__39410));
    Span12Mux_s3_v I__7732 (
            .O(N__39413),
            .I(N__39407));
    Span4Mux_h I__7731 (
            .O(N__39410),
            .I(N__39404));
    Odrv12 I__7730 (
            .O(N__39407),
            .I(reg_B_1));
    Odrv4 I__7729 (
            .O(N__39404),
            .I(reg_B_1));
    InMux I__7728 (
            .O(N__39399),
            .I(N__39396));
    LocalMux I__7727 (
            .O(N__39396),
            .I(N__39392));
    InMux I__7726 (
            .O(N__39395),
            .I(N__39389));
    Odrv4 I__7725 (
            .O(N__39392),
            .I(pwm_setpoint_15));
    LocalMux I__7724 (
            .O(N__39389),
            .I(pwm_setpoint_15));
    InMux I__7723 (
            .O(N__39384),
            .I(N__39379));
    InMux I__7722 (
            .O(N__39383),
            .I(N__39374));
    InMux I__7721 (
            .O(N__39382),
            .I(N__39374));
    LocalMux I__7720 (
            .O(N__39379),
            .I(N__39369));
    LocalMux I__7719 (
            .O(N__39374),
            .I(N__39369));
    Odrv12 I__7718 (
            .O(N__39369),
            .I(n31_adj_674));
    InMux I__7717 (
            .O(N__39366),
            .I(N__39363));
    LocalMux I__7716 (
            .O(N__39363),
            .I(n15121));
    InMux I__7715 (
            .O(N__39360),
            .I(N__39357));
    LocalMux I__7714 (
            .O(N__39357),
            .I(n15182));
    InMux I__7713 (
            .O(N__39354),
            .I(N__39351));
    LocalMux I__7712 (
            .O(N__39351),
            .I(N__39347));
    InMux I__7711 (
            .O(N__39350),
            .I(N__39344));
    Odrv4 I__7710 (
            .O(N__39347),
            .I(n29_adj_672));
    LocalMux I__7709 (
            .O(N__39344),
            .I(n29_adj_672));
    CascadeMux I__7708 (
            .O(N__39339),
            .I(n30_adj_673_cascade_));
    InMux I__7707 (
            .O(N__39336),
            .I(N__39333));
    LocalMux I__7706 (
            .O(N__39333),
            .I(n10_adj_659));
    CascadeMux I__7705 (
            .O(N__39330),
            .I(N__39327));
    InMux I__7704 (
            .O(N__39327),
            .I(N__39324));
    LocalMux I__7703 (
            .O(N__39324),
            .I(n15267));
    InMux I__7702 (
            .O(N__39321),
            .I(N__39318));
    LocalMux I__7701 (
            .O(N__39318),
            .I(n20_adj_600));
    InMux I__7700 (
            .O(N__39315),
            .I(N__39312));
    LocalMux I__7699 (
            .O(N__39312),
            .I(n16_adj_596));
    InMux I__7698 (
            .O(N__39309),
            .I(N__39306));
    LocalMux I__7697 (
            .O(N__39306),
            .I(n15_adj_595));
    InMux I__7696 (
            .O(N__39303),
            .I(N__39300));
    LocalMux I__7695 (
            .O(N__39300),
            .I(n21_adj_601));
    InMux I__7694 (
            .O(N__39297),
            .I(N__39294));
    LocalMux I__7693 (
            .O(N__39294),
            .I(pwm_setpoint_23_N_171_5));
    CascadeMux I__7692 (
            .O(N__39291),
            .I(n29_adj_672_cascade_));
    InMux I__7691 (
            .O(N__39288),
            .I(N__39285));
    LocalMux I__7690 (
            .O(N__39285),
            .I(n15233));
    InMux I__7689 (
            .O(N__39282),
            .I(N__39279));
    LocalMux I__7688 (
            .O(N__39279),
            .I(n15234));
    InMux I__7687 (
            .O(N__39276),
            .I(N__39273));
    LocalMux I__7686 (
            .O(N__39273),
            .I(N__39270));
    Span4Mux_v I__7685 (
            .O(N__39270),
            .I(N__39267));
    Odrv4 I__7684 (
            .O(N__39267),
            .I(encoder0_position_scaled_16));
    CascadeMux I__7683 (
            .O(N__39264),
            .I(n33_adj_675_cascade_));
    InMux I__7682 (
            .O(N__39261),
            .I(N__39258));
    LocalMux I__7681 (
            .O(N__39258),
            .I(N__39255));
    Odrv4 I__7680 (
            .O(N__39255),
            .I(n12_adj_592));
    InMux I__7679 (
            .O(N__39252),
            .I(N__39249));
    LocalMux I__7678 (
            .O(N__39249),
            .I(N__39246));
    Span4Mux_h I__7677 (
            .O(N__39246),
            .I(N__39243));
    Odrv4 I__7676 (
            .O(N__39243),
            .I(pwm_setpoint_23_N_171_16));
    CascadeMux I__7675 (
            .O(N__39240),
            .I(N__39237));
    InMux I__7674 (
            .O(N__39237),
            .I(N__39234));
    LocalMux I__7673 (
            .O(N__39234),
            .I(N__39231));
    Odrv4 I__7672 (
            .O(N__39231),
            .I(pwm_setpoint_23_N_171_2));
    CascadeMux I__7671 (
            .O(N__39228),
            .I(N__39225));
    InMux I__7670 (
            .O(N__39225),
            .I(N__39222));
    LocalMux I__7669 (
            .O(N__39222),
            .I(N__39219));
    Span4Mux_v I__7668 (
            .O(N__39219),
            .I(N__39216));
    Odrv4 I__7667 (
            .O(N__39216),
            .I(pwm_setpoint_23_N_171_14));
    InMux I__7666 (
            .O(N__39213),
            .I(N__39207));
    InMux I__7665 (
            .O(N__39212),
            .I(N__39207));
    LocalMux I__7664 (
            .O(N__39207),
            .I(N__39204));
    Odrv4 I__7663 (
            .O(N__39204),
            .I(pwm_setpoint_14));
    CascadeMux I__7662 (
            .O(N__39201),
            .I(N__39198));
    InMux I__7661 (
            .O(N__39198),
            .I(N__39195));
    LocalMux I__7660 (
            .O(N__39195),
            .I(N__39192));
    Odrv4 I__7659 (
            .O(N__39192),
            .I(n3_adj_624));
    InMux I__7658 (
            .O(N__39189),
            .I(N__39186));
    LocalMux I__7657 (
            .O(N__39186),
            .I(N__39183));
    Span4Mux_h I__7656 (
            .O(N__39183),
            .I(N__39180));
    Odrv4 I__7655 (
            .O(N__39180),
            .I(encoder0_position_scaled_2));
    InMux I__7654 (
            .O(N__39177),
            .I(N__39174));
    LocalMux I__7653 (
            .O(N__39174),
            .I(n4_adj_655));
    CascadeMux I__7652 (
            .O(N__39171),
            .I(N__39168));
    InMux I__7651 (
            .O(N__39168),
            .I(N__39165));
    LocalMux I__7650 (
            .O(N__39165),
            .I(\quad_counter0.a_prev_N_543 ));
    InMux I__7649 (
            .O(N__39162),
            .I(N__39152));
    InMux I__7648 (
            .O(N__39161),
            .I(N__39152));
    InMux I__7647 (
            .O(N__39160),
            .I(N__39152));
    InMux I__7646 (
            .O(N__39159),
            .I(N__39149));
    LocalMux I__7645 (
            .O(N__39152),
            .I(\quad_counter0.b_new_1 ));
    LocalMux I__7644 (
            .O(N__39149),
            .I(\quad_counter0.b_new_1 ));
    InMux I__7643 (
            .O(N__39144),
            .I(N__39138));
    InMux I__7642 (
            .O(N__39143),
            .I(N__39138));
    LocalMux I__7641 (
            .O(N__39138),
            .I(\quad_counter0.a_prev ));
    InMux I__7640 (
            .O(N__39135),
            .I(N__39130));
    InMux I__7639 (
            .O(N__39134),
            .I(N__39125));
    InMux I__7638 (
            .O(N__39133),
            .I(N__39125));
    LocalMux I__7637 (
            .O(N__39130),
            .I(\quad_counter0.debounce_cnt ));
    LocalMux I__7636 (
            .O(N__39125),
            .I(\quad_counter0.debounce_cnt ));
    CascadeMux I__7635 (
            .O(N__39120),
            .I(\quad_counter0.direction_N_540_cascade_ ));
    CEMux I__7634 (
            .O(N__39117),
            .I(N__39114));
    LocalMux I__7633 (
            .O(N__39114),
            .I(N__39108));
    CEMux I__7632 (
            .O(N__39113),
            .I(N__39105));
    CEMux I__7631 (
            .O(N__39112),
            .I(N__39102));
    CEMux I__7630 (
            .O(N__39111),
            .I(N__39099));
    Span4Mux_h I__7629 (
            .O(N__39108),
            .I(N__39092));
    LocalMux I__7628 (
            .O(N__39105),
            .I(N__39092));
    LocalMux I__7627 (
            .O(N__39102),
            .I(N__39092));
    LocalMux I__7626 (
            .O(N__39099),
            .I(N__39089));
    Span4Mux_v I__7625 (
            .O(N__39092),
            .I(N__39086));
    Odrv4 I__7624 (
            .O(N__39089),
            .I(direction_N_537));
    Odrv4 I__7623 (
            .O(N__39086),
            .I(direction_N_537));
    CascadeMux I__7622 (
            .O(N__39081),
            .I(N__39077));
    CascadeMux I__7621 (
            .O(N__39080),
            .I(N__39071));
    InMux I__7620 (
            .O(N__39077),
            .I(N__39067));
    InMux I__7619 (
            .O(N__39076),
            .I(N__39060));
    InMux I__7618 (
            .O(N__39075),
            .I(N__39060));
    InMux I__7617 (
            .O(N__39074),
            .I(N__39060));
    InMux I__7616 (
            .O(N__39071),
            .I(N__39055));
    InMux I__7615 (
            .O(N__39070),
            .I(N__39055));
    LocalMux I__7614 (
            .O(N__39067),
            .I(a_new_1));
    LocalMux I__7613 (
            .O(N__39060),
            .I(a_new_1));
    LocalMux I__7612 (
            .O(N__39055),
            .I(a_new_1));
    CascadeMux I__7611 (
            .O(N__39048),
            .I(direction_N_537_cascade_));
    InMux I__7610 (
            .O(N__39045),
            .I(N__39039));
    InMux I__7609 (
            .O(N__39044),
            .I(N__39034));
    InMux I__7608 (
            .O(N__39043),
            .I(N__39034));
    InMux I__7607 (
            .O(N__39042),
            .I(N__39031));
    LocalMux I__7606 (
            .O(N__39039),
            .I(b_prev));
    LocalMux I__7605 (
            .O(N__39034),
            .I(b_prev));
    LocalMux I__7604 (
            .O(N__39031),
            .I(b_prev));
    InMux I__7603 (
            .O(N__39024),
            .I(N__39021));
    LocalMux I__7602 (
            .O(N__39021),
            .I(n1302));
    CascadeMux I__7601 (
            .O(N__39018),
            .I(N__39015));
    InMux I__7600 (
            .O(N__39015),
            .I(N__39012));
    LocalMux I__7599 (
            .O(N__39012),
            .I(n4_adj_625));
    InMux I__7598 (
            .O(N__39009),
            .I(N__39006));
    LocalMux I__7597 (
            .O(N__39006),
            .I(pwm_setpoint_1));
    InMux I__7596 (
            .O(N__39003),
            .I(N__39000));
    LocalMux I__7595 (
            .O(N__39000),
            .I(pwm_setpoint_0));
    InMux I__7594 (
            .O(N__38997),
            .I(N__38994));
    LocalMux I__7593 (
            .O(N__38994),
            .I(N__38991));
    Odrv12 I__7592 (
            .O(N__38991),
            .I(n28));
    InMux I__7591 (
            .O(N__38988),
            .I(N__38984));
    CascadeMux I__7590 (
            .O(N__38987),
            .I(N__38981));
    LocalMux I__7589 (
            .O(N__38984),
            .I(N__38978));
    InMux I__7588 (
            .O(N__38981),
            .I(N__38974));
    Span4Mux_v I__7587 (
            .O(N__38978),
            .I(N__38971));
    InMux I__7586 (
            .O(N__38977),
            .I(N__38968));
    LocalMux I__7585 (
            .O(N__38974),
            .I(encoder0_position_5));
    Odrv4 I__7584 (
            .O(N__38971),
            .I(encoder0_position_5));
    LocalMux I__7583 (
            .O(N__38968),
            .I(encoder0_position_5));
    CascadeMux I__7582 (
            .O(N__38961),
            .I(N__38958));
    InMux I__7581 (
            .O(N__38958),
            .I(N__38953));
    InMux I__7580 (
            .O(N__38957),
            .I(N__38950));
    InMux I__7579 (
            .O(N__38956),
            .I(N__38947));
    LocalMux I__7578 (
            .O(N__38953),
            .I(N__38942));
    LocalMux I__7577 (
            .O(N__38950),
            .I(N__38942));
    LocalMux I__7576 (
            .O(N__38947),
            .I(N__38937));
    Span4Mux_v I__7575 (
            .O(N__38942),
            .I(N__38937));
    Span4Mux_h I__7574 (
            .O(N__38937),
            .I(N__38934));
    Span4Mux_h I__7573 (
            .O(N__38934),
            .I(N__38931));
    Odrv4 I__7572 (
            .O(N__38931),
            .I(n314));
    InMux I__7571 (
            .O(N__38928),
            .I(N__38923));
    InMux I__7570 (
            .O(N__38927),
            .I(N__38920));
    InMux I__7569 (
            .O(N__38926),
            .I(N__38917));
    LocalMux I__7568 (
            .O(N__38923),
            .I(N__38914));
    LocalMux I__7567 (
            .O(N__38920),
            .I(N__38909));
    LocalMux I__7566 (
            .O(N__38917),
            .I(N__38909));
    Span4Mux_v I__7565 (
            .O(N__38914),
            .I(N__38906));
    Span4Mux_h I__7564 (
            .O(N__38909),
            .I(N__38903));
    Span4Mux_h I__7563 (
            .O(N__38906),
            .I(N__38900));
    Span4Mux_h I__7562 (
            .O(N__38903),
            .I(N__38897));
    Odrv4 I__7561 (
            .O(N__38900),
            .I(\quad_counter0.b_new_0 ));
    Odrv4 I__7560 (
            .O(N__38897),
            .I(\quad_counter0.b_new_0 ));
    InMux I__7559 (
            .O(N__38892),
            .I(N__38889));
    LocalMux I__7558 (
            .O(N__38889),
            .I(N__38886));
    Span4Mux_v I__7557 (
            .O(N__38886),
            .I(N__38883));
    Odrv4 I__7556 (
            .O(N__38883),
            .I(encoder0_position_scaled_0));
    InMux I__7555 (
            .O(N__38880),
            .I(N__38877));
    LocalMux I__7554 (
            .O(N__38877),
            .I(N__38874));
    Span4Mux_v I__7553 (
            .O(N__38874),
            .I(N__38871));
    Odrv4 I__7552 (
            .O(N__38871),
            .I(encoder0_position_scaled_15));
    InMux I__7551 (
            .O(N__38868),
            .I(N__38865));
    LocalMux I__7550 (
            .O(N__38865),
            .I(N__38862));
    Span4Mux_h I__7549 (
            .O(N__38862),
            .I(N__38859));
    Odrv4 I__7548 (
            .O(N__38859),
            .I(encoder0_position_scaled_13));
    InMux I__7547 (
            .O(N__38856),
            .I(n12994));
    InMux I__7546 (
            .O(N__38853),
            .I(n12995));
    InMux I__7545 (
            .O(N__38850),
            .I(n12996));
    InMux I__7544 (
            .O(N__38847),
            .I(n12997));
    InMux I__7543 (
            .O(N__38844),
            .I(n12998));
    CascadeMux I__7542 (
            .O(N__38841),
            .I(N__38838));
    InMux I__7541 (
            .O(N__38838),
            .I(N__38835));
    LocalMux I__7540 (
            .O(N__38835),
            .I(n5_adj_626));
    CascadeMux I__7539 (
            .O(N__38832),
            .I(N__38829));
    InMux I__7538 (
            .O(N__38829),
            .I(N__38826));
    LocalMux I__7537 (
            .O(N__38826),
            .I(n6_adj_627));
    CascadeMux I__7536 (
            .O(N__38823),
            .I(N__38820));
    InMux I__7535 (
            .O(N__38820),
            .I(N__38817));
    LocalMux I__7534 (
            .O(N__38817),
            .I(n8_adj_629));
    CascadeMux I__7533 (
            .O(N__38814),
            .I(N__38811));
    InMux I__7532 (
            .O(N__38811),
            .I(N__38808));
    LocalMux I__7531 (
            .O(N__38808),
            .I(n7_adj_628));
    CascadeMux I__7530 (
            .O(N__38805),
            .I(N__38802));
    InMux I__7529 (
            .O(N__38802),
            .I(N__38799));
    LocalMux I__7528 (
            .O(N__38799),
            .I(N__38796));
    Odrv4 I__7527 (
            .O(N__38796),
            .I(n15_adj_636));
    InMux I__7526 (
            .O(N__38793),
            .I(n12985));
    InMux I__7525 (
            .O(N__38790),
            .I(n12986));
    CascadeMux I__7524 (
            .O(N__38787),
            .I(N__38784));
    InMux I__7523 (
            .O(N__38784),
            .I(N__38781));
    LocalMux I__7522 (
            .O(N__38781),
            .I(N__38778));
    Odrv4 I__7521 (
            .O(N__38778),
            .I(n13_adj_634));
    InMux I__7520 (
            .O(N__38775),
            .I(n12987));
    InMux I__7519 (
            .O(N__38772),
            .I(n12988));
    InMux I__7518 (
            .O(N__38769),
            .I(n12989));
    InMux I__7517 (
            .O(N__38766),
            .I(n12990));
    InMux I__7516 (
            .O(N__38763),
            .I(bfn_10_24_0_));
    InMux I__7515 (
            .O(N__38760),
            .I(n12992));
    InMux I__7514 (
            .O(N__38757),
            .I(n12993));
    InMux I__7513 (
            .O(N__38754),
            .I(N__38751));
    LocalMux I__7512 (
            .O(N__38751),
            .I(N__38748));
    Span4Mux_h I__7511 (
            .O(N__38748),
            .I(N__38745));
    Span4Mux_h I__7510 (
            .O(N__38745),
            .I(N__38742));
    Odrv4 I__7509 (
            .O(N__38742),
            .I(n23));
    InMux I__7508 (
            .O(N__38739),
            .I(n12977));
    InMux I__7507 (
            .O(N__38736),
            .I(N__38733));
    LocalMux I__7506 (
            .O(N__38733),
            .I(N__38730));
    Odrv4 I__7505 (
            .O(N__38730),
            .I(n22_adj_643));
    InMux I__7504 (
            .O(N__38727),
            .I(N__38724));
    LocalMux I__7503 (
            .O(N__38724),
            .I(N__38721));
    Odrv4 I__7502 (
            .O(N__38721),
            .I(n22));
    InMux I__7501 (
            .O(N__38718),
            .I(n12978));
    CascadeMux I__7500 (
            .O(N__38715),
            .I(N__38712));
    InMux I__7499 (
            .O(N__38712),
            .I(N__38709));
    LocalMux I__7498 (
            .O(N__38709),
            .I(N__38706));
    Span4Mux_v I__7497 (
            .O(N__38706),
            .I(N__38703));
    Span4Mux_h I__7496 (
            .O(N__38703),
            .I(N__38700));
    Odrv4 I__7495 (
            .O(N__38700),
            .I(n21_adj_642));
    InMux I__7494 (
            .O(N__38697),
            .I(N__38694));
    LocalMux I__7493 (
            .O(N__38694),
            .I(N__38691));
    Span4Mux_h I__7492 (
            .O(N__38691),
            .I(N__38688));
    Span4Mux_h I__7491 (
            .O(N__38688),
            .I(N__38685));
    Odrv4 I__7490 (
            .O(N__38685),
            .I(n21));
    InMux I__7489 (
            .O(N__38682),
            .I(n12979));
    CascadeMux I__7488 (
            .O(N__38679),
            .I(N__38676));
    InMux I__7487 (
            .O(N__38676),
            .I(N__38673));
    LocalMux I__7486 (
            .O(N__38673),
            .I(N__38670));
    Span4Mux_h I__7485 (
            .O(N__38670),
            .I(N__38667));
    Span4Mux_h I__7484 (
            .O(N__38667),
            .I(N__38664));
    Odrv4 I__7483 (
            .O(N__38664),
            .I(n20_adj_641));
    InMux I__7482 (
            .O(N__38661),
            .I(N__38658));
    LocalMux I__7481 (
            .O(N__38658),
            .I(N__38655));
    Span4Mux_v I__7480 (
            .O(N__38655),
            .I(N__38652));
    Span4Mux_h I__7479 (
            .O(N__38652),
            .I(N__38649));
    Odrv4 I__7478 (
            .O(N__38649),
            .I(n20));
    InMux I__7477 (
            .O(N__38646),
            .I(n12980));
    CascadeMux I__7476 (
            .O(N__38643),
            .I(N__38640));
    InMux I__7475 (
            .O(N__38640),
            .I(N__38637));
    LocalMux I__7474 (
            .O(N__38637),
            .I(N__38634));
    Span4Mux_h I__7473 (
            .O(N__38634),
            .I(N__38631));
    Odrv4 I__7472 (
            .O(N__38631),
            .I(n19_adj_640));
    InMux I__7471 (
            .O(N__38628),
            .I(N__38625));
    LocalMux I__7470 (
            .O(N__38625),
            .I(N__38622));
    Span4Mux_v I__7469 (
            .O(N__38622),
            .I(N__38619));
    Odrv4 I__7468 (
            .O(N__38619),
            .I(n19));
    InMux I__7467 (
            .O(N__38616),
            .I(n12981));
    InMux I__7466 (
            .O(N__38613),
            .I(n12982));
    CascadeMux I__7465 (
            .O(N__38610),
            .I(N__38607));
    InMux I__7464 (
            .O(N__38607),
            .I(N__38604));
    LocalMux I__7463 (
            .O(N__38604),
            .I(N__38601));
    Odrv12 I__7462 (
            .O(N__38601),
            .I(n17_adj_638));
    InMux I__7461 (
            .O(N__38598),
            .I(bfn_10_23_0_));
    InMux I__7460 (
            .O(N__38595),
            .I(n12984));
    CascadeMux I__7459 (
            .O(N__38592),
            .I(N__38589));
    InMux I__7458 (
            .O(N__38589),
            .I(N__38586));
    LocalMux I__7457 (
            .O(N__38586),
            .I(n31_adj_652));
    InMux I__7456 (
            .O(N__38583),
            .I(n12969));
    InMux I__7455 (
            .O(N__38580),
            .I(n12970));
    CascadeMux I__7454 (
            .O(N__38577),
            .I(N__38574));
    InMux I__7453 (
            .O(N__38574),
            .I(N__38571));
    LocalMux I__7452 (
            .O(N__38571),
            .I(n29_adj_650));
    InMux I__7451 (
            .O(N__38568),
            .I(N__38565));
    LocalMux I__7450 (
            .O(N__38565),
            .I(N__38562));
    Span4Mux_v I__7449 (
            .O(N__38562),
            .I(N__38559));
    Odrv4 I__7448 (
            .O(N__38559),
            .I(n29));
    InMux I__7447 (
            .O(N__38556),
            .I(n12971));
    CascadeMux I__7446 (
            .O(N__38553),
            .I(N__38550));
    InMux I__7445 (
            .O(N__38550),
            .I(N__38547));
    LocalMux I__7444 (
            .O(N__38547),
            .I(n28_adj_649));
    InMux I__7443 (
            .O(N__38544),
            .I(n12972));
    CascadeMux I__7442 (
            .O(N__38541),
            .I(N__38538));
    InMux I__7441 (
            .O(N__38538),
            .I(N__38535));
    LocalMux I__7440 (
            .O(N__38535),
            .I(n27_adj_648));
    InMux I__7439 (
            .O(N__38532),
            .I(n12973));
    CascadeMux I__7438 (
            .O(N__38529),
            .I(N__38526));
    InMux I__7437 (
            .O(N__38526),
            .I(N__38523));
    LocalMux I__7436 (
            .O(N__38523),
            .I(n26_adj_647));
    InMux I__7435 (
            .O(N__38520),
            .I(n12974));
    CascadeMux I__7434 (
            .O(N__38517),
            .I(N__38514));
    InMux I__7433 (
            .O(N__38514),
            .I(N__38511));
    LocalMux I__7432 (
            .O(N__38511),
            .I(N__38508));
    Span4Mux_v I__7431 (
            .O(N__38508),
            .I(N__38505));
    Span4Mux_h I__7430 (
            .O(N__38505),
            .I(N__38502));
    Odrv4 I__7429 (
            .O(N__38502),
            .I(n25_adj_646));
    InMux I__7428 (
            .O(N__38499),
            .I(N__38496));
    LocalMux I__7427 (
            .O(N__38496),
            .I(N__38493));
    Span4Mux_h I__7426 (
            .O(N__38493),
            .I(N__38490));
    Span4Mux_h I__7425 (
            .O(N__38490),
            .I(N__38487));
    Odrv4 I__7424 (
            .O(N__38487),
            .I(n25_adj_551));
    InMux I__7423 (
            .O(N__38484),
            .I(bfn_10_22_0_));
    CascadeMux I__7422 (
            .O(N__38481),
            .I(N__38478));
    InMux I__7421 (
            .O(N__38478),
            .I(N__38475));
    LocalMux I__7420 (
            .O(N__38475),
            .I(N__38472));
    Odrv4 I__7419 (
            .O(N__38472),
            .I(n24_adj_645));
    InMux I__7418 (
            .O(N__38469),
            .I(N__38466));
    LocalMux I__7417 (
            .O(N__38466),
            .I(N__38463));
    Odrv12 I__7416 (
            .O(N__38463),
            .I(n24));
    InMux I__7415 (
            .O(N__38460),
            .I(n12976));
    CascadeMux I__7414 (
            .O(N__38457),
            .I(N__38453));
    InMux I__7413 (
            .O(N__38456),
            .I(N__38450));
    InMux I__7412 (
            .O(N__38453),
            .I(N__38447));
    LocalMux I__7411 (
            .O(N__38450),
            .I(N__38444));
    LocalMux I__7410 (
            .O(N__38447),
            .I(n1932));
    Odrv4 I__7409 (
            .O(N__38444),
            .I(n1932));
    CascadeMux I__7408 (
            .O(N__38439),
            .I(n1932_cascade_));
    InMux I__7407 (
            .O(N__38436),
            .I(N__38433));
    LocalMux I__7406 (
            .O(N__38433),
            .I(N__38430));
    Odrv4 I__7405 (
            .O(N__38430),
            .I(n1999));
    CascadeMux I__7404 (
            .O(N__38427),
            .I(N__38424));
    InMux I__7403 (
            .O(N__38424),
            .I(N__38420));
    InMux I__7402 (
            .O(N__38423),
            .I(N__38417));
    LocalMux I__7401 (
            .O(N__38420),
            .I(N__38414));
    LocalMux I__7400 (
            .O(N__38417),
            .I(N__38411));
    Span4Mux_h I__7399 (
            .O(N__38414),
            .I(N__38408));
    Odrv4 I__7398 (
            .O(N__38411),
            .I(n2031));
    Odrv4 I__7397 (
            .O(N__38408),
            .I(n2031));
    InMux I__7396 (
            .O(N__38403),
            .I(N__38399));
    InMux I__7395 (
            .O(N__38402),
            .I(N__38395));
    LocalMux I__7394 (
            .O(N__38399),
            .I(N__38392));
    InMux I__7393 (
            .O(N__38398),
            .I(N__38389));
    LocalMux I__7392 (
            .O(N__38395),
            .I(N__38386));
    Span4Mux_v I__7391 (
            .O(N__38392),
            .I(N__38383));
    LocalMux I__7390 (
            .O(N__38389),
            .I(N__38378));
    Span4Mux_v I__7389 (
            .O(N__38386),
            .I(N__38378));
    Span4Mux_h I__7388 (
            .O(N__38383),
            .I(N__38375));
    Odrv4 I__7387 (
            .O(N__38378),
            .I(n306));
    Odrv4 I__7386 (
            .O(N__38375),
            .I(n306));
    CascadeMux I__7385 (
            .O(N__38370),
            .I(n2031_cascade_));
    InMux I__7384 (
            .O(N__38367),
            .I(N__38364));
    LocalMux I__7383 (
            .O(N__38364),
            .I(n11964));
    InMux I__7382 (
            .O(N__38361),
            .I(N__38354));
    InMux I__7381 (
            .O(N__38360),
            .I(N__38354));
    InMux I__7380 (
            .O(N__38359),
            .I(N__38351));
    LocalMux I__7379 (
            .O(N__38354),
            .I(N__38348));
    LocalMux I__7378 (
            .O(N__38351),
            .I(N__38345));
    Span4Mux_v I__7377 (
            .O(N__38348),
            .I(N__38342));
    Sp12to4 I__7376 (
            .O(N__38345),
            .I(N__38339));
    Odrv4 I__7375 (
            .O(N__38342),
            .I(n305));
    Odrv12 I__7374 (
            .O(N__38339),
            .I(n305));
    InMux I__7373 (
            .O(N__38334),
            .I(N__38331));
    LocalMux I__7372 (
            .O(N__38331),
            .I(N__38328));
    Span4Mux_v I__7371 (
            .O(N__38328),
            .I(N__38325));
    Odrv4 I__7370 (
            .O(N__38325),
            .I(n2001));
    CascadeMux I__7369 (
            .O(N__38322),
            .I(N__38318));
    CascadeMux I__7368 (
            .O(N__38321),
            .I(N__38315));
    InMux I__7367 (
            .O(N__38318),
            .I(N__38312));
    InMux I__7366 (
            .O(N__38315),
            .I(N__38309));
    LocalMux I__7365 (
            .O(N__38312),
            .I(N__38306));
    LocalMux I__7364 (
            .O(N__38309),
            .I(N__38303));
    Span4Mux_v I__7363 (
            .O(N__38306),
            .I(N__38297));
    Span4Mux_v I__7362 (
            .O(N__38303),
            .I(N__38297));
    InMux I__7361 (
            .O(N__38302),
            .I(N__38294));
    Odrv4 I__7360 (
            .O(N__38297),
            .I(n2033));
    LocalMux I__7359 (
            .O(N__38294),
            .I(n2033));
    InMux I__7358 (
            .O(N__38289),
            .I(N__38286));
    LocalMux I__7357 (
            .O(N__38286),
            .I(N__38283));
    Odrv4 I__7356 (
            .O(N__38283),
            .I(n1996));
    CascadeMux I__7355 (
            .O(N__38280),
            .I(N__38276));
    InMux I__7354 (
            .O(N__38279),
            .I(N__38273));
    InMux I__7353 (
            .O(N__38276),
            .I(N__38270));
    LocalMux I__7352 (
            .O(N__38273),
            .I(N__38264));
    LocalMux I__7351 (
            .O(N__38270),
            .I(N__38264));
    CascadeMux I__7350 (
            .O(N__38269),
            .I(N__38261));
    Span4Mux_v I__7349 (
            .O(N__38264),
            .I(N__38258));
    InMux I__7348 (
            .O(N__38261),
            .I(N__38255));
    Odrv4 I__7347 (
            .O(N__38258),
            .I(n2028));
    LocalMux I__7346 (
            .O(N__38255),
            .I(n2028));
    InMux I__7345 (
            .O(N__38250),
            .I(N__38247));
    LocalMux I__7344 (
            .O(N__38247),
            .I(N__38244));
    Span4Mux_v I__7343 (
            .O(N__38244),
            .I(N__38241));
    Odrv4 I__7342 (
            .O(N__38241),
            .I(n2000));
    CascadeMux I__7341 (
            .O(N__38238),
            .I(N__38235));
    InMux I__7340 (
            .O(N__38235),
            .I(N__38228));
    InMux I__7339 (
            .O(N__38234),
            .I(N__38228));
    InMux I__7338 (
            .O(N__38233),
            .I(N__38225));
    LocalMux I__7337 (
            .O(N__38228),
            .I(N__38222));
    LocalMux I__7336 (
            .O(N__38225),
            .I(n1933));
    Odrv4 I__7335 (
            .O(N__38222),
            .I(n1933));
    InMux I__7334 (
            .O(N__38217),
            .I(N__38214));
    LocalMux I__7333 (
            .O(N__38214),
            .I(N__38211));
    Span4Mux_v I__7332 (
            .O(N__38211),
            .I(N__38202));
    InMux I__7331 (
            .O(N__38210),
            .I(N__38199));
    CascadeMux I__7330 (
            .O(N__38209),
            .I(N__38192));
    CascadeMux I__7329 (
            .O(N__38208),
            .I(N__38188));
    CascadeMux I__7328 (
            .O(N__38207),
            .I(N__38185));
    CascadeMux I__7327 (
            .O(N__38206),
            .I(N__38181));
    CascadeMux I__7326 (
            .O(N__38205),
            .I(N__38175));
    Span4Mux_v I__7325 (
            .O(N__38202),
            .I(N__38168));
    LocalMux I__7324 (
            .O(N__38199),
            .I(N__38168));
    InMux I__7323 (
            .O(N__38198),
            .I(N__38161));
    InMux I__7322 (
            .O(N__38197),
            .I(N__38161));
    InMux I__7321 (
            .O(N__38196),
            .I(N__38161));
    InMux I__7320 (
            .O(N__38195),
            .I(N__38148));
    InMux I__7319 (
            .O(N__38192),
            .I(N__38148));
    InMux I__7318 (
            .O(N__38191),
            .I(N__38148));
    InMux I__7317 (
            .O(N__38188),
            .I(N__38148));
    InMux I__7316 (
            .O(N__38185),
            .I(N__38148));
    InMux I__7315 (
            .O(N__38184),
            .I(N__38148));
    InMux I__7314 (
            .O(N__38181),
            .I(N__38143));
    InMux I__7313 (
            .O(N__38180),
            .I(N__38143));
    InMux I__7312 (
            .O(N__38179),
            .I(N__38134));
    InMux I__7311 (
            .O(N__38178),
            .I(N__38134));
    InMux I__7310 (
            .O(N__38175),
            .I(N__38134));
    InMux I__7309 (
            .O(N__38174),
            .I(N__38134));
    InMux I__7308 (
            .O(N__38173),
            .I(N__38131));
    Odrv4 I__7307 (
            .O(N__38168),
            .I(n1950));
    LocalMux I__7306 (
            .O(N__38161),
            .I(n1950));
    LocalMux I__7305 (
            .O(N__38148),
            .I(n1950));
    LocalMux I__7304 (
            .O(N__38143),
            .I(n1950));
    LocalMux I__7303 (
            .O(N__38134),
            .I(n1950));
    LocalMux I__7302 (
            .O(N__38131),
            .I(n1950));
    CascadeMux I__7301 (
            .O(N__38118),
            .I(N__38114));
    CascadeMux I__7300 (
            .O(N__38117),
            .I(N__38111));
    InMux I__7299 (
            .O(N__38114),
            .I(N__38108));
    InMux I__7298 (
            .O(N__38111),
            .I(N__38105));
    LocalMux I__7297 (
            .O(N__38108),
            .I(N__38100));
    LocalMux I__7296 (
            .O(N__38105),
            .I(N__38100));
    Span4Mux_h I__7295 (
            .O(N__38100),
            .I(N__38096));
    InMux I__7294 (
            .O(N__38099),
            .I(N__38093));
    Odrv4 I__7293 (
            .O(N__38096),
            .I(n2032));
    LocalMux I__7292 (
            .O(N__38093),
            .I(n2032));
    CascadeMux I__7291 (
            .O(N__38088),
            .I(N__38085));
    InMux I__7290 (
            .O(N__38085),
            .I(N__38082));
    LocalMux I__7289 (
            .O(N__38082),
            .I(n33_adj_654));
    InMux I__7288 (
            .O(N__38079),
            .I(N__38076));
    LocalMux I__7287 (
            .O(N__38076),
            .I(N__38073));
    Span4Mux_h I__7286 (
            .O(N__38073),
            .I(N__38070));
    Odrv4 I__7285 (
            .O(N__38070),
            .I(n33));
    InMux I__7284 (
            .O(N__38067),
            .I(bfn_10_21_0_));
    CascadeMux I__7283 (
            .O(N__38064),
            .I(N__38061));
    InMux I__7282 (
            .O(N__38061),
            .I(N__38058));
    LocalMux I__7281 (
            .O(N__38058),
            .I(n32_adj_653));
    InMux I__7280 (
            .O(N__38055),
            .I(n12968));
    CascadeMux I__7279 (
            .O(N__38052),
            .I(N__38049));
    InMux I__7278 (
            .O(N__38049),
            .I(N__38045));
    InMux I__7277 (
            .O(N__38048),
            .I(N__38042));
    LocalMux I__7276 (
            .O(N__38045),
            .I(n1922));
    LocalMux I__7275 (
            .O(N__38042),
            .I(n1922));
    InMux I__7274 (
            .O(N__38037),
            .I(N__38034));
    LocalMux I__7273 (
            .O(N__38034),
            .I(n1989));
    CascadeMux I__7272 (
            .O(N__38031),
            .I(n1922_cascade_));
    CascadeMux I__7271 (
            .O(N__38028),
            .I(N__38025));
    InMux I__7270 (
            .O(N__38025),
            .I(N__38021));
    InMux I__7269 (
            .O(N__38024),
            .I(N__38018));
    LocalMux I__7268 (
            .O(N__38021),
            .I(N__38015));
    LocalMux I__7267 (
            .O(N__38018),
            .I(N__38012));
    Span4Mux_h I__7266 (
            .O(N__38015),
            .I(N__38006));
    Span4Mux_v I__7265 (
            .O(N__38012),
            .I(N__38006));
    InMux I__7264 (
            .O(N__38011),
            .I(N__38003));
    Odrv4 I__7263 (
            .O(N__38006),
            .I(n2021));
    LocalMux I__7262 (
            .O(N__38003),
            .I(n2021));
    InMux I__7261 (
            .O(N__37998),
            .I(N__37995));
    LocalMux I__7260 (
            .O(N__37995),
            .I(n14416));
    CascadeMux I__7259 (
            .O(N__37992),
            .I(n14420_cascade_));
    CascadeMux I__7258 (
            .O(N__37989),
            .I(n1950_cascade_));
    InMux I__7257 (
            .O(N__37986),
            .I(N__37983));
    LocalMux I__7256 (
            .O(N__37983),
            .I(N__37980));
    Span4Mux_v I__7255 (
            .O(N__37980),
            .I(N__37977));
    Odrv4 I__7254 (
            .O(N__37977),
            .I(n1998));
    CascadeMux I__7253 (
            .O(N__37974),
            .I(N__37970));
    CascadeMux I__7252 (
            .O(N__37973),
            .I(N__37967));
    InMux I__7251 (
            .O(N__37970),
            .I(N__37963));
    InMux I__7250 (
            .O(N__37967),
            .I(N__37960));
    InMux I__7249 (
            .O(N__37966),
            .I(N__37957));
    LocalMux I__7248 (
            .O(N__37963),
            .I(N__37952));
    LocalMux I__7247 (
            .O(N__37960),
            .I(N__37952));
    LocalMux I__7246 (
            .O(N__37957),
            .I(N__37947));
    Span4Mux_h I__7245 (
            .O(N__37952),
            .I(N__37947));
    Odrv4 I__7244 (
            .O(N__37947),
            .I(n2030));
    InMux I__7243 (
            .O(N__37944),
            .I(N__37941));
    LocalMux I__7242 (
            .O(N__37941),
            .I(N__37938));
    Span12Mux_s9_h I__7241 (
            .O(N__37938),
            .I(N__37934));
    InMux I__7240 (
            .O(N__37937),
            .I(N__37931));
    Odrv12 I__7239 (
            .O(N__37934),
            .I(n15666));
    LocalMux I__7238 (
            .O(N__37931),
            .I(n15666));
    CascadeMux I__7237 (
            .O(N__37926),
            .I(N__37923));
    InMux I__7236 (
            .O(N__37923),
            .I(N__37919));
    InMux I__7235 (
            .O(N__37922),
            .I(N__37916));
    LocalMux I__7234 (
            .O(N__37919),
            .I(n1917));
    LocalMux I__7233 (
            .O(N__37916),
            .I(n1917));
    InMux I__7232 (
            .O(N__37911),
            .I(N__37908));
    LocalMux I__7231 (
            .O(N__37908),
            .I(n1988));
    CascadeMux I__7230 (
            .O(N__37905),
            .I(N__37901));
    CascadeMux I__7229 (
            .O(N__37904),
            .I(N__37898));
    InMux I__7228 (
            .O(N__37901),
            .I(N__37895));
    InMux I__7227 (
            .O(N__37898),
            .I(N__37892));
    LocalMux I__7226 (
            .O(N__37895),
            .I(n1921));
    LocalMux I__7225 (
            .O(N__37892),
            .I(n1921));
    CascadeMux I__7224 (
            .O(N__37887),
            .I(N__37883));
    InMux I__7223 (
            .O(N__37886),
            .I(N__37880));
    InMux I__7222 (
            .O(N__37883),
            .I(N__37877));
    LocalMux I__7221 (
            .O(N__37880),
            .I(N__37874));
    LocalMux I__7220 (
            .O(N__37877),
            .I(N__37871));
    Span4Mux_h I__7219 (
            .O(N__37874),
            .I(N__37867));
    Span4Mux_h I__7218 (
            .O(N__37871),
            .I(N__37864));
    InMux I__7217 (
            .O(N__37870),
            .I(N__37861));
    Odrv4 I__7216 (
            .O(N__37867),
            .I(n2020));
    Odrv4 I__7215 (
            .O(N__37864),
            .I(n2020));
    LocalMux I__7214 (
            .O(N__37861),
            .I(n2020));
    InMux I__7213 (
            .O(N__37854),
            .I(N__37851));
    LocalMux I__7212 (
            .O(N__37851),
            .I(n11966));
    InMux I__7211 (
            .O(N__37848),
            .I(N__37844));
    InMux I__7210 (
            .O(N__37847),
            .I(N__37841));
    LocalMux I__7209 (
            .O(N__37844),
            .I(N__37837));
    LocalMux I__7208 (
            .O(N__37841),
            .I(N__37834));
    InMux I__7207 (
            .O(N__37840),
            .I(N__37831));
    Span4Mux_v I__7206 (
            .O(N__37837),
            .I(N__37828));
    Span4Mux_v I__7205 (
            .O(N__37834),
            .I(N__37825));
    LocalMux I__7204 (
            .O(N__37831),
            .I(encoder0_position_9));
    Odrv4 I__7203 (
            .O(N__37828),
            .I(encoder0_position_9));
    Odrv4 I__7202 (
            .O(N__37825),
            .I(encoder0_position_9));
    InMux I__7201 (
            .O(N__37818),
            .I(N__37813));
    InMux I__7200 (
            .O(N__37817),
            .I(N__37810));
    InMux I__7199 (
            .O(N__37816),
            .I(N__37807));
    LocalMux I__7198 (
            .O(N__37813),
            .I(N__37800));
    LocalMux I__7197 (
            .O(N__37810),
            .I(N__37800));
    LocalMux I__7196 (
            .O(N__37807),
            .I(N__37800));
    Odrv12 I__7195 (
            .O(N__37800),
            .I(n310));
    CascadeMux I__7194 (
            .O(N__37797),
            .I(N__37794));
    InMux I__7193 (
            .O(N__37794),
            .I(N__37791));
    LocalMux I__7192 (
            .O(N__37791),
            .I(N__37788));
    Span4Mux_h I__7191 (
            .O(N__37788),
            .I(N__37783));
    InMux I__7190 (
            .O(N__37787),
            .I(N__37780));
    InMux I__7189 (
            .O(N__37786),
            .I(N__37777));
    Odrv4 I__7188 (
            .O(N__37783),
            .I(n1927));
    LocalMux I__7187 (
            .O(N__37780),
            .I(n1927));
    LocalMux I__7186 (
            .O(N__37777),
            .I(n1927));
    InMux I__7185 (
            .O(N__37770),
            .I(N__37766));
    CascadeMux I__7184 (
            .O(N__37769),
            .I(N__37763));
    LocalMux I__7183 (
            .O(N__37766),
            .I(N__37760));
    InMux I__7182 (
            .O(N__37763),
            .I(N__37757));
    Odrv4 I__7181 (
            .O(N__37760),
            .I(n1923));
    LocalMux I__7180 (
            .O(N__37757),
            .I(n1923));
    CascadeMux I__7179 (
            .O(N__37752),
            .I(N__37749));
    InMux I__7178 (
            .O(N__37749),
            .I(N__37745));
    CascadeMux I__7177 (
            .O(N__37748),
            .I(N__37742));
    LocalMux I__7176 (
            .O(N__37745),
            .I(N__37738));
    InMux I__7175 (
            .O(N__37742),
            .I(N__37735));
    InMux I__7174 (
            .O(N__37741),
            .I(N__37732));
    Odrv4 I__7173 (
            .O(N__37738),
            .I(n1926));
    LocalMux I__7172 (
            .O(N__37735),
            .I(n1926));
    LocalMux I__7171 (
            .O(N__37732),
            .I(n1926));
    CascadeMux I__7170 (
            .O(N__37725),
            .I(n1923_cascade_));
    InMux I__7169 (
            .O(N__37722),
            .I(N__37718));
    CascadeMux I__7168 (
            .O(N__37721),
            .I(N__37715));
    LocalMux I__7167 (
            .O(N__37718),
            .I(N__37711));
    InMux I__7166 (
            .O(N__37715),
            .I(N__37708));
    InMux I__7165 (
            .O(N__37714),
            .I(N__37705));
    Odrv4 I__7164 (
            .O(N__37711),
            .I(n1924));
    LocalMux I__7163 (
            .O(N__37708),
            .I(n1924));
    LocalMux I__7162 (
            .O(N__37705),
            .I(n1924));
    InMux I__7161 (
            .O(N__37698),
            .I(N__37695));
    LocalMux I__7160 (
            .O(N__37695),
            .I(n14408));
    CascadeMux I__7159 (
            .O(N__37692),
            .I(n1921_cascade_));
    InMux I__7158 (
            .O(N__37689),
            .I(N__37686));
    LocalMux I__7157 (
            .O(N__37686),
            .I(n14410));
    InMux I__7156 (
            .O(N__37683),
            .I(N__37680));
    LocalMux I__7155 (
            .O(N__37680),
            .I(n1995));
    CascadeMux I__7154 (
            .O(N__37677),
            .I(N__37673));
    CascadeMux I__7153 (
            .O(N__37676),
            .I(N__37670));
    InMux I__7152 (
            .O(N__37673),
            .I(N__37667));
    InMux I__7151 (
            .O(N__37670),
            .I(N__37664));
    LocalMux I__7150 (
            .O(N__37667),
            .I(N__37660));
    LocalMux I__7149 (
            .O(N__37664),
            .I(N__37657));
    InMux I__7148 (
            .O(N__37663),
            .I(N__37654));
    Span4Mux_h I__7147 (
            .O(N__37660),
            .I(N__37651));
    Span4Mux_h I__7146 (
            .O(N__37657),
            .I(N__37646));
    LocalMux I__7145 (
            .O(N__37654),
            .I(N__37646));
    Odrv4 I__7144 (
            .O(N__37651),
            .I(n2027));
    Odrv4 I__7143 (
            .O(N__37646),
            .I(n2027));
    CascadeMux I__7142 (
            .O(N__37641),
            .I(N__37636));
    CascadeMux I__7141 (
            .O(N__37640),
            .I(N__37633));
    InMux I__7140 (
            .O(N__37639),
            .I(N__37630));
    InMux I__7139 (
            .O(N__37636),
            .I(N__37627));
    InMux I__7138 (
            .O(N__37633),
            .I(N__37624));
    LocalMux I__7137 (
            .O(N__37630),
            .I(n1925));
    LocalMux I__7136 (
            .O(N__37627),
            .I(n1925));
    LocalMux I__7135 (
            .O(N__37624),
            .I(n1925));
    InMux I__7134 (
            .O(N__37617),
            .I(N__37614));
    LocalMux I__7133 (
            .O(N__37614),
            .I(N__37611));
    Odrv12 I__7132 (
            .O(N__37611),
            .I(n6_adj_586));
    InMux I__7131 (
            .O(N__37608),
            .I(n12430));
    InMux I__7130 (
            .O(N__37605),
            .I(n12431));
    InMux I__7129 (
            .O(N__37602),
            .I(n12432));
    InMux I__7128 (
            .O(N__37599),
            .I(n12433));
    InMux I__7127 (
            .O(N__37596),
            .I(n12434));
    InMux I__7126 (
            .O(N__37593),
            .I(n12421));
    InMux I__7125 (
            .O(N__37590),
            .I(N__37587));
    LocalMux I__7124 (
            .O(N__37587),
            .I(N__37584));
    Odrv4 I__7123 (
            .O(N__37584),
            .I(n14_adj_594));
    InMux I__7122 (
            .O(N__37581),
            .I(n12422));
    InMux I__7121 (
            .O(N__37578),
            .I(N__37575));
    LocalMux I__7120 (
            .O(N__37575),
            .I(N__37572));
    Odrv4 I__7119 (
            .O(N__37572),
            .I(n13_adj_593));
    InMux I__7118 (
            .O(N__37569),
            .I(n12423));
    InMux I__7117 (
            .O(N__37566),
            .I(n12424));
    InMux I__7116 (
            .O(N__37563),
            .I(n12425));
    InMux I__7115 (
            .O(N__37560),
            .I(N__37557));
    LocalMux I__7114 (
            .O(N__37557),
            .I(N__37554));
    Odrv4 I__7113 (
            .O(N__37554),
            .I(n10_adj_590));
    InMux I__7112 (
            .O(N__37551),
            .I(n12426));
    InMux I__7111 (
            .O(N__37548),
            .I(bfn_9_32_0_));
    InMux I__7110 (
            .O(N__37545),
            .I(n12428));
    InMux I__7109 (
            .O(N__37542),
            .I(n12429));
    InMux I__7108 (
            .O(N__37539),
            .I(N__37536));
    LocalMux I__7107 (
            .O(N__37536),
            .I(N__37533));
    Odrv4 I__7106 (
            .O(N__37533),
            .I(n24_adj_604));
    InMux I__7105 (
            .O(N__37530),
            .I(N__37527));
    LocalMux I__7104 (
            .O(N__37527),
            .I(N__37524));
    Odrv12 I__7103 (
            .O(N__37524),
            .I(pwm_setpoint_23_N_171_1));
    InMux I__7102 (
            .O(N__37521),
            .I(n12412));
    InMux I__7101 (
            .O(N__37518),
            .I(N__37515));
    LocalMux I__7100 (
            .O(N__37515),
            .I(N__37512));
    Odrv4 I__7099 (
            .O(N__37512),
            .I(n23_adj_603));
    InMux I__7098 (
            .O(N__37509),
            .I(n12413));
    InMux I__7097 (
            .O(N__37506),
            .I(N__37503));
    LocalMux I__7096 (
            .O(N__37503),
            .I(n22_adj_602));
    InMux I__7095 (
            .O(N__37500),
            .I(n12414));
    InMux I__7094 (
            .O(N__37497),
            .I(n12415));
    InMux I__7093 (
            .O(N__37494),
            .I(n12416));
    InMux I__7092 (
            .O(N__37491),
            .I(n12417));
    InMux I__7091 (
            .O(N__37488),
            .I(N__37485));
    LocalMux I__7090 (
            .O(N__37485),
            .I(N__37482));
    Odrv4 I__7089 (
            .O(N__37482),
            .I(n18_adj_598));
    InMux I__7088 (
            .O(N__37479),
            .I(n12418));
    InMux I__7087 (
            .O(N__37476),
            .I(N__37473));
    LocalMux I__7086 (
            .O(N__37473),
            .I(N__37470));
    Odrv4 I__7085 (
            .O(N__37470),
            .I(n17_adj_597));
    InMux I__7084 (
            .O(N__37467),
            .I(bfn_9_31_0_));
    InMux I__7083 (
            .O(N__37464),
            .I(n12420));
    InMux I__7082 (
            .O(N__37461),
            .I(N__37458));
    LocalMux I__7081 (
            .O(N__37458),
            .I(N__37455));
    Span4Mux_v I__7080 (
            .O(N__37455),
            .I(N__37452));
    Odrv4 I__7079 (
            .O(N__37452),
            .I(encoder0_position_scaled_19));
    InMux I__7078 (
            .O(N__37449),
            .I(N__37446));
    LocalMux I__7077 (
            .O(N__37446),
            .I(N__37443));
    Odrv4 I__7076 (
            .O(N__37443),
            .I(n25_adj_605));
    InMux I__7075 (
            .O(N__37440),
            .I(N__37437));
    LocalMux I__7074 (
            .O(N__37437),
            .I(N__37434));
    Odrv12 I__7073 (
            .O(N__37434),
            .I(pwm_setpoint_23_N_171_0));
    InMux I__7072 (
            .O(N__37431),
            .I(bfn_9_30_0_));
    CascadeMux I__7071 (
            .O(N__37428),
            .I(\quad_counter0.a_prev_N_543_cascade_ ));
    CascadeMux I__7070 (
            .O(N__37425),
            .I(N__37408));
    CascadeMux I__7069 (
            .O(N__37424),
            .I(N__37404));
    CascadeMux I__7068 (
            .O(N__37423),
            .I(N__37400));
    CascadeMux I__7067 (
            .O(N__37422),
            .I(N__37396));
    CascadeMux I__7066 (
            .O(N__37421),
            .I(N__37393));
    CascadeMux I__7065 (
            .O(N__37420),
            .I(N__37389));
    CascadeMux I__7064 (
            .O(N__37419),
            .I(N__37385));
    CascadeMux I__7063 (
            .O(N__37418),
            .I(N__37381));
    CascadeMux I__7062 (
            .O(N__37417),
            .I(N__37376));
    CascadeMux I__7061 (
            .O(N__37416),
            .I(N__37372));
    CascadeMux I__7060 (
            .O(N__37415),
            .I(N__37368));
    CascadeMux I__7059 (
            .O(N__37414),
            .I(N__37362));
    CascadeMux I__7058 (
            .O(N__37413),
            .I(N__37358));
    CascadeMux I__7057 (
            .O(N__37412),
            .I(N__37354));
    InMux I__7056 (
            .O(N__37411),
            .I(N__37336));
    InMux I__7055 (
            .O(N__37408),
            .I(N__37336));
    InMux I__7054 (
            .O(N__37407),
            .I(N__37336));
    InMux I__7053 (
            .O(N__37404),
            .I(N__37336));
    InMux I__7052 (
            .O(N__37403),
            .I(N__37336));
    InMux I__7051 (
            .O(N__37400),
            .I(N__37336));
    InMux I__7050 (
            .O(N__37399),
            .I(N__37336));
    InMux I__7049 (
            .O(N__37396),
            .I(N__37336));
    InMux I__7048 (
            .O(N__37393),
            .I(N__37319));
    InMux I__7047 (
            .O(N__37392),
            .I(N__37319));
    InMux I__7046 (
            .O(N__37389),
            .I(N__37319));
    InMux I__7045 (
            .O(N__37388),
            .I(N__37319));
    InMux I__7044 (
            .O(N__37385),
            .I(N__37319));
    InMux I__7043 (
            .O(N__37384),
            .I(N__37319));
    InMux I__7042 (
            .O(N__37381),
            .I(N__37319));
    InMux I__7041 (
            .O(N__37380),
            .I(N__37319));
    InMux I__7040 (
            .O(N__37379),
            .I(N__37304));
    InMux I__7039 (
            .O(N__37376),
            .I(N__37304));
    InMux I__7038 (
            .O(N__37375),
            .I(N__37304));
    InMux I__7037 (
            .O(N__37372),
            .I(N__37304));
    InMux I__7036 (
            .O(N__37371),
            .I(N__37304));
    InMux I__7035 (
            .O(N__37368),
            .I(N__37304));
    InMux I__7034 (
            .O(N__37367),
            .I(N__37304));
    InMux I__7033 (
            .O(N__37366),
            .I(N__37287));
    InMux I__7032 (
            .O(N__37365),
            .I(N__37287));
    InMux I__7031 (
            .O(N__37362),
            .I(N__37287));
    InMux I__7030 (
            .O(N__37361),
            .I(N__37287));
    InMux I__7029 (
            .O(N__37358),
            .I(N__37287));
    InMux I__7028 (
            .O(N__37357),
            .I(N__37287));
    InMux I__7027 (
            .O(N__37354),
            .I(N__37287));
    InMux I__7026 (
            .O(N__37353),
            .I(N__37287));
    LocalMux I__7025 (
            .O(N__37336),
            .I(N__37280));
    LocalMux I__7024 (
            .O(N__37319),
            .I(N__37280));
    LocalMux I__7023 (
            .O(N__37304),
            .I(N__37280));
    LocalMux I__7022 (
            .O(N__37287),
            .I(N__37277));
    Span4Mux_v I__7021 (
            .O(N__37280),
            .I(N__37274));
    Odrv4 I__7020 (
            .O(N__37277),
            .I(\quad_counter0.direction_N_536 ));
    Odrv4 I__7019 (
            .O(N__37274),
            .I(\quad_counter0.direction_N_536 ));
    CascadeMux I__7018 (
            .O(N__37269),
            .I(N__37266));
    InMux I__7017 (
            .O(N__37266),
            .I(N__37262));
    InMux I__7016 (
            .O(N__37265),
            .I(N__37259));
    LocalMux I__7015 (
            .O(N__37262),
            .I(N__37256));
    LocalMux I__7014 (
            .O(N__37259),
            .I(N__37252));
    Span4Mux_h I__7013 (
            .O(N__37256),
            .I(N__37249));
    InMux I__7012 (
            .O(N__37255),
            .I(N__37246));
    Odrv12 I__7011 (
            .O(N__37252),
            .I(n3024));
    Odrv4 I__7010 (
            .O(N__37249),
            .I(n3024));
    LocalMux I__7009 (
            .O(N__37246),
            .I(n3024));
    CascadeMux I__7008 (
            .O(N__37239),
            .I(N__37236));
    InMux I__7007 (
            .O(N__37236),
            .I(N__37233));
    LocalMux I__7006 (
            .O(N__37233),
            .I(N__37230));
    Span12Mux_h I__7005 (
            .O(N__37230),
            .I(N__37227));
    Odrv12 I__7004 (
            .O(N__37227),
            .I(n3091));
    CascadeMux I__7003 (
            .O(N__37224),
            .I(N__37220));
    CascadeMux I__7002 (
            .O(N__37223),
            .I(N__37212));
    InMux I__7001 (
            .O(N__37220),
            .I(N__37207));
    InMux I__7000 (
            .O(N__37219),
            .I(N__37200));
    CascadeMux I__6999 (
            .O(N__37218),
            .I(N__37197));
    CascadeMux I__6998 (
            .O(N__37217),
            .I(N__37190));
    InMux I__6997 (
            .O(N__37216),
            .I(N__37187));
    InMux I__6996 (
            .O(N__37215),
            .I(N__37184));
    InMux I__6995 (
            .O(N__37212),
            .I(N__37179));
    InMux I__6994 (
            .O(N__37211),
            .I(N__37179));
    InMux I__6993 (
            .O(N__37210),
            .I(N__37176));
    LocalMux I__6992 (
            .O(N__37207),
            .I(N__37173));
    CascadeMux I__6991 (
            .O(N__37206),
            .I(N__37166));
    CascadeMux I__6990 (
            .O(N__37205),
            .I(N__37163));
    CascadeMux I__6989 (
            .O(N__37204),
            .I(N__37159));
    CascadeMux I__6988 (
            .O(N__37203),
            .I(N__37150));
    LocalMux I__6987 (
            .O(N__37200),
            .I(N__37146));
    InMux I__6986 (
            .O(N__37197),
            .I(N__37141));
    InMux I__6985 (
            .O(N__37196),
            .I(N__37141));
    InMux I__6984 (
            .O(N__37195),
            .I(N__37132));
    InMux I__6983 (
            .O(N__37194),
            .I(N__37132));
    InMux I__6982 (
            .O(N__37193),
            .I(N__37132));
    InMux I__6981 (
            .O(N__37190),
            .I(N__37132));
    LocalMux I__6980 (
            .O(N__37187),
            .I(N__37127));
    LocalMux I__6979 (
            .O(N__37184),
            .I(N__37127));
    LocalMux I__6978 (
            .O(N__37179),
            .I(N__37124));
    LocalMux I__6977 (
            .O(N__37176),
            .I(N__37121));
    Span12Mux_v I__6976 (
            .O(N__37173),
            .I(N__37118));
    InMux I__6975 (
            .O(N__37172),
            .I(N__37113));
    InMux I__6974 (
            .O(N__37171),
            .I(N__37113));
    InMux I__6973 (
            .O(N__37170),
            .I(N__37110));
    InMux I__6972 (
            .O(N__37169),
            .I(N__37101));
    InMux I__6971 (
            .O(N__37166),
            .I(N__37101));
    InMux I__6970 (
            .O(N__37163),
            .I(N__37101));
    InMux I__6969 (
            .O(N__37162),
            .I(N__37101));
    InMux I__6968 (
            .O(N__37159),
            .I(N__37096));
    InMux I__6967 (
            .O(N__37158),
            .I(N__37096));
    InMux I__6966 (
            .O(N__37157),
            .I(N__37093));
    InMux I__6965 (
            .O(N__37156),
            .I(N__37088));
    InMux I__6964 (
            .O(N__37155),
            .I(N__37088));
    InMux I__6963 (
            .O(N__37154),
            .I(N__37079));
    InMux I__6962 (
            .O(N__37153),
            .I(N__37079));
    InMux I__6961 (
            .O(N__37150),
            .I(N__37079));
    InMux I__6960 (
            .O(N__37149),
            .I(N__37079));
    Span4Mux_h I__6959 (
            .O(N__37146),
            .I(N__37070));
    LocalMux I__6958 (
            .O(N__37141),
            .I(N__37070));
    LocalMux I__6957 (
            .O(N__37132),
            .I(N__37070));
    Span4Mux_h I__6956 (
            .O(N__37127),
            .I(N__37070));
    Span4Mux_h I__6955 (
            .O(N__37124),
            .I(N__37065));
    Span4Mux_v I__6954 (
            .O(N__37121),
            .I(N__37065));
    Odrv12 I__6953 (
            .O(N__37118),
            .I(n3039));
    LocalMux I__6952 (
            .O(N__37113),
            .I(n3039));
    LocalMux I__6951 (
            .O(N__37110),
            .I(n3039));
    LocalMux I__6950 (
            .O(N__37101),
            .I(n3039));
    LocalMux I__6949 (
            .O(N__37096),
            .I(n3039));
    LocalMux I__6948 (
            .O(N__37093),
            .I(n3039));
    LocalMux I__6947 (
            .O(N__37088),
            .I(n3039));
    LocalMux I__6946 (
            .O(N__37079),
            .I(n3039));
    Odrv4 I__6945 (
            .O(N__37070),
            .I(n3039));
    Odrv4 I__6944 (
            .O(N__37065),
            .I(n3039));
    CascadeMux I__6943 (
            .O(N__37044),
            .I(N__37040));
    InMux I__6942 (
            .O(N__37043),
            .I(N__37036));
    InMux I__6941 (
            .O(N__37040),
            .I(N__37033));
    InMux I__6940 (
            .O(N__37039),
            .I(N__37030));
    LocalMux I__6939 (
            .O(N__37036),
            .I(N__37025));
    LocalMux I__6938 (
            .O(N__37033),
            .I(N__37025));
    LocalMux I__6937 (
            .O(N__37030),
            .I(N__37022));
    Span4Mux_h I__6936 (
            .O(N__37025),
            .I(N__37019));
    Span12Mux_s4_v I__6935 (
            .O(N__37022),
            .I(N__37016));
    Odrv4 I__6934 (
            .O(N__37019),
            .I(n3123));
    Odrv12 I__6933 (
            .O(N__37016),
            .I(n3123));
    InMux I__6932 (
            .O(N__37011),
            .I(N__37008));
    LocalMux I__6931 (
            .O(N__37008),
            .I(N__37005));
    Span4Mux_v I__6930 (
            .O(N__37005),
            .I(N__37002));
    IoSpan4Mux I__6929 (
            .O(N__37002),
            .I(N__36999));
    IoSpan4Mux I__6928 (
            .O(N__36999),
            .I(N__36996));
    Odrv4 I__6927 (
            .O(N__36996),
            .I(ENCODER0_A_N));
    InMux I__6926 (
            .O(N__36993),
            .I(N__36984));
    InMux I__6925 (
            .O(N__36992),
            .I(N__36984));
    InMux I__6924 (
            .O(N__36991),
            .I(N__36984));
    LocalMux I__6923 (
            .O(N__36984),
            .I(\quad_counter0.a_new_0 ));
    InMux I__6922 (
            .O(N__36981),
            .I(N__36978));
    LocalMux I__6921 (
            .O(N__36978),
            .I(N__36975));
    Span4Mux_v I__6920 (
            .O(N__36975),
            .I(N__36972));
    Odrv4 I__6919 (
            .O(N__36972),
            .I(encoder0_position_scaled_21));
    InMux I__6918 (
            .O(N__36969),
            .I(N__36966));
    LocalMux I__6917 (
            .O(N__36966),
            .I(N__36963));
    Span4Mux_h I__6916 (
            .O(N__36963),
            .I(N__36960));
    Odrv4 I__6915 (
            .O(N__36960),
            .I(encoder0_position_scaled_4));
    InMux I__6914 (
            .O(N__36957),
            .I(N__36954));
    LocalMux I__6913 (
            .O(N__36954),
            .I(N__36951));
    Span4Mux_h I__6912 (
            .O(N__36951),
            .I(N__36948));
    Odrv4 I__6911 (
            .O(N__36948),
            .I(encoder0_position_scaled_5));
    InMux I__6910 (
            .O(N__36945),
            .I(N__36942));
    LocalMux I__6909 (
            .O(N__36942),
            .I(N__36939));
    Span4Mux_h I__6908 (
            .O(N__36939),
            .I(N__36936));
    Odrv4 I__6907 (
            .O(N__36936),
            .I(encoder0_position_scaled_22));
    CascadeMux I__6906 (
            .O(N__36933),
            .I(N__36929));
    CascadeMux I__6905 (
            .O(N__36932),
            .I(N__36926));
    InMux I__6904 (
            .O(N__36929),
            .I(N__36923));
    InMux I__6903 (
            .O(N__36926),
            .I(N__36920));
    LocalMux I__6902 (
            .O(N__36923),
            .I(N__36917));
    LocalMux I__6901 (
            .O(N__36920),
            .I(N__36914));
    Span4Mux_v I__6900 (
            .O(N__36917),
            .I(N__36909));
    Span4Mux_h I__6899 (
            .O(N__36914),
            .I(N__36909));
    Odrv4 I__6898 (
            .O(N__36909),
            .I(n3133));
    CascadeMux I__6897 (
            .O(N__36906),
            .I(N__36902));
    InMux I__6896 (
            .O(N__36905),
            .I(N__36899));
    InMux I__6895 (
            .O(N__36902),
            .I(N__36895));
    LocalMux I__6894 (
            .O(N__36899),
            .I(N__36892));
    InMux I__6893 (
            .O(N__36898),
            .I(N__36889));
    LocalMux I__6892 (
            .O(N__36895),
            .I(N__36886));
    Span4Mux_h I__6891 (
            .O(N__36892),
            .I(N__36883));
    LocalMux I__6890 (
            .O(N__36889),
            .I(n3132));
    Odrv12 I__6889 (
            .O(N__36886),
            .I(n3132));
    Odrv4 I__6888 (
            .O(N__36883),
            .I(n3132));
    CascadeMux I__6887 (
            .O(N__36876),
            .I(N__36871));
    InMux I__6886 (
            .O(N__36875),
            .I(N__36868));
    InMux I__6885 (
            .O(N__36874),
            .I(N__36865));
    InMux I__6884 (
            .O(N__36871),
            .I(N__36862));
    LocalMux I__6883 (
            .O(N__36868),
            .I(N__36859));
    LocalMux I__6882 (
            .O(N__36865),
            .I(N__36856));
    LocalMux I__6881 (
            .O(N__36862),
            .I(N__36853));
    Span4Mux_v I__6880 (
            .O(N__36859),
            .I(N__36850));
    Span4Mux_h I__6879 (
            .O(N__36856),
            .I(N__36845));
    Span4Mux_v I__6878 (
            .O(N__36853),
            .I(N__36845));
    Span4Mux_h I__6877 (
            .O(N__36850),
            .I(N__36842));
    Odrv4 I__6876 (
            .O(N__36845),
            .I(n3129));
    Odrv4 I__6875 (
            .O(N__36842),
            .I(n3129));
    InMux I__6874 (
            .O(N__36837),
            .I(N__36832));
    CascadeMux I__6873 (
            .O(N__36836),
            .I(N__36829));
    InMux I__6872 (
            .O(N__36835),
            .I(N__36826));
    LocalMux I__6871 (
            .O(N__36832),
            .I(N__36823));
    InMux I__6870 (
            .O(N__36829),
            .I(N__36820));
    LocalMux I__6869 (
            .O(N__36826),
            .I(N__36817));
    Span4Mux_h I__6868 (
            .O(N__36823),
            .I(N__36814));
    LocalMux I__6867 (
            .O(N__36820),
            .I(N__36811));
    Span4Mux_v I__6866 (
            .O(N__36817),
            .I(N__36808));
    Odrv4 I__6865 (
            .O(N__36814),
            .I(n3130));
    Odrv12 I__6864 (
            .O(N__36811),
            .I(n3130));
    Odrv4 I__6863 (
            .O(N__36808),
            .I(n3130));
    CascadeMux I__6862 (
            .O(N__36801),
            .I(n11930_cascade_));
    CascadeMux I__6861 (
            .O(N__36798),
            .I(N__36795));
    InMux I__6860 (
            .O(N__36795),
            .I(N__36791));
    InMux I__6859 (
            .O(N__36794),
            .I(N__36788));
    LocalMux I__6858 (
            .O(N__36791),
            .I(N__36784));
    LocalMux I__6857 (
            .O(N__36788),
            .I(N__36781));
    InMux I__6856 (
            .O(N__36787),
            .I(N__36778));
    Span4Mux_v I__6855 (
            .O(N__36784),
            .I(N__36773));
    Span4Mux_h I__6854 (
            .O(N__36781),
            .I(N__36773));
    LocalMux I__6853 (
            .O(N__36778),
            .I(n3131));
    Odrv4 I__6852 (
            .O(N__36773),
            .I(n3131));
    CascadeMux I__6851 (
            .O(N__36768),
            .I(N__36765));
    InMux I__6850 (
            .O(N__36765),
            .I(N__36762));
    LocalMux I__6849 (
            .O(N__36762),
            .I(N__36759));
    Span4Mux_h I__6848 (
            .O(N__36759),
            .I(N__36756));
    Odrv4 I__6847 (
            .O(N__36756),
            .I(n13819));
    InMux I__6846 (
            .O(N__36753),
            .I(\quad_counter0.n13049 ));
    InMux I__6845 (
            .O(N__36750),
            .I(\quad_counter0.n13050 ));
    InMux I__6844 (
            .O(N__36747),
            .I(\quad_counter0.n13051 ));
    InMux I__6843 (
            .O(N__36744),
            .I(\quad_counter0.n13052 ));
    InMux I__6842 (
            .O(N__36741),
            .I(\quad_counter0.n13053 ));
    InMux I__6841 (
            .O(N__36738),
            .I(\quad_counter0.n13054 ));
    InMux I__6840 (
            .O(N__36735),
            .I(\quad_counter0.n13055 ));
    InMux I__6839 (
            .O(N__36732),
            .I(N__36729));
    LocalMux I__6838 (
            .O(N__36729),
            .I(N__36726));
    Span4Mux_v I__6837 (
            .O(N__36726),
            .I(N__36723));
    Odrv4 I__6836 (
            .O(N__36723),
            .I(encoder0_position_scaled_17));
    CascadeMux I__6835 (
            .O(N__36720),
            .I(N__36715));
    InMux I__6834 (
            .O(N__36719),
            .I(N__36712));
    InMux I__6833 (
            .O(N__36718),
            .I(N__36709));
    InMux I__6832 (
            .O(N__36715),
            .I(N__36706));
    LocalMux I__6831 (
            .O(N__36712),
            .I(N__36703));
    LocalMux I__6830 (
            .O(N__36709),
            .I(N__36700));
    LocalMux I__6829 (
            .O(N__36706),
            .I(encoder0_position_14));
    Odrv4 I__6828 (
            .O(N__36703),
            .I(encoder0_position_14));
    Odrv4 I__6827 (
            .O(N__36700),
            .I(encoder0_position_14));
    InMux I__6826 (
            .O(N__36693),
            .I(bfn_9_24_0_));
    InMux I__6825 (
            .O(N__36690),
            .I(\quad_counter0.n13041 ));
    InMux I__6824 (
            .O(N__36687),
            .I(\quad_counter0.n13042 ));
    InMux I__6823 (
            .O(N__36684),
            .I(\quad_counter0.n13043 ));
    InMux I__6822 (
            .O(N__36681),
            .I(\quad_counter0.n13044 ));
    InMux I__6821 (
            .O(N__36678),
            .I(\quad_counter0.n13045 ));
    InMux I__6820 (
            .O(N__36675),
            .I(\quad_counter0.n13046 ));
    InMux I__6819 (
            .O(N__36672),
            .I(\quad_counter0.n13047 ));
    InMux I__6818 (
            .O(N__36669),
            .I(bfn_9_25_0_));
    InMux I__6817 (
            .O(N__36666),
            .I(N__36659));
    InMux I__6816 (
            .O(N__36665),
            .I(N__36659));
    CascadeMux I__6815 (
            .O(N__36664),
            .I(N__36656));
    LocalMux I__6814 (
            .O(N__36659),
            .I(N__36653));
    InMux I__6813 (
            .O(N__36656),
            .I(N__36650));
    Span4Mux_h I__6812 (
            .O(N__36653),
            .I(N__36647));
    LocalMux I__6811 (
            .O(N__36650),
            .I(encoder0_position_8));
    Odrv4 I__6810 (
            .O(N__36647),
            .I(encoder0_position_8));
    InMux I__6809 (
            .O(N__36642),
            .I(bfn_9_23_0_));
    InMux I__6808 (
            .O(N__36639),
            .I(\quad_counter0.n13033 ));
    InMux I__6807 (
            .O(N__36636),
            .I(\quad_counter0.n13034 ));
    InMux I__6806 (
            .O(N__36633),
            .I(N__36627));
    InMux I__6805 (
            .O(N__36632),
            .I(N__36627));
    LocalMux I__6804 (
            .O(N__36627),
            .I(N__36623));
    InMux I__6803 (
            .O(N__36626),
            .I(N__36620));
    Span4Mux_h I__6802 (
            .O(N__36623),
            .I(N__36617));
    LocalMux I__6801 (
            .O(N__36620),
            .I(encoder0_position_11));
    Odrv4 I__6800 (
            .O(N__36617),
            .I(encoder0_position_11));
    InMux I__6799 (
            .O(N__36612),
            .I(\quad_counter0.n13035 ));
    InMux I__6798 (
            .O(N__36609),
            .I(N__36605));
    InMux I__6797 (
            .O(N__36608),
            .I(N__36602));
    LocalMux I__6796 (
            .O(N__36605),
            .I(N__36598));
    LocalMux I__6795 (
            .O(N__36602),
            .I(N__36595));
    CascadeMux I__6794 (
            .O(N__36601),
            .I(N__36592));
    Span4Mux_v I__6793 (
            .O(N__36598),
            .I(N__36589));
    Span4Mux_h I__6792 (
            .O(N__36595),
            .I(N__36586));
    InMux I__6791 (
            .O(N__36592),
            .I(N__36583));
    Span4Mux_h I__6790 (
            .O(N__36589),
            .I(N__36578));
    Span4Mux_v I__6789 (
            .O(N__36586),
            .I(N__36578));
    LocalMux I__6788 (
            .O(N__36583),
            .I(encoder0_position_12));
    Odrv4 I__6787 (
            .O(N__36578),
            .I(encoder0_position_12));
    InMux I__6786 (
            .O(N__36573),
            .I(\quad_counter0.n13036 ));
    InMux I__6785 (
            .O(N__36570),
            .I(N__36566));
    InMux I__6784 (
            .O(N__36569),
            .I(N__36562));
    LocalMux I__6783 (
            .O(N__36566),
            .I(N__36559));
    InMux I__6782 (
            .O(N__36565),
            .I(N__36556));
    LocalMux I__6781 (
            .O(N__36562),
            .I(N__36551));
    Span4Mux_v I__6780 (
            .O(N__36559),
            .I(N__36551));
    LocalMux I__6779 (
            .O(N__36556),
            .I(encoder0_position_13));
    Odrv4 I__6778 (
            .O(N__36551),
            .I(encoder0_position_13));
    InMux I__6777 (
            .O(N__36546),
            .I(\quad_counter0.n13037 ));
    InMux I__6776 (
            .O(N__36543),
            .I(\quad_counter0.n13038 ));
    InMux I__6775 (
            .O(N__36540),
            .I(\quad_counter0.n13039 ));
    InMux I__6774 (
            .O(N__36537),
            .I(N__36533));
    InMux I__6773 (
            .O(N__36536),
            .I(N__36529));
    LocalMux I__6772 (
            .O(N__36533),
            .I(N__36526));
    InMux I__6771 (
            .O(N__36532),
            .I(N__36523));
    LocalMux I__6770 (
            .O(N__36529),
            .I(encoder0_position_0));
    Odrv4 I__6769 (
            .O(N__36526),
            .I(encoder0_position_0));
    LocalMux I__6768 (
            .O(N__36523),
            .I(encoder0_position_0));
    InMux I__6767 (
            .O(N__36516),
            .I(bfn_9_22_0_));
    InMux I__6766 (
            .O(N__36513),
            .I(\quad_counter0.n13025 ));
    InMux I__6765 (
            .O(N__36510),
            .I(\quad_counter0.n13026 ));
    InMux I__6764 (
            .O(N__36507),
            .I(\quad_counter0.n13027 ));
    InMux I__6763 (
            .O(N__36504),
            .I(N__36500));
    InMux I__6762 (
            .O(N__36503),
            .I(N__36496));
    LocalMux I__6761 (
            .O(N__36500),
            .I(N__36493));
    InMux I__6760 (
            .O(N__36499),
            .I(N__36490));
    LocalMux I__6759 (
            .O(N__36496),
            .I(encoder0_position_4));
    Odrv4 I__6758 (
            .O(N__36493),
            .I(encoder0_position_4));
    LocalMux I__6757 (
            .O(N__36490),
            .I(encoder0_position_4));
    InMux I__6756 (
            .O(N__36483),
            .I(\quad_counter0.n13028 ));
    InMux I__6755 (
            .O(N__36480),
            .I(\quad_counter0.n13029 ));
    InMux I__6754 (
            .O(N__36477),
            .I(\quad_counter0.n13030 ));
    InMux I__6753 (
            .O(N__36474),
            .I(\quad_counter0.n13031 ));
    CascadeMux I__6752 (
            .O(N__36471),
            .I(n14558_cascade_));
    CascadeMux I__6751 (
            .O(N__36468),
            .I(N__36465));
    InMux I__6750 (
            .O(N__36465),
            .I(N__36461));
    InMux I__6749 (
            .O(N__36464),
            .I(N__36458));
    LocalMux I__6748 (
            .O(N__36461),
            .I(N__36455));
    LocalMux I__6747 (
            .O(N__36458),
            .I(N__36452));
    Span4Mux_h I__6746 (
            .O(N__36455),
            .I(N__36448));
    Span4Mux_h I__6745 (
            .O(N__36452),
            .I(N__36445));
    InMux I__6744 (
            .O(N__36451),
            .I(N__36442));
    Odrv4 I__6743 (
            .O(N__36448),
            .I(n2019));
    Odrv4 I__6742 (
            .O(N__36445),
            .I(n2019));
    LocalMux I__6741 (
            .O(N__36442),
            .I(n2019));
    InMux I__6740 (
            .O(N__36435),
            .I(N__36432));
    LocalMux I__6739 (
            .O(N__36432),
            .I(N__36429));
    Span4Mux_h I__6738 (
            .O(N__36429),
            .I(N__36426));
    Odrv4 I__6737 (
            .O(N__36426),
            .I(n14564));
    InMux I__6736 (
            .O(N__36423),
            .I(N__36420));
    LocalMux I__6735 (
            .O(N__36420),
            .I(N__36417));
    Odrv4 I__6734 (
            .O(N__36417),
            .I(n1991));
    CascadeMux I__6733 (
            .O(N__36414),
            .I(N__36410));
    CascadeMux I__6732 (
            .O(N__36413),
            .I(N__36407));
    InMux I__6731 (
            .O(N__36410),
            .I(N__36404));
    InMux I__6730 (
            .O(N__36407),
            .I(N__36401));
    LocalMux I__6729 (
            .O(N__36404),
            .I(N__36398));
    LocalMux I__6728 (
            .O(N__36401),
            .I(N__36394));
    Span4Mux_h I__6727 (
            .O(N__36398),
            .I(N__36391));
    InMux I__6726 (
            .O(N__36397),
            .I(N__36388));
    Odrv4 I__6725 (
            .O(N__36394),
            .I(n2023));
    Odrv4 I__6724 (
            .O(N__36391),
            .I(n2023));
    LocalMux I__6723 (
            .O(N__36388),
            .I(n2023));
    InMux I__6722 (
            .O(N__36381),
            .I(N__36378));
    LocalMux I__6721 (
            .O(N__36378),
            .I(N__36375));
    Odrv4 I__6720 (
            .O(N__36375),
            .I(n1994));
    CascadeMux I__6719 (
            .O(N__36372),
            .I(N__36368));
    CascadeMux I__6718 (
            .O(N__36371),
            .I(N__36365));
    InMux I__6717 (
            .O(N__36368),
            .I(N__36362));
    InMux I__6716 (
            .O(N__36365),
            .I(N__36359));
    LocalMux I__6715 (
            .O(N__36362),
            .I(N__36356));
    LocalMux I__6714 (
            .O(N__36359),
            .I(N__36353));
    Span4Mux_h I__6713 (
            .O(N__36356),
            .I(N__36349));
    Span4Mux_h I__6712 (
            .O(N__36353),
            .I(N__36346));
    InMux I__6711 (
            .O(N__36352),
            .I(N__36343));
    Odrv4 I__6710 (
            .O(N__36349),
            .I(n2026));
    Odrv4 I__6709 (
            .O(N__36346),
            .I(n2026));
    LocalMux I__6708 (
            .O(N__36343),
            .I(n2026));
    InMux I__6707 (
            .O(N__36336),
            .I(N__36333));
    LocalMux I__6706 (
            .O(N__36333),
            .I(n1993));
    InMux I__6705 (
            .O(N__36330),
            .I(N__36327));
    LocalMux I__6704 (
            .O(N__36327),
            .I(n1990));
    InMux I__6703 (
            .O(N__36324),
            .I(N__36321));
    LocalMux I__6702 (
            .O(N__36321),
            .I(n1985));
    InMux I__6701 (
            .O(N__36318),
            .I(N__36313));
    InMux I__6700 (
            .O(N__36317),
            .I(N__36308));
    InMux I__6699 (
            .O(N__36316),
            .I(N__36308));
    LocalMux I__6698 (
            .O(N__36313),
            .I(N__36305));
    LocalMux I__6697 (
            .O(N__36308),
            .I(N__36302));
    Odrv4 I__6696 (
            .O(N__36305),
            .I(n2017));
    Odrv12 I__6695 (
            .O(N__36302),
            .I(n2017));
    InMux I__6694 (
            .O(N__36297),
            .I(N__36294));
    LocalMux I__6693 (
            .O(N__36294),
            .I(n1992));
    CascadeMux I__6692 (
            .O(N__36291),
            .I(N__36288));
    InMux I__6691 (
            .O(N__36288),
            .I(N__36285));
    LocalMux I__6690 (
            .O(N__36285),
            .I(N__36282));
    Odrv4 I__6689 (
            .O(N__36282),
            .I(n1997));
    InMux I__6688 (
            .O(N__36279),
            .I(N__36276));
    LocalMux I__6687 (
            .O(N__36276),
            .I(n1987));
    CascadeMux I__6686 (
            .O(N__36273),
            .I(N__36270));
    InMux I__6685 (
            .O(N__36270),
            .I(N__36266));
    InMux I__6684 (
            .O(N__36269),
            .I(N__36263));
    LocalMux I__6683 (
            .O(N__36266),
            .I(N__36260));
    LocalMux I__6682 (
            .O(N__36263),
            .I(N__36256));
    Span4Mux_h I__6681 (
            .O(N__36260),
            .I(N__36253));
    InMux I__6680 (
            .O(N__36259),
            .I(N__36250));
    Odrv4 I__6679 (
            .O(N__36256),
            .I(n2025));
    Odrv4 I__6678 (
            .O(N__36253),
            .I(n2025));
    LocalMux I__6677 (
            .O(N__36250),
            .I(n2025));
    CascadeMux I__6676 (
            .O(N__36243),
            .I(N__36239));
    CascadeMux I__6675 (
            .O(N__36242),
            .I(N__36236));
    InMux I__6674 (
            .O(N__36239),
            .I(N__36233));
    InMux I__6673 (
            .O(N__36236),
            .I(N__36230));
    LocalMux I__6672 (
            .O(N__36233),
            .I(N__36227));
    LocalMux I__6671 (
            .O(N__36230),
            .I(N__36224));
    Span4Mux_h I__6670 (
            .O(N__36227),
            .I(N__36220));
    Span4Mux_h I__6669 (
            .O(N__36224),
            .I(N__36217));
    InMux I__6668 (
            .O(N__36223),
            .I(N__36214));
    Odrv4 I__6667 (
            .O(N__36220),
            .I(n2022));
    Odrv4 I__6666 (
            .O(N__36217),
            .I(n2022));
    LocalMux I__6665 (
            .O(N__36214),
            .I(n2022));
    CascadeMux I__6664 (
            .O(N__36207),
            .I(N__36204));
    InMux I__6663 (
            .O(N__36204),
            .I(N__36200));
    InMux I__6662 (
            .O(N__36203),
            .I(N__36196));
    LocalMux I__6661 (
            .O(N__36200),
            .I(N__36193));
    InMux I__6660 (
            .O(N__36199),
            .I(N__36190));
    LocalMux I__6659 (
            .O(N__36196),
            .I(N__36187));
    Span4Mux_h I__6658 (
            .O(N__36193),
            .I(N__36182));
    LocalMux I__6657 (
            .O(N__36190),
            .I(N__36182));
    Odrv4 I__6656 (
            .O(N__36187),
            .I(n2024));
    Odrv4 I__6655 (
            .O(N__36182),
            .I(n2024));
    CascadeMux I__6654 (
            .O(N__36177),
            .I(n14550_cascade_));
    CascadeMux I__6653 (
            .O(N__36174),
            .I(N__36170));
    CascadeMux I__6652 (
            .O(N__36173),
            .I(N__36167));
    InMux I__6651 (
            .O(N__36170),
            .I(N__36164));
    InMux I__6650 (
            .O(N__36167),
            .I(N__36161));
    LocalMux I__6649 (
            .O(N__36164),
            .I(N__36158));
    LocalMux I__6648 (
            .O(N__36161),
            .I(N__36155));
    Span4Mux_h I__6647 (
            .O(N__36158),
            .I(N__36151));
    Span4Mux_h I__6646 (
            .O(N__36155),
            .I(N__36148));
    InMux I__6645 (
            .O(N__36154),
            .I(N__36145));
    Odrv4 I__6644 (
            .O(N__36151),
            .I(n2029));
    Odrv4 I__6643 (
            .O(N__36148),
            .I(n2029));
    LocalMux I__6642 (
            .O(N__36145),
            .I(n2029));
    CascadeMux I__6641 (
            .O(N__36138),
            .I(n14556_cascade_));
    InMux I__6640 (
            .O(N__36135),
            .I(n12616));
    InMux I__6639 (
            .O(N__36132),
            .I(n12617));
    InMux I__6638 (
            .O(N__36129),
            .I(n12618));
    InMux I__6637 (
            .O(N__36126),
            .I(n12619));
    InMux I__6636 (
            .O(N__36123),
            .I(n12620));
    InMux I__6635 (
            .O(N__36120),
            .I(n12621));
    CascadeMux I__6634 (
            .O(N__36117),
            .I(N__36114));
    InMux I__6633 (
            .O(N__36114),
            .I(N__36111));
    LocalMux I__6632 (
            .O(N__36111),
            .I(N__36108));
    Span4Mux_h I__6631 (
            .O(N__36108),
            .I(N__36105));
    Odrv4 I__6630 (
            .O(N__36105),
            .I(n1986));
    InMux I__6629 (
            .O(N__36102),
            .I(n12622));
    InMux I__6628 (
            .O(N__36099),
            .I(bfn_9_19_0_));
    InMux I__6627 (
            .O(N__36096),
            .I(n12624));
    InMux I__6626 (
            .O(N__36093),
            .I(N__36089));
    InMux I__6625 (
            .O(N__36092),
            .I(N__36086));
    LocalMux I__6624 (
            .O(N__36089),
            .I(N__36081));
    LocalMux I__6623 (
            .O(N__36086),
            .I(N__36081));
    Odrv12 I__6622 (
            .O(N__36081),
            .I(n2016));
    InMux I__6621 (
            .O(N__36078),
            .I(bfn_9_17_0_));
    InMux I__6620 (
            .O(N__36075),
            .I(n12608));
    InMux I__6619 (
            .O(N__36072),
            .I(n12609));
    InMux I__6618 (
            .O(N__36069),
            .I(n12610));
    InMux I__6617 (
            .O(N__36066),
            .I(n12611));
    InMux I__6616 (
            .O(N__36063),
            .I(n12612));
    InMux I__6615 (
            .O(N__36060),
            .I(n12613));
    InMux I__6614 (
            .O(N__36057),
            .I(n12614));
    InMux I__6613 (
            .O(N__36054),
            .I(bfn_9_18_0_));
    InMux I__6612 (
            .O(N__36051),
            .I(N__36048));
    LocalMux I__6611 (
            .O(N__36048),
            .I(N__36044));
    InMux I__6610 (
            .O(N__36047),
            .I(N__36041));
    Sp12to4 I__6609 (
            .O(N__36044),
            .I(N__36036));
    LocalMux I__6608 (
            .O(N__36041),
            .I(N__36036));
    Span12Mux_s5_v I__6607 (
            .O(N__36036),
            .I(N__36032));
    InMux I__6606 (
            .O(N__36035),
            .I(N__36029));
    Odrv12 I__6605 (
            .O(N__36032),
            .I(n3211));
    LocalMux I__6604 (
            .O(N__36029),
            .I(n3211));
    InMux I__6603 (
            .O(N__36024),
            .I(N__36021));
    LocalMux I__6602 (
            .O(N__36021),
            .I(n3278));
    InMux I__6601 (
            .O(N__36018),
            .I(bfn_7_32_0_));
    InMux I__6600 (
            .O(N__36015),
            .I(N__36010));
    InMux I__6599 (
            .O(N__36014),
            .I(N__36007));
    CascadeMux I__6598 (
            .O(N__36013),
            .I(N__36004));
    LocalMux I__6597 (
            .O(N__36010),
            .I(N__36001));
    LocalMux I__6596 (
            .O(N__36007),
            .I(N__35998));
    InMux I__6595 (
            .O(N__36004),
            .I(N__35995));
    Span4Mux_s1_v I__6594 (
            .O(N__36001),
            .I(N__35992));
    Span4Mux_s3_v I__6593 (
            .O(N__35998),
            .I(N__35987));
    LocalMux I__6592 (
            .O(N__35995),
            .I(N__35987));
    Odrv4 I__6591 (
            .O(N__35992),
            .I(n3210));
    Odrv4 I__6590 (
            .O(N__35987),
            .I(n3210));
    InMux I__6589 (
            .O(N__35982),
            .I(N__35979));
    LocalMux I__6588 (
            .O(N__35979),
            .I(n3277));
    InMux I__6587 (
            .O(N__35976),
            .I(n12931));
    InMux I__6586 (
            .O(N__35973),
            .I(N__35970));
    LocalMux I__6585 (
            .O(N__35970),
            .I(N__35965));
    InMux I__6584 (
            .O(N__35969),
            .I(N__35960));
    InMux I__6583 (
            .O(N__35968),
            .I(N__35960));
    Odrv12 I__6582 (
            .O(N__35965),
            .I(n3209));
    LocalMux I__6581 (
            .O(N__35960),
            .I(n3209));
    InMux I__6580 (
            .O(N__35955),
            .I(N__35952));
    LocalMux I__6579 (
            .O(N__35952),
            .I(N__35949));
    Span4Mux_v I__6578 (
            .O(N__35949),
            .I(N__35946));
    Odrv4 I__6577 (
            .O(N__35946),
            .I(n3276));
    InMux I__6576 (
            .O(N__35943),
            .I(n12932));
    InMux I__6575 (
            .O(N__35940),
            .I(N__35937));
    LocalMux I__6574 (
            .O(N__35937),
            .I(N__35934));
    Span4Mux_v I__6573 (
            .O(N__35934),
            .I(N__35931));
    Odrv4 I__6572 (
            .O(N__35931),
            .I(n3275));
    InMux I__6571 (
            .O(N__35928),
            .I(n12933));
    InMux I__6570 (
            .O(N__35925),
            .I(N__35922));
    LocalMux I__6569 (
            .O(N__35922),
            .I(N__35919));
    Span4Mux_s1_v I__6568 (
            .O(N__35919),
            .I(N__35914));
    InMux I__6567 (
            .O(N__35918),
            .I(N__35909));
    InMux I__6566 (
            .O(N__35917),
            .I(N__35909));
    Span4Mux_v I__6565 (
            .O(N__35914),
            .I(N__35906));
    LocalMux I__6564 (
            .O(N__35909),
            .I(N__35903));
    Odrv4 I__6563 (
            .O(N__35906),
            .I(n3207));
    Odrv4 I__6562 (
            .O(N__35903),
            .I(n3207));
    InMux I__6561 (
            .O(N__35898),
            .I(N__35895));
    LocalMux I__6560 (
            .O(N__35895),
            .I(N__35892));
    Span4Mux_v I__6559 (
            .O(N__35892),
            .I(N__35889));
    Span4Mux_v I__6558 (
            .O(N__35889),
            .I(N__35886));
    Odrv4 I__6557 (
            .O(N__35886),
            .I(n3274));
    InMux I__6556 (
            .O(N__35883),
            .I(n12934));
    InMux I__6555 (
            .O(N__35880),
            .I(N__35876));
    InMux I__6554 (
            .O(N__35879),
            .I(N__35872));
    LocalMux I__6553 (
            .O(N__35876),
            .I(N__35869));
    InMux I__6552 (
            .O(N__35875),
            .I(N__35866));
    LocalMux I__6551 (
            .O(N__35872),
            .I(N__35863));
    Span4Mux_v I__6550 (
            .O(N__35869),
            .I(N__35860));
    LocalMux I__6549 (
            .O(N__35866),
            .I(N__35857));
    Odrv12 I__6548 (
            .O(N__35863),
            .I(n3206));
    Odrv4 I__6547 (
            .O(N__35860),
            .I(n3206));
    Odrv4 I__6546 (
            .O(N__35857),
            .I(n3206));
    InMux I__6545 (
            .O(N__35850),
            .I(N__35847));
    LocalMux I__6544 (
            .O(N__35847),
            .I(n3273));
    InMux I__6543 (
            .O(N__35844),
            .I(n12935));
    InMux I__6542 (
            .O(N__35841),
            .I(N__35838));
    LocalMux I__6541 (
            .O(N__35838),
            .I(N__35835));
    Span4Mux_v I__6540 (
            .O(N__35835),
            .I(N__35830));
    InMux I__6539 (
            .O(N__35834),
            .I(N__35825));
    InMux I__6538 (
            .O(N__35833),
            .I(N__35825));
    Odrv4 I__6537 (
            .O(N__35830),
            .I(n3205));
    LocalMux I__6536 (
            .O(N__35825),
            .I(n3205));
    InMux I__6535 (
            .O(N__35820),
            .I(N__35817));
    LocalMux I__6534 (
            .O(N__35817),
            .I(N__35814));
    Span4Mux_h I__6533 (
            .O(N__35814),
            .I(N__35811));
    Span4Mux_v I__6532 (
            .O(N__35811),
            .I(N__35808));
    Odrv4 I__6531 (
            .O(N__35808),
            .I(n3272));
    InMux I__6530 (
            .O(N__35805),
            .I(n12936));
    InMux I__6529 (
            .O(N__35802),
            .I(N__35798));
    InMux I__6528 (
            .O(N__35801),
            .I(N__35795));
    LocalMux I__6527 (
            .O(N__35798),
            .I(N__35792));
    LocalMux I__6526 (
            .O(N__35795),
            .I(N__35789));
    Span4Mux_s1_v I__6525 (
            .O(N__35792),
            .I(N__35786));
    Odrv12 I__6524 (
            .O(N__35789),
            .I(n15450));
    Odrv4 I__6523 (
            .O(N__35786),
            .I(n15450));
    CascadeMux I__6522 (
            .O(N__35781),
            .I(N__35778));
    InMux I__6521 (
            .O(N__35778),
            .I(N__35775));
    LocalMux I__6520 (
            .O(N__35775),
            .I(N__35771));
    InMux I__6519 (
            .O(N__35774),
            .I(N__35768));
    Span4Mux_v I__6518 (
            .O(N__35771),
            .I(N__35765));
    LocalMux I__6517 (
            .O(N__35768),
            .I(N__35762));
    Odrv4 I__6516 (
            .O(N__35765),
            .I(n3204));
    Odrv4 I__6515 (
            .O(N__35762),
            .I(n3204));
    InMux I__6514 (
            .O(N__35757),
            .I(n12937));
    InMux I__6513 (
            .O(N__35754),
            .I(N__35751));
    LocalMux I__6512 (
            .O(N__35751),
            .I(N__35748));
    Span4Mux_v I__6511 (
            .O(N__35748),
            .I(N__35745));
    Span4Mux_v I__6510 (
            .O(N__35745),
            .I(N__35742));
    Odrv4 I__6509 (
            .O(N__35742),
            .I(n14873));
    InMux I__6508 (
            .O(N__35739),
            .I(N__35736));
    LocalMux I__6507 (
            .O(N__35736),
            .I(N__35732));
    InMux I__6506 (
            .O(N__35735),
            .I(N__35729));
    Span4Mux_h I__6505 (
            .O(N__35732),
            .I(N__35726));
    LocalMux I__6504 (
            .O(N__35729),
            .I(N__35723));
    Odrv4 I__6503 (
            .O(N__35726),
            .I(n3218));
    Odrv12 I__6502 (
            .O(N__35723),
            .I(n3218));
    InMux I__6501 (
            .O(N__35718),
            .I(N__35715));
    LocalMux I__6500 (
            .O(N__35715),
            .I(n3285));
    InMux I__6499 (
            .O(N__35712),
            .I(n12923));
    CascadeMux I__6498 (
            .O(N__35709),
            .I(N__35706));
    InMux I__6497 (
            .O(N__35706),
            .I(N__35701));
    InMux I__6496 (
            .O(N__35705),
            .I(N__35698));
    InMux I__6495 (
            .O(N__35704),
            .I(N__35695));
    LocalMux I__6494 (
            .O(N__35701),
            .I(N__35692));
    LocalMux I__6493 (
            .O(N__35698),
            .I(N__35689));
    LocalMux I__6492 (
            .O(N__35695),
            .I(N__35686));
    Odrv4 I__6491 (
            .O(N__35692),
            .I(n3217));
    Odrv4 I__6490 (
            .O(N__35689),
            .I(n3217));
    Odrv4 I__6489 (
            .O(N__35686),
            .I(n3217));
    InMux I__6488 (
            .O(N__35679),
            .I(N__35676));
    LocalMux I__6487 (
            .O(N__35676),
            .I(n3284));
    InMux I__6486 (
            .O(N__35673),
            .I(n12924));
    InMux I__6485 (
            .O(N__35670),
            .I(N__35667));
    LocalMux I__6484 (
            .O(N__35667),
            .I(N__35663));
    InMux I__6483 (
            .O(N__35666),
            .I(N__35660));
    Span4Mux_v I__6482 (
            .O(N__35663),
            .I(N__35656));
    LocalMux I__6481 (
            .O(N__35660),
            .I(N__35653));
    InMux I__6480 (
            .O(N__35659),
            .I(N__35650));
    Odrv4 I__6479 (
            .O(N__35656),
            .I(n3216));
    Odrv12 I__6478 (
            .O(N__35653),
            .I(n3216));
    LocalMux I__6477 (
            .O(N__35650),
            .I(n3216));
    InMux I__6476 (
            .O(N__35643),
            .I(N__35640));
    LocalMux I__6475 (
            .O(N__35640),
            .I(n3283));
    InMux I__6474 (
            .O(N__35637),
            .I(n12925));
    CascadeMux I__6473 (
            .O(N__35634),
            .I(N__35631));
    InMux I__6472 (
            .O(N__35631),
            .I(N__35627));
    InMux I__6471 (
            .O(N__35630),
            .I(N__35624));
    LocalMux I__6470 (
            .O(N__35627),
            .I(N__35619));
    LocalMux I__6469 (
            .O(N__35624),
            .I(N__35619));
    Span4Mux_s3_v I__6468 (
            .O(N__35619),
            .I(N__35615));
    InMux I__6467 (
            .O(N__35618),
            .I(N__35612));
    Odrv4 I__6466 (
            .O(N__35615),
            .I(n3215));
    LocalMux I__6465 (
            .O(N__35612),
            .I(n3215));
    InMux I__6464 (
            .O(N__35607),
            .I(N__35604));
    LocalMux I__6463 (
            .O(N__35604),
            .I(n3282));
    InMux I__6462 (
            .O(N__35601),
            .I(n12926));
    InMux I__6461 (
            .O(N__35598),
            .I(N__35594));
    InMux I__6460 (
            .O(N__35597),
            .I(N__35591));
    LocalMux I__6459 (
            .O(N__35594),
            .I(N__35588));
    LocalMux I__6458 (
            .O(N__35591),
            .I(N__35585));
    Span4Mux_v I__6457 (
            .O(N__35588),
            .I(N__35582));
    Odrv12 I__6456 (
            .O(N__35585),
            .I(n3214));
    Odrv4 I__6455 (
            .O(N__35582),
            .I(n3214));
    InMux I__6454 (
            .O(N__35577),
            .I(N__35574));
    LocalMux I__6453 (
            .O(N__35574),
            .I(n3281));
    InMux I__6452 (
            .O(N__35571),
            .I(n12927));
    InMux I__6451 (
            .O(N__35568),
            .I(N__35564));
    InMux I__6450 (
            .O(N__35567),
            .I(N__35561));
    LocalMux I__6449 (
            .O(N__35564),
            .I(N__35557));
    LocalMux I__6448 (
            .O(N__35561),
            .I(N__35554));
    InMux I__6447 (
            .O(N__35560),
            .I(N__35551));
    Span4Mux_s1_v I__6446 (
            .O(N__35557),
            .I(N__35546));
    Span4Mux_h I__6445 (
            .O(N__35554),
            .I(N__35546));
    LocalMux I__6444 (
            .O(N__35551),
            .I(N__35543));
    Odrv4 I__6443 (
            .O(N__35546),
            .I(n3213));
    Odrv4 I__6442 (
            .O(N__35543),
            .I(n3213));
    CascadeMux I__6441 (
            .O(N__35538),
            .I(N__35535));
    InMux I__6440 (
            .O(N__35535),
            .I(N__35532));
    LocalMux I__6439 (
            .O(N__35532),
            .I(n3280));
    InMux I__6438 (
            .O(N__35529),
            .I(n12928));
    InMux I__6437 (
            .O(N__35526),
            .I(N__35521));
    InMux I__6436 (
            .O(N__35525),
            .I(N__35518));
    InMux I__6435 (
            .O(N__35524),
            .I(N__35515));
    LocalMux I__6434 (
            .O(N__35521),
            .I(N__35512));
    LocalMux I__6433 (
            .O(N__35518),
            .I(N__35509));
    LocalMux I__6432 (
            .O(N__35515),
            .I(N__35506));
    Span4Mux_s2_v I__6431 (
            .O(N__35512),
            .I(N__35503));
    Span12Mux_s4_v I__6430 (
            .O(N__35509),
            .I(N__35500));
    Span4Mux_h I__6429 (
            .O(N__35506),
            .I(N__35497));
    Odrv4 I__6428 (
            .O(N__35503),
            .I(n3212));
    Odrv12 I__6427 (
            .O(N__35500),
            .I(n3212));
    Odrv4 I__6426 (
            .O(N__35497),
            .I(n3212));
    InMux I__6425 (
            .O(N__35490),
            .I(N__35487));
    LocalMux I__6424 (
            .O(N__35487),
            .I(n3279));
    InMux I__6423 (
            .O(N__35484),
            .I(n12929));
    InMux I__6422 (
            .O(N__35481),
            .I(N__35478));
    LocalMux I__6421 (
            .O(N__35478),
            .I(N__35474));
    InMux I__6420 (
            .O(N__35477),
            .I(N__35471));
    Span4Mux_v I__6419 (
            .O(N__35474),
            .I(N__35465));
    LocalMux I__6418 (
            .O(N__35471),
            .I(N__35465));
    InMux I__6417 (
            .O(N__35470),
            .I(N__35462));
    Odrv4 I__6416 (
            .O(N__35465),
            .I(n3226));
    LocalMux I__6415 (
            .O(N__35462),
            .I(n3226));
    CascadeMux I__6414 (
            .O(N__35457),
            .I(N__35454));
    InMux I__6413 (
            .O(N__35454),
            .I(N__35451));
    LocalMux I__6412 (
            .O(N__35451),
            .I(N__35448));
    Span4Mux_h I__6411 (
            .O(N__35448),
            .I(N__35445));
    Span4Mux_v I__6410 (
            .O(N__35445),
            .I(N__35442));
    Odrv4 I__6409 (
            .O(N__35442),
            .I(n3293));
    InMux I__6408 (
            .O(N__35439),
            .I(n12915));
    InMux I__6407 (
            .O(N__35436),
            .I(N__35432));
    InMux I__6406 (
            .O(N__35435),
            .I(N__35429));
    LocalMux I__6405 (
            .O(N__35432),
            .I(N__35426));
    LocalMux I__6404 (
            .O(N__35429),
            .I(N__35423));
    Span4Mux_s3_v I__6403 (
            .O(N__35426),
            .I(N__35420));
    Odrv4 I__6402 (
            .O(N__35423),
            .I(n3225));
    Odrv4 I__6401 (
            .O(N__35420),
            .I(n3225));
    InMux I__6400 (
            .O(N__35415),
            .I(N__35412));
    LocalMux I__6399 (
            .O(N__35412),
            .I(N__35409));
    Span4Mux_v I__6398 (
            .O(N__35409),
            .I(N__35406));
    Odrv4 I__6397 (
            .O(N__35406),
            .I(n3292));
    InMux I__6396 (
            .O(N__35403),
            .I(n12916));
    InMux I__6395 (
            .O(N__35400),
            .I(N__35396));
    InMux I__6394 (
            .O(N__35399),
            .I(N__35393));
    LocalMux I__6393 (
            .O(N__35396),
            .I(N__35389));
    LocalMux I__6392 (
            .O(N__35393),
            .I(N__35386));
    InMux I__6391 (
            .O(N__35392),
            .I(N__35383));
    Odrv4 I__6390 (
            .O(N__35389),
            .I(n3224));
    Odrv4 I__6389 (
            .O(N__35386),
            .I(n3224));
    LocalMux I__6388 (
            .O(N__35383),
            .I(n3224));
    InMux I__6387 (
            .O(N__35376),
            .I(N__35373));
    LocalMux I__6386 (
            .O(N__35373),
            .I(N__35370));
    Span4Mux_v I__6385 (
            .O(N__35370),
            .I(N__35367));
    Span4Mux_v I__6384 (
            .O(N__35367),
            .I(N__35364));
    Odrv4 I__6383 (
            .O(N__35364),
            .I(n3291));
    InMux I__6382 (
            .O(N__35361),
            .I(n12917));
    InMux I__6381 (
            .O(N__35358),
            .I(N__35354));
    InMux I__6380 (
            .O(N__35357),
            .I(N__35351));
    LocalMux I__6379 (
            .O(N__35354),
            .I(N__35345));
    LocalMux I__6378 (
            .O(N__35351),
            .I(N__35345));
    InMux I__6377 (
            .O(N__35350),
            .I(N__35342));
    Odrv4 I__6376 (
            .O(N__35345),
            .I(n3223));
    LocalMux I__6375 (
            .O(N__35342),
            .I(n3223));
    InMux I__6374 (
            .O(N__35337),
            .I(N__35334));
    LocalMux I__6373 (
            .O(N__35334),
            .I(n3290));
    InMux I__6372 (
            .O(N__35331),
            .I(n12918));
    InMux I__6371 (
            .O(N__35328),
            .I(N__35325));
    LocalMux I__6370 (
            .O(N__35325),
            .I(N__35322));
    Span4Mux_s3_v I__6369 (
            .O(N__35322),
            .I(N__35318));
    InMux I__6368 (
            .O(N__35321),
            .I(N__35315));
    Odrv4 I__6367 (
            .O(N__35318),
            .I(n3222));
    LocalMux I__6366 (
            .O(N__35315),
            .I(n3222));
    InMux I__6365 (
            .O(N__35310),
            .I(N__35307));
    LocalMux I__6364 (
            .O(N__35307),
            .I(N__35304));
    Span4Mux_h I__6363 (
            .O(N__35304),
            .I(N__35301));
    Odrv4 I__6362 (
            .O(N__35301),
            .I(n3289));
    InMux I__6361 (
            .O(N__35298),
            .I(n12919));
    CascadeMux I__6360 (
            .O(N__35295),
            .I(N__35292));
    InMux I__6359 (
            .O(N__35292),
            .I(N__35288));
    InMux I__6358 (
            .O(N__35291),
            .I(N__35285));
    LocalMux I__6357 (
            .O(N__35288),
            .I(N__35282));
    LocalMux I__6356 (
            .O(N__35285),
            .I(n3221));
    Odrv4 I__6355 (
            .O(N__35282),
            .I(n3221));
    InMux I__6354 (
            .O(N__35277),
            .I(N__35274));
    LocalMux I__6353 (
            .O(N__35274),
            .I(N__35271));
    Odrv12 I__6352 (
            .O(N__35271),
            .I(n3288));
    InMux I__6351 (
            .O(N__35268),
            .I(n12920));
    InMux I__6350 (
            .O(N__35265),
            .I(N__35262));
    LocalMux I__6349 (
            .O(N__35262),
            .I(N__35257));
    InMux I__6348 (
            .O(N__35261),
            .I(N__35252));
    InMux I__6347 (
            .O(N__35260),
            .I(N__35252));
    Odrv4 I__6346 (
            .O(N__35257),
            .I(n3220));
    LocalMux I__6345 (
            .O(N__35252),
            .I(n3220));
    CascadeMux I__6344 (
            .O(N__35247),
            .I(N__35244));
    InMux I__6343 (
            .O(N__35244),
            .I(N__35241));
    LocalMux I__6342 (
            .O(N__35241),
            .I(N__35238));
    Odrv12 I__6341 (
            .O(N__35238),
            .I(n3287));
    InMux I__6340 (
            .O(N__35235),
            .I(n12921));
    InMux I__6339 (
            .O(N__35232),
            .I(N__35228));
    InMux I__6338 (
            .O(N__35231),
            .I(N__35225));
    LocalMux I__6337 (
            .O(N__35228),
            .I(N__35222));
    LocalMux I__6336 (
            .O(N__35225),
            .I(N__35218));
    Span4Mux_s3_v I__6335 (
            .O(N__35222),
            .I(N__35215));
    InMux I__6334 (
            .O(N__35221),
            .I(N__35212));
    Odrv4 I__6333 (
            .O(N__35218),
            .I(n3219));
    Odrv4 I__6332 (
            .O(N__35215),
            .I(n3219));
    LocalMux I__6331 (
            .O(N__35212),
            .I(n3219));
    InMux I__6330 (
            .O(N__35205),
            .I(N__35202));
    LocalMux I__6329 (
            .O(N__35202),
            .I(N__35199));
    Span4Mux_v I__6328 (
            .O(N__35199),
            .I(N__35196));
    Odrv4 I__6327 (
            .O(N__35196),
            .I(n3286));
    InMux I__6326 (
            .O(N__35193),
            .I(bfn_7_31_0_));
    InMux I__6325 (
            .O(N__35190),
            .I(N__35187));
    LocalMux I__6324 (
            .O(N__35187),
            .I(N__35184));
    Span4Mux_h I__6323 (
            .O(N__35184),
            .I(N__35181));
    Odrv4 I__6322 (
            .O(N__35181),
            .I(n3301));
    InMux I__6321 (
            .O(N__35178),
            .I(n12907));
    InMux I__6320 (
            .O(N__35175),
            .I(N__35171));
    InMux I__6319 (
            .O(N__35174),
            .I(N__35168));
    LocalMux I__6318 (
            .O(N__35171),
            .I(n3233));
    LocalMux I__6317 (
            .O(N__35168),
            .I(n3233));
    InMux I__6316 (
            .O(N__35163),
            .I(N__35160));
    LocalMux I__6315 (
            .O(N__35160),
            .I(n3300));
    InMux I__6314 (
            .O(N__35157),
            .I(n12908));
    InMux I__6313 (
            .O(N__35154),
            .I(N__35151));
    LocalMux I__6312 (
            .O(N__35151),
            .I(N__35147));
    InMux I__6311 (
            .O(N__35150),
            .I(N__35144));
    Odrv12 I__6310 (
            .O(N__35147),
            .I(n3232));
    LocalMux I__6309 (
            .O(N__35144),
            .I(n3232));
    InMux I__6308 (
            .O(N__35139),
            .I(N__35136));
    LocalMux I__6307 (
            .O(N__35136),
            .I(N__35133));
    Odrv4 I__6306 (
            .O(N__35133),
            .I(n3299));
    InMux I__6305 (
            .O(N__35130),
            .I(n12909));
    InMux I__6304 (
            .O(N__35127),
            .I(N__35122));
    InMux I__6303 (
            .O(N__35126),
            .I(N__35119));
    InMux I__6302 (
            .O(N__35125),
            .I(N__35116));
    LocalMux I__6301 (
            .O(N__35122),
            .I(n3231));
    LocalMux I__6300 (
            .O(N__35119),
            .I(n3231));
    LocalMux I__6299 (
            .O(N__35116),
            .I(n3231));
    InMux I__6298 (
            .O(N__35109),
            .I(n12910));
    InMux I__6297 (
            .O(N__35106),
            .I(N__35103));
    LocalMux I__6296 (
            .O(N__35103),
            .I(n3298));
    InMux I__6295 (
            .O(N__35100),
            .I(N__35095));
    InMux I__6294 (
            .O(N__35099),
            .I(N__35092));
    InMux I__6293 (
            .O(N__35098),
            .I(N__35089));
    LocalMux I__6292 (
            .O(N__35095),
            .I(N__35086));
    LocalMux I__6291 (
            .O(N__35092),
            .I(n3230));
    LocalMux I__6290 (
            .O(N__35089),
            .I(n3230));
    Odrv4 I__6289 (
            .O(N__35086),
            .I(n3230));
    InMux I__6288 (
            .O(N__35079),
            .I(N__35076));
    LocalMux I__6287 (
            .O(N__35076),
            .I(n15097));
    InMux I__6286 (
            .O(N__35073),
            .I(n12911));
    CascadeMux I__6285 (
            .O(N__35070),
            .I(N__35066));
    InMux I__6284 (
            .O(N__35069),
            .I(N__35063));
    InMux I__6283 (
            .O(N__35066),
            .I(N__35060));
    LocalMux I__6282 (
            .O(N__35063),
            .I(n3229));
    LocalMux I__6281 (
            .O(N__35060),
            .I(n3229));
    InMux I__6280 (
            .O(N__35055),
            .I(N__35052));
    LocalMux I__6279 (
            .O(N__35052),
            .I(n3296));
    InMux I__6278 (
            .O(N__35049),
            .I(n12912));
    InMux I__6277 (
            .O(N__35046),
            .I(N__35043));
    LocalMux I__6276 (
            .O(N__35043),
            .I(N__35038));
    InMux I__6275 (
            .O(N__35042),
            .I(N__35035));
    InMux I__6274 (
            .O(N__35041),
            .I(N__35032));
    Odrv4 I__6273 (
            .O(N__35038),
            .I(n3228));
    LocalMux I__6272 (
            .O(N__35035),
            .I(n3228));
    LocalMux I__6271 (
            .O(N__35032),
            .I(n3228));
    InMux I__6270 (
            .O(N__35025),
            .I(N__35022));
    LocalMux I__6269 (
            .O(N__35022),
            .I(n3295));
    InMux I__6268 (
            .O(N__35019),
            .I(n12913));
    InMux I__6267 (
            .O(N__35016),
            .I(N__35012));
    InMux I__6266 (
            .O(N__35015),
            .I(N__35009));
    LocalMux I__6265 (
            .O(N__35012),
            .I(N__35005));
    LocalMux I__6264 (
            .O(N__35009),
            .I(N__35002));
    InMux I__6263 (
            .O(N__35008),
            .I(N__34999));
    Odrv4 I__6262 (
            .O(N__35005),
            .I(n3227));
    Odrv12 I__6261 (
            .O(N__35002),
            .I(n3227));
    LocalMux I__6260 (
            .O(N__34999),
            .I(n3227));
    CascadeMux I__6259 (
            .O(N__34992),
            .I(N__34989));
    InMux I__6258 (
            .O(N__34989),
            .I(N__34986));
    LocalMux I__6257 (
            .O(N__34986),
            .I(N__34983));
    Span4Mux_h I__6256 (
            .O(N__34983),
            .I(N__34980));
    Span4Mux_v I__6255 (
            .O(N__34980),
            .I(N__34977));
    Odrv4 I__6254 (
            .O(N__34977),
            .I(n3294));
    InMux I__6253 (
            .O(N__34974),
            .I(bfn_7_30_0_));
    CascadeMux I__6252 (
            .O(N__34971),
            .I(N__34968));
    InMux I__6251 (
            .O(N__34968),
            .I(N__34965));
    LocalMux I__6250 (
            .O(N__34965),
            .I(N__34962));
    Span4Mux_v I__6249 (
            .O(N__34962),
            .I(N__34959));
    Odrv4 I__6248 (
            .O(N__34959),
            .I(n3080));
    InMux I__6247 (
            .O(N__34956),
            .I(N__34953));
    LocalMux I__6246 (
            .O(N__34953),
            .I(N__34949));
    InMux I__6245 (
            .O(N__34952),
            .I(N__34945));
    Span4Mux_v I__6244 (
            .O(N__34949),
            .I(N__34942));
    InMux I__6243 (
            .O(N__34948),
            .I(N__34939));
    LocalMux I__6242 (
            .O(N__34945),
            .I(n3112));
    Odrv4 I__6241 (
            .O(N__34942),
            .I(n3112));
    LocalMux I__6240 (
            .O(N__34939),
            .I(n3112));
    InMux I__6239 (
            .O(N__34932),
            .I(N__34929));
    LocalMux I__6238 (
            .O(N__34929),
            .I(N__34926));
    Span4Mux_h I__6237 (
            .O(N__34926),
            .I(N__34923));
    Odrv4 I__6236 (
            .O(N__34923),
            .I(n3192));
    CascadeMux I__6235 (
            .O(N__34920),
            .I(N__34917));
    InMux I__6234 (
            .O(N__34917),
            .I(N__34913));
    InMux I__6233 (
            .O(N__34916),
            .I(N__34910));
    LocalMux I__6232 (
            .O(N__34913),
            .I(N__34907));
    LocalMux I__6231 (
            .O(N__34910),
            .I(N__34903));
    Span4Mux_v I__6230 (
            .O(N__34907),
            .I(N__34900));
    InMux I__6229 (
            .O(N__34906),
            .I(N__34897));
    Odrv4 I__6228 (
            .O(N__34903),
            .I(n3125));
    Odrv4 I__6227 (
            .O(N__34900),
            .I(n3125));
    LocalMux I__6226 (
            .O(N__34897),
            .I(n3125));
    CascadeMux I__6225 (
            .O(N__34890),
            .I(N__34887));
    InMux I__6224 (
            .O(N__34887),
            .I(N__34884));
    LocalMux I__6223 (
            .O(N__34884),
            .I(N__34881));
    Span4Mux_h I__6222 (
            .O(N__34881),
            .I(N__34878));
    Odrv4 I__6221 (
            .O(N__34878),
            .I(n3196));
    InMux I__6220 (
            .O(N__34875),
            .I(N__34871));
    InMux I__6219 (
            .O(N__34874),
            .I(N__34868));
    LocalMux I__6218 (
            .O(N__34871),
            .I(N__34865));
    LocalMux I__6217 (
            .O(N__34868),
            .I(N__34860));
    Span4Mux_h I__6216 (
            .O(N__34865),
            .I(N__34860));
    Span4Mux_h I__6215 (
            .O(N__34860),
            .I(N__34857));
    Odrv4 I__6214 (
            .O(N__34857),
            .I(\debounce.reg_A_0 ));
    InMux I__6213 (
            .O(N__34854),
            .I(N__34850));
    CascadeMux I__6212 (
            .O(N__34853),
            .I(N__34847));
    LocalMux I__6211 (
            .O(N__34850),
            .I(N__34844));
    InMux I__6210 (
            .O(N__34847),
            .I(N__34841));
    Span4Mux_s3_h I__6209 (
            .O(N__34844),
            .I(N__34838));
    LocalMux I__6208 (
            .O(N__34841),
            .I(N__34835));
    Span4Mux_v I__6207 (
            .O(N__34838),
            .I(N__34832));
    Span4Mux_h I__6206 (
            .O(N__34835),
            .I(N__34829));
    Odrv4 I__6205 (
            .O(N__34832),
            .I(reg_B_0));
    Odrv4 I__6204 (
            .O(N__34829),
            .I(reg_B_0));
    InMux I__6203 (
            .O(N__34824),
            .I(N__34820));
    InMux I__6202 (
            .O(N__34823),
            .I(N__34817));
    LocalMux I__6201 (
            .O(N__34820),
            .I(N__34814));
    LocalMux I__6200 (
            .O(N__34817),
            .I(\debounce.reg_A_1 ));
    Odrv12 I__6199 (
            .O(N__34814),
            .I(\debounce.reg_A_1 ));
    CascadeMux I__6198 (
            .O(N__34809),
            .I(N__34806));
    InMux I__6197 (
            .O(N__34806),
            .I(N__34803));
    LocalMux I__6196 (
            .O(N__34803),
            .I(N__34800));
    Span4Mux_v I__6195 (
            .O(N__34800),
            .I(N__34797));
    Odrv4 I__6194 (
            .O(N__34797),
            .I(\debounce.n6 ));
    InMux I__6193 (
            .O(N__34794),
            .I(N__34791));
    LocalMux I__6192 (
            .O(N__34791),
            .I(N__34788));
    Span4Mux_h I__6191 (
            .O(N__34788),
            .I(N__34785));
    Odrv4 I__6190 (
            .O(N__34785),
            .I(n3185));
    CascadeMux I__6189 (
            .O(N__34782),
            .I(N__34777));
    InMux I__6188 (
            .O(N__34781),
            .I(N__34774));
    InMux I__6187 (
            .O(N__34780),
            .I(N__34771));
    InMux I__6186 (
            .O(N__34777),
            .I(N__34768));
    LocalMux I__6185 (
            .O(N__34774),
            .I(N__34765));
    LocalMux I__6184 (
            .O(N__34771),
            .I(N__34762));
    LocalMux I__6183 (
            .O(N__34768),
            .I(N__34759));
    Span4Mux_h I__6182 (
            .O(N__34765),
            .I(N__34752));
    Span4Mux_v I__6181 (
            .O(N__34762),
            .I(N__34752));
    Span4Mux_v I__6180 (
            .O(N__34759),
            .I(N__34752));
    Odrv4 I__6179 (
            .O(N__34752),
            .I(n3118));
    CascadeMux I__6178 (
            .O(N__34749),
            .I(N__34746));
    InMux I__6177 (
            .O(N__34746),
            .I(N__34743));
    LocalMux I__6176 (
            .O(N__34743),
            .I(N__34740));
    Span4Mux_h I__6175 (
            .O(N__34740),
            .I(N__34737));
    Odrv4 I__6174 (
            .O(N__34737),
            .I(n3197));
    CascadeMux I__6173 (
            .O(N__34734),
            .I(n3229_cascade_));
    CascadeMux I__6172 (
            .O(N__34731),
            .I(N__34722));
    CascadeMux I__6171 (
            .O(N__34730),
            .I(N__34717));
    CascadeMux I__6170 (
            .O(N__34729),
            .I(N__34712));
    CascadeMux I__6169 (
            .O(N__34728),
            .I(N__34709));
    CascadeMux I__6168 (
            .O(N__34727),
            .I(N__34704));
    InMux I__6167 (
            .O(N__34726),
            .I(N__34696));
    InMux I__6166 (
            .O(N__34725),
            .I(N__34687));
    InMux I__6165 (
            .O(N__34722),
            .I(N__34687));
    InMux I__6164 (
            .O(N__34721),
            .I(N__34687));
    InMux I__6163 (
            .O(N__34720),
            .I(N__34687));
    InMux I__6162 (
            .O(N__34717),
            .I(N__34678));
    InMux I__6161 (
            .O(N__34716),
            .I(N__34678));
    InMux I__6160 (
            .O(N__34715),
            .I(N__34678));
    InMux I__6159 (
            .O(N__34712),
            .I(N__34678));
    InMux I__6158 (
            .O(N__34709),
            .I(N__34665));
    InMux I__6157 (
            .O(N__34708),
            .I(N__34665));
    InMux I__6156 (
            .O(N__34707),
            .I(N__34665));
    InMux I__6155 (
            .O(N__34704),
            .I(N__34665));
    InMux I__6154 (
            .O(N__34703),
            .I(N__34665));
    InMux I__6153 (
            .O(N__34702),
            .I(N__34665));
    InMux I__6152 (
            .O(N__34701),
            .I(N__34660));
    CascadeMux I__6151 (
            .O(N__34700),
            .I(N__34657));
    CascadeMux I__6150 (
            .O(N__34699),
            .I(N__34652));
    LocalMux I__6149 (
            .O(N__34696),
            .I(N__34648));
    LocalMux I__6148 (
            .O(N__34687),
            .I(N__34641));
    LocalMux I__6147 (
            .O(N__34678),
            .I(N__34641));
    LocalMux I__6146 (
            .O(N__34665),
            .I(N__34641));
    InMux I__6145 (
            .O(N__34664),
            .I(N__34636));
    InMux I__6144 (
            .O(N__34663),
            .I(N__34636));
    LocalMux I__6143 (
            .O(N__34660),
            .I(N__34626));
    InMux I__6142 (
            .O(N__34657),
            .I(N__34615));
    InMux I__6141 (
            .O(N__34656),
            .I(N__34615));
    InMux I__6140 (
            .O(N__34655),
            .I(N__34615));
    InMux I__6139 (
            .O(N__34652),
            .I(N__34615));
    InMux I__6138 (
            .O(N__34651),
            .I(N__34615));
    Span4Mux_h I__6137 (
            .O(N__34648),
            .I(N__34608));
    Span4Mux_v I__6136 (
            .O(N__34641),
            .I(N__34608));
    LocalMux I__6135 (
            .O(N__34636),
            .I(N__34608));
    InMux I__6134 (
            .O(N__34635),
            .I(N__34599));
    InMux I__6133 (
            .O(N__34634),
            .I(N__34599));
    InMux I__6132 (
            .O(N__34633),
            .I(N__34599));
    InMux I__6131 (
            .O(N__34632),
            .I(N__34599));
    InMux I__6130 (
            .O(N__34631),
            .I(N__34594));
    InMux I__6129 (
            .O(N__34630),
            .I(N__34594));
    InMux I__6128 (
            .O(N__34629),
            .I(N__34591));
    Odrv4 I__6127 (
            .O(N__34626),
            .I(n3237));
    LocalMux I__6126 (
            .O(N__34615),
            .I(n3237));
    Odrv4 I__6125 (
            .O(N__34608),
            .I(n3237));
    LocalMux I__6124 (
            .O(N__34599),
            .I(n3237));
    LocalMux I__6123 (
            .O(N__34594),
            .I(n3237));
    LocalMux I__6122 (
            .O(N__34591),
            .I(n3237));
    CascadeMux I__6121 (
            .O(N__34578),
            .I(N__34575));
    InMux I__6120 (
            .O(N__34575),
            .I(N__34572));
    LocalMux I__6119 (
            .O(N__34572),
            .I(N__34569));
    Odrv4 I__6118 (
            .O(N__34569),
            .I(n13_adj_709));
    InMux I__6117 (
            .O(N__34566),
            .I(N__34562));
    InMux I__6116 (
            .O(N__34565),
            .I(N__34559));
    LocalMux I__6115 (
            .O(N__34562),
            .I(N__34556));
    LocalMux I__6114 (
            .O(N__34559),
            .I(N__34551));
    Span4Mux_v I__6113 (
            .O(N__34556),
            .I(N__34551));
    Odrv4 I__6112 (
            .O(N__34551),
            .I(n319));
    CascadeMux I__6111 (
            .O(N__34548),
            .I(n14780_cascade_));
    CascadeMux I__6110 (
            .O(N__34545),
            .I(N__34541));
    InMux I__6109 (
            .O(N__34544),
            .I(N__34538));
    InMux I__6108 (
            .O(N__34541),
            .I(N__34535));
    LocalMux I__6107 (
            .O(N__34538),
            .I(N__34531));
    LocalMux I__6106 (
            .O(N__34535),
            .I(N__34528));
    InMux I__6105 (
            .O(N__34534),
            .I(N__34525));
    Span4Mux_h I__6104 (
            .O(N__34531),
            .I(N__34522));
    Span4Mux_v I__6103 (
            .O(N__34528),
            .I(N__34517));
    LocalMux I__6102 (
            .O(N__34525),
            .I(N__34517));
    Odrv4 I__6101 (
            .O(N__34522),
            .I(n3128));
    Odrv4 I__6100 (
            .O(N__34517),
            .I(n3128));
    CascadeMux I__6099 (
            .O(N__34512),
            .I(N__34509));
    InMux I__6098 (
            .O(N__34509),
            .I(N__34506));
    LocalMux I__6097 (
            .O(N__34506),
            .I(N__34503));
    Span4Mux_h I__6096 (
            .O(N__34503),
            .I(N__34500));
    Odrv4 I__6095 (
            .O(N__34500),
            .I(n3195));
    InMux I__6094 (
            .O(N__34497),
            .I(N__34493));
    CascadeMux I__6093 (
            .O(N__34496),
            .I(N__34490));
    LocalMux I__6092 (
            .O(N__34493),
            .I(N__34487));
    InMux I__6091 (
            .O(N__34490),
            .I(N__34484));
    Span4Mux_h I__6090 (
            .O(N__34487),
            .I(N__34481));
    LocalMux I__6089 (
            .O(N__34484),
            .I(N__34478));
    Span4Mux_v I__6088 (
            .O(N__34481),
            .I(N__34475));
    Span4Mux_v I__6087 (
            .O(N__34478),
            .I(N__34472));
    Odrv4 I__6086 (
            .O(N__34475),
            .I(n3117));
    Odrv4 I__6085 (
            .O(N__34472),
            .I(n3117));
    InMux I__6084 (
            .O(N__34467),
            .I(N__34464));
    LocalMux I__6083 (
            .O(N__34464),
            .I(N__34461));
    Odrv4 I__6082 (
            .O(N__34461),
            .I(n3184));
    InMux I__6081 (
            .O(N__34458),
            .I(N__34454));
    InMux I__6080 (
            .O(N__34457),
            .I(N__34451));
    LocalMux I__6079 (
            .O(N__34454),
            .I(N__34448));
    LocalMux I__6078 (
            .O(N__34451),
            .I(N__34445));
    Span4Mux_h I__6077 (
            .O(N__34448),
            .I(N__34441));
    Span4Mux_v I__6076 (
            .O(N__34445),
            .I(N__34438));
    InMux I__6075 (
            .O(N__34444),
            .I(N__34435));
    Odrv4 I__6074 (
            .O(N__34441),
            .I(n3119));
    Odrv4 I__6073 (
            .O(N__34438),
            .I(n3119));
    LocalMux I__6072 (
            .O(N__34435),
            .I(n3119));
    CascadeMux I__6071 (
            .O(N__34428),
            .I(N__34425));
    InMux I__6070 (
            .O(N__34425),
            .I(N__34422));
    LocalMux I__6069 (
            .O(N__34422),
            .I(N__34419));
    Span4Mux_h I__6068 (
            .O(N__34419),
            .I(N__34416));
    Odrv4 I__6067 (
            .O(N__34416),
            .I(n3186));
    CascadeMux I__6066 (
            .O(N__34413),
            .I(n3218_cascade_));
    InMux I__6065 (
            .O(N__34410),
            .I(N__34407));
    LocalMux I__6064 (
            .O(N__34407),
            .I(n14778));
    InMux I__6063 (
            .O(N__34404),
            .I(N__34401));
    LocalMux I__6062 (
            .O(N__34401),
            .I(N__34398));
    Odrv4 I__6061 (
            .O(N__34398),
            .I(n12030));
    InMux I__6060 (
            .O(N__34395),
            .I(N__34392));
    LocalMux I__6059 (
            .O(N__34392),
            .I(n14786));
    InMux I__6058 (
            .O(N__34389),
            .I(N__34386));
    LocalMux I__6057 (
            .O(N__34386),
            .I(n14788));
    InMux I__6056 (
            .O(N__34383),
            .I(N__34380));
    LocalMux I__6055 (
            .O(N__34380),
            .I(N__34377));
    Odrv4 I__6054 (
            .O(N__34377),
            .I(encoder0_position_scaled_12));
    InMux I__6053 (
            .O(N__34374),
            .I(N__34371));
    LocalMux I__6052 (
            .O(N__34371),
            .I(N__34368));
    Span4Mux_h I__6051 (
            .O(N__34368),
            .I(N__34365));
    Odrv4 I__6050 (
            .O(N__34365),
            .I(n3194));
    InMux I__6049 (
            .O(N__34362),
            .I(N__34358));
    CascadeMux I__6048 (
            .O(N__34361),
            .I(N__34355));
    LocalMux I__6047 (
            .O(N__34358),
            .I(N__34352));
    InMux I__6046 (
            .O(N__34355),
            .I(N__34349));
    Span4Mux_h I__6045 (
            .O(N__34352),
            .I(N__34346));
    LocalMux I__6044 (
            .O(N__34349),
            .I(N__34343));
    Odrv4 I__6043 (
            .O(N__34346),
            .I(n3127));
    Odrv12 I__6042 (
            .O(N__34343),
            .I(n3127));
    InMux I__6041 (
            .O(N__34338),
            .I(N__34335));
    LocalMux I__6040 (
            .O(N__34335),
            .I(N__34332));
    Span4Mux_h I__6039 (
            .O(N__34332),
            .I(N__34327));
    InMux I__6038 (
            .O(N__34331),
            .I(N__34324));
    InMux I__6037 (
            .O(N__34330),
            .I(N__34321));
    Odrv4 I__6036 (
            .O(N__34327),
            .I(n3013));
    LocalMux I__6035 (
            .O(N__34324),
            .I(n3013));
    LocalMux I__6034 (
            .O(N__34321),
            .I(n3013));
    InMux I__6033 (
            .O(N__34314),
            .I(n12958));
    InMux I__6032 (
            .O(N__34311),
            .I(n12959));
    InMux I__6031 (
            .O(N__34308),
            .I(n12960));
    InMux I__6030 (
            .O(N__34305),
            .I(N__34302));
    LocalMux I__6029 (
            .O(N__34302),
            .I(N__34299));
    Span4Mux_h I__6028 (
            .O(N__34299),
            .I(N__34296));
    Odrv4 I__6027 (
            .O(N__34296),
            .I(n3177));
    InMux I__6026 (
            .O(N__34293),
            .I(N__34289));
    CascadeMux I__6025 (
            .O(N__34292),
            .I(N__34286));
    LocalMux I__6024 (
            .O(N__34289),
            .I(N__34282));
    InMux I__6023 (
            .O(N__34286),
            .I(N__34279));
    InMux I__6022 (
            .O(N__34285),
            .I(N__34276));
    Span4Mux_h I__6021 (
            .O(N__34282),
            .I(N__34273));
    LocalMux I__6020 (
            .O(N__34279),
            .I(N__34268));
    LocalMux I__6019 (
            .O(N__34276),
            .I(N__34268));
    Span4Mux_v I__6018 (
            .O(N__34273),
            .I(N__34265));
    Span4Mux_h I__6017 (
            .O(N__34268),
            .I(N__34262));
    Odrv4 I__6016 (
            .O(N__34265),
            .I(n3110));
    Odrv4 I__6015 (
            .O(N__34262),
            .I(n3110));
    CascadeMux I__6014 (
            .O(N__34257),
            .I(n31_adj_714_cascade_));
    InMux I__6013 (
            .O(N__34254),
            .I(N__34251));
    LocalMux I__6012 (
            .O(N__34251),
            .I(N__34248));
    Odrv4 I__6011 (
            .O(N__34248),
            .I(n14232));
    InMux I__6010 (
            .O(N__34245),
            .I(N__34240));
    InMux I__6009 (
            .O(N__34244),
            .I(N__34237));
    CascadeMux I__6008 (
            .O(N__34243),
            .I(N__34234));
    LocalMux I__6007 (
            .O(N__34240),
            .I(N__34231));
    LocalMux I__6006 (
            .O(N__34237),
            .I(N__34228));
    InMux I__6005 (
            .O(N__34234),
            .I(N__34225));
    Span4Mux_s3_v I__6004 (
            .O(N__34231),
            .I(N__34222));
    Odrv4 I__6003 (
            .O(N__34228),
            .I(n3126));
    LocalMux I__6002 (
            .O(N__34225),
            .I(n3126));
    Odrv4 I__6001 (
            .O(N__34222),
            .I(n3126));
    CascadeMux I__6000 (
            .O(N__34215),
            .I(N__34212));
    InMux I__5999 (
            .O(N__34212),
            .I(N__34209));
    LocalMux I__5998 (
            .O(N__34209),
            .I(N__34206));
    Odrv4 I__5997 (
            .O(N__34206),
            .I(n3193));
    CascadeMux I__5996 (
            .O(N__34203),
            .I(n3225_cascade_));
    CascadeMux I__5995 (
            .O(N__34200),
            .I(n14776_cascade_));
    InMux I__5994 (
            .O(N__34197),
            .I(N__34194));
    LocalMux I__5993 (
            .O(N__34194),
            .I(n14764));
    InMux I__5992 (
            .O(N__34191),
            .I(N__34188));
    LocalMux I__5991 (
            .O(N__34188),
            .I(N__34185));
    Span4Mux_h I__5990 (
            .O(N__34185),
            .I(N__34181));
    InMux I__5989 (
            .O(N__34184),
            .I(N__34178));
    Span4Mux_v I__5988 (
            .O(N__34181),
            .I(N__34173));
    LocalMux I__5987 (
            .O(N__34178),
            .I(N__34173));
    Odrv4 I__5986 (
            .O(N__34173),
            .I(n15714));
    InMux I__5985 (
            .O(N__34170),
            .I(N__34164));
    CascadeMux I__5984 (
            .O(N__34169),
            .I(N__34156));
    CascadeMux I__5983 (
            .O(N__34168),
            .I(N__34149));
    CascadeMux I__5982 (
            .O(N__34167),
            .I(N__34145));
    LocalMux I__5981 (
            .O(N__34164),
            .I(N__34141));
    InMux I__5980 (
            .O(N__34163),
            .I(N__34138));
    CascadeMux I__5979 (
            .O(N__34162),
            .I(N__34134));
    CascadeMux I__5978 (
            .O(N__34161),
            .I(N__34130));
    InMux I__5977 (
            .O(N__34160),
            .I(N__34122));
    InMux I__5976 (
            .O(N__34159),
            .I(N__34122));
    InMux I__5975 (
            .O(N__34156),
            .I(N__34119));
    InMux I__5974 (
            .O(N__34155),
            .I(N__34114));
    InMux I__5973 (
            .O(N__34154),
            .I(N__34114));
    InMux I__5972 (
            .O(N__34153),
            .I(N__34109));
    InMux I__5971 (
            .O(N__34152),
            .I(N__34109));
    InMux I__5970 (
            .O(N__34149),
            .I(N__34104));
    InMux I__5969 (
            .O(N__34148),
            .I(N__34104));
    InMux I__5968 (
            .O(N__34145),
            .I(N__34099));
    InMux I__5967 (
            .O(N__34144),
            .I(N__34099));
    Span4Mux_v I__5966 (
            .O(N__34141),
            .I(N__34094));
    LocalMux I__5965 (
            .O(N__34138),
            .I(N__34094));
    InMux I__5964 (
            .O(N__34137),
            .I(N__34081));
    InMux I__5963 (
            .O(N__34134),
            .I(N__34081));
    InMux I__5962 (
            .O(N__34133),
            .I(N__34081));
    InMux I__5961 (
            .O(N__34130),
            .I(N__34081));
    InMux I__5960 (
            .O(N__34129),
            .I(N__34081));
    InMux I__5959 (
            .O(N__34128),
            .I(N__34081));
    InMux I__5958 (
            .O(N__34127),
            .I(N__34078));
    LocalMux I__5957 (
            .O(N__34122),
            .I(N__34075));
    LocalMux I__5956 (
            .O(N__34119),
            .I(N__34070));
    LocalMux I__5955 (
            .O(N__34114),
            .I(N__34070));
    LocalMux I__5954 (
            .O(N__34109),
            .I(n2148));
    LocalMux I__5953 (
            .O(N__34104),
            .I(n2148));
    LocalMux I__5952 (
            .O(N__34099),
            .I(n2148));
    Odrv4 I__5951 (
            .O(N__34094),
            .I(n2148));
    LocalMux I__5950 (
            .O(N__34081),
            .I(n2148));
    LocalMux I__5949 (
            .O(N__34078),
            .I(n2148));
    Odrv4 I__5948 (
            .O(N__34075),
            .I(n2148));
    Odrv4 I__5947 (
            .O(N__34070),
            .I(n2148));
    InMux I__5946 (
            .O(N__34053),
            .I(n12949));
    InMux I__5945 (
            .O(N__34050),
            .I(N__34047));
    LocalMux I__5944 (
            .O(N__34047),
            .I(N__34043));
    CascadeMux I__5943 (
            .O(N__34046),
            .I(N__34040));
    Span4Mux_v I__5942 (
            .O(N__34043),
            .I(N__34037));
    InMux I__5941 (
            .O(N__34040),
            .I(N__34034));
    Odrv4 I__5940 (
            .O(N__34037),
            .I(n15689));
    LocalMux I__5939 (
            .O(N__34034),
            .I(n15689));
    InMux I__5938 (
            .O(N__34029),
            .I(N__34021));
    CascadeMux I__5937 (
            .O(N__34028),
            .I(N__34012));
    CascadeMux I__5936 (
            .O(N__34027),
            .I(N__34007));
    CascadeMux I__5935 (
            .O(N__34026),
            .I(N__34004));
    InMux I__5934 (
            .O(N__34025),
            .I(N__33997));
    InMux I__5933 (
            .O(N__34024),
            .I(N__33997));
    LocalMux I__5932 (
            .O(N__34021),
            .I(N__33994));
    InMux I__5931 (
            .O(N__34020),
            .I(N__33989));
    InMux I__5930 (
            .O(N__34019),
            .I(N__33989));
    InMux I__5929 (
            .O(N__34018),
            .I(N__33986));
    CascadeMux I__5928 (
            .O(N__34017),
            .I(N__33981));
    CascadeMux I__5927 (
            .O(N__34016),
            .I(N__33978));
    InMux I__5926 (
            .O(N__34015),
            .I(N__33974));
    InMux I__5925 (
            .O(N__34012),
            .I(N__33967));
    InMux I__5924 (
            .O(N__34011),
            .I(N__33967));
    InMux I__5923 (
            .O(N__34010),
            .I(N__33967));
    InMux I__5922 (
            .O(N__34007),
            .I(N__33958));
    InMux I__5921 (
            .O(N__34004),
            .I(N__33958));
    InMux I__5920 (
            .O(N__34003),
            .I(N__33958));
    InMux I__5919 (
            .O(N__34002),
            .I(N__33958));
    LocalMux I__5918 (
            .O(N__33997),
            .I(N__33955));
    Span4Mux_v I__5917 (
            .O(N__33994),
            .I(N__33948));
    LocalMux I__5916 (
            .O(N__33989),
            .I(N__33948));
    LocalMux I__5915 (
            .O(N__33986),
            .I(N__33948));
    InMux I__5914 (
            .O(N__33985),
            .I(N__33943));
    InMux I__5913 (
            .O(N__33984),
            .I(N__33943));
    InMux I__5912 (
            .O(N__33981),
            .I(N__33936));
    InMux I__5911 (
            .O(N__33978),
            .I(N__33936));
    InMux I__5910 (
            .O(N__33977),
            .I(N__33936));
    LocalMux I__5909 (
            .O(N__33974),
            .I(n2049));
    LocalMux I__5908 (
            .O(N__33967),
            .I(n2049));
    LocalMux I__5907 (
            .O(N__33958),
            .I(n2049));
    Odrv4 I__5906 (
            .O(N__33955),
            .I(n2049));
    Odrv4 I__5905 (
            .O(N__33948),
            .I(n2049));
    LocalMux I__5904 (
            .O(N__33943),
            .I(n2049));
    LocalMux I__5903 (
            .O(N__33936),
            .I(n2049));
    InMux I__5902 (
            .O(N__33921),
            .I(n12950));
    InMux I__5901 (
            .O(N__33918),
            .I(n12951));
    InMux I__5900 (
            .O(N__33915),
            .I(n12952));
    InMux I__5899 (
            .O(N__33912),
            .I(bfn_7_25_0_));
    InMux I__5898 (
            .O(N__33909),
            .I(n12954));
    InMux I__5897 (
            .O(N__33906),
            .I(n12955));
    InMux I__5896 (
            .O(N__33903),
            .I(n12956));
    InMux I__5895 (
            .O(N__33900),
            .I(n12957));
    InMux I__5894 (
            .O(N__33897),
            .I(N__33888));
    InMux I__5893 (
            .O(N__33896),
            .I(N__33881));
    InMux I__5892 (
            .O(N__33895),
            .I(N__33881));
    InMux I__5891 (
            .O(N__33894),
            .I(N__33874));
    InMux I__5890 (
            .O(N__33893),
            .I(N__33874));
    InMux I__5889 (
            .O(N__33892),
            .I(N__33874));
    CascadeMux I__5888 (
            .O(N__33891),
            .I(N__33868));
    LocalMux I__5887 (
            .O(N__33888),
            .I(N__33859));
    CascadeMux I__5886 (
            .O(N__33887),
            .I(N__33855));
    InMux I__5885 (
            .O(N__33886),
            .I(N__33851));
    LocalMux I__5884 (
            .O(N__33881),
            .I(N__33846));
    LocalMux I__5883 (
            .O(N__33874),
            .I(N__33841));
    InMux I__5882 (
            .O(N__33873),
            .I(N__33830));
    InMux I__5881 (
            .O(N__33872),
            .I(N__33830));
    InMux I__5880 (
            .O(N__33871),
            .I(N__33830));
    InMux I__5879 (
            .O(N__33868),
            .I(N__33830));
    InMux I__5878 (
            .O(N__33867),
            .I(N__33830));
    InMux I__5877 (
            .O(N__33866),
            .I(N__33825));
    InMux I__5876 (
            .O(N__33865),
            .I(N__33825));
    InMux I__5875 (
            .O(N__33864),
            .I(N__33818));
    InMux I__5874 (
            .O(N__33863),
            .I(N__33818));
    InMux I__5873 (
            .O(N__33862),
            .I(N__33818));
    Span4Mux_v I__5872 (
            .O(N__33859),
            .I(N__33815));
    InMux I__5871 (
            .O(N__33858),
            .I(N__33808));
    InMux I__5870 (
            .O(N__33855),
            .I(N__33808));
    InMux I__5869 (
            .O(N__33854),
            .I(N__33808));
    LocalMux I__5868 (
            .O(N__33851),
            .I(N__33805));
    CascadeMux I__5867 (
            .O(N__33850),
            .I(N__33800));
    CascadeMux I__5866 (
            .O(N__33849),
            .I(N__33797));
    Span4Mux_v I__5865 (
            .O(N__33846),
            .I(N__33792));
    InMux I__5864 (
            .O(N__33845),
            .I(N__33789));
    InMux I__5863 (
            .O(N__33844),
            .I(N__33786));
    Span4Mux_s1_v I__5862 (
            .O(N__33841),
            .I(N__33777));
    LocalMux I__5861 (
            .O(N__33830),
            .I(N__33777));
    LocalMux I__5860 (
            .O(N__33825),
            .I(N__33777));
    LocalMux I__5859 (
            .O(N__33818),
            .I(N__33777));
    Span4Mux_h I__5858 (
            .O(N__33815),
            .I(N__33770));
    LocalMux I__5857 (
            .O(N__33808),
            .I(N__33770));
    Span4Mux_s3_h I__5856 (
            .O(N__33805),
            .I(N__33770));
    InMux I__5855 (
            .O(N__33804),
            .I(N__33759));
    InMux I__5854 (
            .O(N__33803),
            .I(N__33759));
    InMux I__5853 (
            .O(N__33800),
            .I(N__33759));
    InMux I__5852 (
            .O(N__33797),
            .I(N__33759));
    InMux I__5851 (
            .O(N__33796),
            .I(N__33759));
    InMux I__5850 (
            .O(N__33795),
            .I(N__33756));
    Odrv4 I__5849 (
            .O(N__33792),
            .I(n2940));
    LocalMux I__5848 (
            .O(N__33789),
            .I(n2940));
    LocalMux I__5847 (
            .O(N__33786),
            .I(n2940));
    Odrv4 I__5846 (
            .O(N__33777),
            .I(n2940));
    Odrv4 I__5845 (
            .O(N__33770),
            .I(n2940));
    LocalMux I__5844 (
            .O(N__33759),
            .I(n2940));
    LocalMux I__5843 (
            .O(N__33756),
            .I(n2940));
    InMux I__5842 (
            .O(N__33741),
            .I(n12941));
    InMux I__5841 (
            .O(N__33738),
            .I(N__33735));
    LocalMux I__5840 (
            .O(N__33735),
            .I(N__33732));
    Span4Mux_v I__5839 (
            .O(N__33732),
            .I(N__33728));
    CascadeMux I__5838 (
            .O(N__33731),
            .I(N__33725));
    Span4Mux_h I__5837 (
            .O(N__33728),
            .I(N__33722));
    InMux I__5836 (
            .O(N__33725),
            .I(N__33719));
    Odrv4 I__5835 (
            .O(N__33722),
            .I(n15346));
    LocalMux I__5834 (
            .O(N__33719),
            .I(n15346));
    InMux I__5833 (
            .O(N__33714),
            .I(N__33710));
    InMux I__5832 (
            .O(N__33713),
            .I(N__33702));
    LocalMux I__5831 (
            .O(N__33710),
            .I(N__33693));
    InMux I__5830 (
            .O(N__33709),
            .I(N__33690));
    InMux I__5829 (
            .O(N__33708),
            .I(N__33683));
    InMux I__5828 (
            .O(N__33707),
            .I(N__33683));
    InMux I__5827 (
            .O(N__33706),
            .I(N__33683));
    InMux I__5826 (
            .O(N__33705),
            .I(N__33680));
    LocalMux I__5825 (
            .O(N__33702),
            .I(N__33677));
    CascadeMux I__5824 (
            .O(N__33701),
            .I(N__33673));
    CascadeMux I__5823 (
            .O(N__33700),
            .I(N__33670));
    CascadeMux I__5822 (
            .O(N__33699),
            .I(N__33664));
    CascadeMux I__5821 (
            .O(N__33698),
            .I(N__33658));
    CascadeMux I__5820 (
            .O(N__33697),
            .I(N__33652));
    InMux I__5819 (
            .O(N__33696),
            .I(N__33648));
    Span4Mux_v I__5818 (
            .O(N__33693),
            .I(N__33642));
    LocalMux I__5817 (
            .O(N__33690),
            .I(N__33639));
    LocalMux I__5816 (
            .O(N__33683),
            .I(N__33636));
    LocalMux I__5815 (
            .O(N__33680),
            .I(N__33633));
    Span4Mux_s2_h I__5814 (
            .O(N__33677),
            .I(N__33630));
    InMux I__5813 (
            .O(N__33676),
            .I(N__33627));
    InMux I__5812 (
            .O(N__33673),
            .I(N__33616));
    InMux I__5811 (
            .O(N__33670),
            .I(N__33616));
    InMux I__5810 (
            .O(N__33669),
            .I(N__33616));
    InMux I__5809 (
            .O(N__33668),
            .I(N__33616));
    InMux I__5808 (
            .O(N__33667),
            .I(N__33616));
    InMux I__5807 (
            .O(N__33664),
            .I(N__33607));
    InMux I__5806 (
            .O(N__33663),
            .I(N__33607));
    InMux I__5805 (
            .O(N__33662),
            .I(N__33607));
    InMux I__5804 (
            .O(N__33661),
            .I(N__33607));
    InMux I__5803 (
            .O(N__33658),
            .I(N__33594));
    InMux I__5802 (
            .O(N__33657),
            .I(N__33594));
    InMux I__5801 (
            .O(N__33656),
            .I(N__33594));
    InMux I__5800 (
            .O(N__33655),
            .I(N__33594));
    InMux I__5799 (
            .O(N__33652),
            .I(N__33594));
    InMux I__5798 (
            .O(N__33651),
            .I(N__33594));
    LocalMux I__5797 (
            .O(N__33648),
            .I(N__33591));
    InMux I__5796 (
            .O(N__33647),
            .I(N__33588));
    InMux I__5795 (
            .O(N__33646),
            .I(N__33583));
    InMux I__5794 (
            .O(N__33645),
            .I(N__33583));
    Span4Mux_h I__5793 (
            .O(N__33642),
            .I(N__33574));
    Span4Mux_v I__5792 (
            .O(N__33639),
            .I(N__33574));
    Span4Mux_s3_h I__5791 (
            .O(N__33636),
            .I(N__33574));
    Span4Mux_s2_v I__5790 (
            .O(N__33633),
            .I(N__33574));
    Odrv4 I__5789 (
            .O(N__33630),
            .I(n2841));
    LocalMux I__5788 (
            .O(N__33627),
            .I(n2841));
    LocalMux I__5787 (
            .O(N__33616),
            .I(n2841));
    LocalMux I__5786 (
            .O(N__33607),
            .I(n2841));
    LocalMux I__5785 (
            .O(N__33594),
            .I(n2841));
    Odrv12 I__5784 (
            .O(N__33591),
            .I(n2841));
    LocalMux I__5783 (
            .O(N__33588),
            .I(n2841));
    LocalMux I__5782 (
            .O(N__33583),
            .I(n2841));
    Odrv4 I__5781 (
            .O(N__33574),
            .I(n2841));
    InMux I__5780 (
            .O(N__33555),
            .I(n12942));
    InMux I__5779 (
            .O(N__33552),
            .I(N__33548));
    CascadeMux I__5778 (
            .O(N__33551),
            .I(N__33545));
    LocalMux I__5777 (
            .O(N__33548),
            .I(N__33542));
    InMux I__5776 (
            .O(N__33545),
            .I(N__33539));
    Span4Mux_v I__5775 (
            .O(N__33542),
            .I(N__33536));
    LocalMux I__5774 (
            .O(N__33539),
            .I(N__33533));
    Odrv4 I__5773 (
            .O(N__33536),
            .I(n15310));
    Odrv4 I__5772 (
            .O(N__33533),
            .I(n15310));
    InMux I__5771 (
            .O(N__33528),
            .I(N__33525));
    LocalMux I__5770 (
            .O(N__33525),
            .I(N__33518));
    InMux I__5769 (
            .O(N__33524),
            .I(N__33507));
    CascadeMux I__5768 (
            .O(N__33523),
            .I(N__33499));
    CascadeMux I__5767 (
            .O(N__33522),
            .I(N__33496));
    CascadeMux I__5766 (
            .O(N__33521),
            .I(N__33493));
    Span4Mux_h I__5765 (
            .O(N__33518),
            .I(N__33488));
    InMux I__5764 (
            .O(N__33517),
            .I(N__33483));
    InMux I__5763 (
            .O(N__33516),
            .I(N__33483));
    CascadeMux I__5762 (
            .O(N__33515),
            .I(N__33480));
    CascadeMux I__5761 (
            .O(N__33514),
            .I(N__33477));
    CascadeMux I__5760 (
            .O(N__33513),
            .I(N__33474));
    CascadeMux I__5759 (
            .O(N__33512),
            .I(N__33471));
    InMux I__5758 (
            .O(N__33511),
            .I(N__33465));
    InMux I__5757 (
            .O(N__33510),
            .I(N__33465));
    LocalMux I__5756 (
            .O(N__33507),
            .I(N__33460));
    CascadeMux I__5755 (
            .O(N__33506),
            .I(N__33457));
    CascadeMux I__5754 (
            .O(N__33505),
            .I(N__33453));
    CascadeMux I__5753 (
            .O(N__33504),
            .I(N__33449));
    CascadeMux I__5752 (
            .O(N__33503),
            .I(N__33446));
    InMux I__5751 (
            .O(N__33502),
            .I(N__33432));
    InMux I__5750 (
            .O(N__33499),
            .I(N__33432));
    InMux I__5749 (
            .O(N__33496),
            .I(N__33432));
    InMux I__5748 (
            .O(N__33493),
            .I(N__33432));
    InMux I__5747 (
            .O(N__33492),
            .I(N__33432));
    InMux I__5746 (
            .O(N__33491),
            .I(N__33432));
    Span4Mux_h I__5745 (
            .O(N__33488),
            .I(N__33427));
    LocalMux I__5744 (
            .O(N__33483),
            .I(N__33427));
    InMux I__5743 (
            .O(N__33480),
            .I(N__33416));
    InMux I__5742 (
            .O(N__33477),
            .I(N__33416));
    InMux I__5741 (
            .O(N__33474),
            .I(N__33416));
    InMux I__5740 (
            .O(N__33471),
            .I(N__33416));
    InMux I__5739 (
            .O(N__33470),
            .I(N__33416));
    LocalMux I__5738 (
            .O(N__33465),
            .I(N__33413));
    InMux I__5737 (
            .O(N__33464),
            .I(N__33408));
    InMux I__5736 (
            .O(N__33463),
            .I(N__33408));
    Span4Mux_s3_v I__5735 (
            .O(N__33460),
            .I(N__33405));
    InMux I__5734 (
            .O(N__33457),
            .I(N__33400));
    InMux I__5733 (
            .O(N__33456),
            .I(N__33400));
    InMux I__5732 (
            .O(N__33453),
            .I(N__33389));
    InMux I__5731 (
            .O(N__33452),
            .I(N__33389));
    InMux I__5730 (
            .O(N__33449),
            .I(N__33389));
    InMux I__5729 (
            .O(N__33446),
            .I(N__33389));
    InMux I__5728 (
            .O(N__33445),
            .I(N__33389));
    LocalMux I__5727 (
            .O(N__33432),
            .I(n2742));
    Odrv4 I__5726 (
            .O(N__33427),
            .I(n2742));
    LocalMux I__5725 (
            .O(N__33416),
            .I(n2742));
    Odrv4 I__5724 (
            .O(N__33413),
            .I(n2742));
    LocalMux I__5723 (
            .O(N__33408),
            .I(n2742));
    Odrv4 I__5722 (
            .O(N__33405),
            .I(n2742));
    LocalMux I__5721 (
            .O(N__33400),
            .I(n2742));
    LocalMux I__5720 (
            .O(N__33389),
            .I(n2742));
    InMux I__5719 (
            .O(N__33372),
            .I(n12943));
    InMux I__5718 (
            .O(N__33369),
            .I(N__33366));
    LocalMux I__5717 (
            .O(N__33366),
            .I(N__33363));
    Span4Mux_h I__5716 (
            .O(N__33363),
            .I(N__33359));
    InMux I__5715 (
            .O(N__33362),
            .I(N__33356));
    Odrv4 I__5714 (
            .O(N__33359),
            .I(n15852));
    LocalMux I__5713 (
            .O(N__33356),
            .I(n15852));
    CascadeMux I__5712 (
            .O(N__33351),
            .I(N__33346));
    InMux I__5711 (
            .O(N__33350),
            .I(N__33336));
    InMux I__5710 (
            .O(N__33349),
            .I(N__33331));
    InMux I__5709 (
            .O(N__33346),
            .I(N__33325));
    CascadeMux I__5708 (
            .O(N__33345),
            .I(N__33322));
    InMux I__5707 (
            .O(N__33344),
            .I(N__33318));
    InMux I__5706 (
            .O(N__33343),
            .I(N__33315));
    CascadeMux I__5705 (
            .O(N__33342),
            .I(N__33311));
    CascadeMux I__5704 (
            .O(N__33341),
            .I(N__33307));
    CascadeMux I__5703 (
            .O(N__33340),
            .I(N__33304));
    CascadeMux I__5702 (
            .O(N__33339),
            .I(N__33298));
    LocalMux I__5701 (
            .O(N__33336),
            .I(N__33293));
    InMux I__5700 (
            .O(N__33335),
            .I(N__33288));
    InMux I__5699 (
            .O(N__33334),
            .I(N__33288));
    LocalMux I__5698 (
            .O(N__33331),
            .I(N__33285));
    InMux I__5697 (
            .O(N__33330),
            .I(N__33282));
    CascadeMux I__5696 (
            .O(N__33329),
            .I(N__33279));
    CascadeMux I__5695 (
            .O(N__33328),
            .I(N__33275));
    LocalMux I__5694 (
            .O(N__33325),
            .I(N__33270));
    InMux I__5693 (
            .O(N__33322),
            .I(N__33265));
    InMux I__5692 (
            .O(N__33321),
            .I(N__33265));
    LocalMux I__5691 (
            .O(N__33318),
            .I(N__33260));
    LocalMux I__5690 (
            .O(N__33315),
            .I(N__33260));
    InMux I__5689 (
            .O(N__33314),
            .I(N__33253));
    InMux I__5688 (
            .O(N__33311),
            .I(N__33253));
    InMux I__5687 (
            .O(N__33310),
            .I(N__33253));
    InMux I__5686 (
            .O(N__33307),
            .I(N__33244));
    InMux I__5685 (
            .O(N__33304),
            .I(N__33244));
    InMux I__5684 (
            .O(N__33303),
            .I(N__33244));
    InMux I__5683 (
            .O(N__33302),
            .I(N__33244));
    InMux I__5682 (
            .O(N__33301),
            .I(N__33235));
    InMux I__5681 (
            .O(N__33298),
            .I(N__33235));
    InMux I__5680 (
            .O(N__33297),
            .I(N__33235));
    InMux I__5679 (
            .O(N__33296),
            .I(N__33235));
    Span4Mux_h I__5678 (
            .O(N__33293),
            .I(N__33226));
    LocalMux I__5677 (
            .O(N__33288),
            .I(N__33226));
    Span4Mux_s3_h I__5676 (
            .O(N__33285),
            .I(N__33226));
    LocalMux I__5675 (
            .O(N__33282),
            .I(N__33226));
    InMux I__5674 (
            .O(N__33279),
            .I(N__33215));
    InMux I__5673 (
            .O(N__33278),
            .I(N__33215));
    InMux I__5672 (
            .O(N__33275),
            .I(N__33215));
    InMux I__5671 (
            .O(N__33274),
            .I(N__33215));
    InMux I__5670 (
            .O(N__33273),
            .I(N__33215));
    Odrv4 I__5669 (
            .O(N__33270),
            .I(n2643));
    LocalMux I__5668 (
            .O(N__33265),
            .I(n2643));
    Odrv4 I__5667 (
            .O(N__33260),
            .I(n2643));
    LocalMux I__5666 (
            .O(N__33253),
            .I(n2643));
    LocalMux I__5665 (
            .O(N__33244),
            .I(n2643));
    LocalMux I__5664 (
            .O(N__33235),
            .I(n2643));
    Odrv4 I__5663 (
            .O(N__33226),
            .I(n2643));
    LocalMux I__5662 (
            .O(N__33215),
            .I(n2643));
    InMux I__5661 (
            .O(N__33198),
            .I(n12944));
    InMux I__5660 (
            .O(N__33195),
            .I(N__33192));
    LocalMux I__5659 (
            .O(N__33192),
            .I(N__33189));
    Span4Mux_h I__5658 (
            .O(N__33189),
            .I(N__33185));
    CascadeMux I__5657 (
            .O(N__33188),
            .I(N__33182));
    Span4Mux_h I__5656 (
            .O(N__33185),
            .I(N__33179));
    InMux I__5655 (
            .O(N__33182),
            .I(N__33176));
    Odrv4 I__5654 (
            .O(N__33179),
            .I(n15821));
    LocalMux I__5653 (
            .O(N__33176),
            .I(n15821));
    InMux I__5652 (
            .O(N__33171),
            .I(N__33167));
    InMux I__5651 (
            .O(N__33170),
            .I(N__33160));
    LocalMux I__5650 (
            .O(N__33167),
            .I(N__33152));
    InMux I__5649 (
            .O(N__33166),
            .I(N__33149));
    CascadeMux I__5648 (
            .O(N__33165),
            .I(N__33145));
    InMux I__5647 (
            .O(N__33164),
            .I(N__33140));
    InMux I__5646 (
            .O(N__33163),
            .I(N__33140));
    LocalMux I__5645 (
            .O(N__33160),
            .I(N__33137));
    CascadeMux I__5644 (
            .O(N__33159),
            .I(N__33132));
    CascadeMux I__5643 (
            .O(N__33158),
            .I(N__33128));
    CascadeMux I__5642 (
            .O(N__33157),
            .I(N__33122));
    CascadeMux I__5641 (
            .O(N__33156),
            .I(N__33115));
    CascadeMux I__5640 (
            .O(N__33155),
            .I(N__33111));
    Span4Mux_h I__5639 (
            .O(N__33152),
            .I(N__33105));
    LocalMux I__5638 (
            .O(N__33149),
            .I(N__33105));
    InMux I__5637 (
            .O(N__33148),
            .I(N__33102));
    InMux I__5636 (
            .O(N__33145),
            .I(N__33099));
    LocalMux I__5635 (
            .O(N__33140),
            .I(N__33096));
    Span4Mux_s2_h I__5634 (
            .O(N__33137),
            .I(N__33092));
    InMux I__5633 (
            .O(N__33136),
            .I(N__33083));
    InMux I__5632 (
            .O(N__33135),
            .I(N__33083));
    InMux I__5631 (
            .O(N__33132),
            .I(N__33083));
    InMux I__5630 (
            .O(N__33131),
            .I(N__33083));
    InMux I__5629 (
            .O(N__33128),
            .I(N__33070));
    InMux I__5628 (
            .O(N__33127),
            .I(N__33070));
    InMux I__5627 (
            .O(N__33126),
            .I(N__33070));
    InMux I__5626 (
            .O(N__33125),
            .I(N__33070));
    InMux I__5625 (
            .O(N__33122),
            .I(N__33070));
    InMux I__5624 (
            .O(N__33121),
            .I(N__33070));
    InMux I__5623 (
            .O(N__33120),
            .I(N__33065));
    InMux I__5622 (
            .O(N__33119),
            .I(N__33065));
    InMux I__5621 (
            .O(N__33118),
            .I(N__33054));
    InMux I__5620 (
            .O(N__33115),
            .I(N__33054));
    InMux I__5619 (
            .O(N__33114),
            .I(N__33054));
    InMux I__5618 (
            .O(N__33111),
            .I(N__33054));
    InMux I__5617 (
            .O(N__33110),
            .I(N__33054));
    Span4Mux_h I__5616 (
            .O(N__33105),
            .I(N__33045));
    LocalMux I__5615 (
            .O(N__33102),
            .I(N__33045));
    LocalMux I__5614 (
            .O(N__33099),
            .I(N__33045));
    Span4Mux_h I__5613 (
            .O(N__33096),
            .I(N__33045));
    InMux I__5612 (
            .O(N__33095),
            .I(N__33042));
    Odrv4 I__5611 (
            .O(N__33092),
            .I(n2544));
    LocalMux I__5610 (
            .O(N__33083),
            .I(n2544));
    LocalMux I__5609 (
            .O(N__33070),
            .I(n2544));
    LocalMux I__5608 (
            .O(N__33065),
            .I(n2544));
    LocalMux I__5607 (
            .O(N__33054),
            .I(n2544));
    Odrv4 I__5606 (
            .O(N__33045),
            .I(n2544));
    LocalMux I__5605 (
            .O(N__33042),
            .I(n2544));
    InMux I__5604 (
            .O(N__33027),
            .I(bfn_7_24_0_));
    InMux I__5603 (
            .O(N__33024),
            .I(N__33021));
    LocalMux I__5602 (
            .O(N__33021),
            .I(N__33017));
    InMux I__5601 (
            .O(N__33020),
            .I(N__33014));
    Span4Mux_v I__5600 (
            .O(N__33017),
            .I(N__33011));
    LocalMux I__5599 (
            .O(N__33014),
            .I(N__33008));
    Span4Mux_h I__5598 (
            .O(N__33011),
            .I(N__33005));
    Odrv4 I__5597 (
            .O(N__33008),
            .I(n15791));
    Odrv4 I__5596 (
            .O(N__33005),
            .I(n15791));
    InMux I__5595 (
            .O(N__33000),
            .I(N__32994));
    InMux I__5594 (
            .O(N__32999),
            .I(N__32991));
    CascadeMux I__5593 (
            .O(N__32998),
            .I(N__32988));
    InMux I__5592 (
            .O(N__32997),
            .I(N__32981));
    LocalMux I__5591 (
            .O(N__32994),
            .I(N__32978));
    LocalMux I__5590 (
            .O(N__32991),
            .I(N__32973));
    InMux I__5589 (
            .O(N__32988),
            .I(N__32970));
    InMux I__5588 (
            .O(N__32987),
            .I(N__32967));
    CascadeMux I__5587 (
            .O(N__32986),
            .I(N__32962));
    CascadeMux I__5586 (
            .O(N__32985),
            .I(N__32959));
    CascadeMux I__5585 (
            .O(N__32984),
            .I(N__32955));
    LocalMux I__5584 (
            .O(N__32981),
            .I(N__32947));
    Span4Mux_s2_h I__5583 (
            .O(N__32978),
            .I(N__32947));
    CascadeMux I__5582 (
            .O(N__32977),
            .I(N__32942));
    CascadeMux I__5581 (
            .O(N__32976),
            .I(N__32937));
    Span4Mux_h I__5580 (
            .O(N__32973),
            .I(N__32930));
    LocalMux I__5579 (
            .O(N__32970),
            .I(N__32930));
    LocalMux I__5578 (
            .O(N__32967),
            .I(N__32930));
    InMux I__5577 (
            .O(N__32966),
            .I(N__32927));
    InMux I__5576 (
            .O(N__32965),
            .I(N__32914));
    InMux I__5575 (
            .O(N__32962),
            .I(N__32914));
    InMux I__5574 (
            .O(N__32959),
            .I(N__32914));
    InMux I__5573 (
            .O(N__32958),
            .I(N__32914));
    InMux I__5572 (
            .O(N__32955),
            .I(N__32914));
    InMux I__5571 (
            .O(N__32954),
            .I(N__32914));
    CascadeMux I__5570 (
            .O(N__32953),
            .I(N__32911));
    CascadeMux I__5569 (
            .O(N__32952),
            .I(N__32908));
    Span4Mux_v I__5568 (
            .O(N__32947),
            .I(N__32901));
    InMux I__5567 (
            .O(N__32946),
            .I(N__32898));
    InMux I__5566 (
            .O(N__32945),
            .I(N__32887));
    InMux I__5565 (
            .O(N__32942),
            .I(N__32887));
    InMux I__5564 (
            .O(N__32941),
            .I(N__32887));
    InMux I__5563 (
            .O(N__32940),
            .I(N__32887));
    InMux I__5562 (
            .O(N__32937),
            .I(N__32887));
    Span4Mux_v I__5561 (
            .O(N__32930),
            .I(N__32882));
    LocalMux I__5560 (
            .O(N__32927),
            .I(N__32882));
    LocalMux I__5559 (
            .O(N__32914),
            .I(N__32879));
    InMux I__5558 (
            .O(N__32911),
            .I(N__32866));
    InMux I__5557 (
            .O(N__32908),
            .I(N__32866));
    InMux I__5556 (
            .O(N__32907),
            .I(N__32866));
    InMux I__5555 (
            .O(N__32906),
            .I(N__32866));
    InMux I__5554 (
            .O(N__32905),
            .I(N__32866));
    InMux I__5553 (
            .O(N__32904),
            .I(N__32866));
    Odrv4 I__5552 (
            .O(N__32901),
            .I(n2445));
    LocalMux I__5551 (
            .O(N__32898),
            .I(n2445));
    LocalMux I__5550 (
            .O(N__32887),
            .I(n2445));
    Odrv4 I__5549 (
            .O(N__32882),
            .I(n2445));
    Odrv4 I__5548 (
            .O(N__32879),
            .I(n2445));
    LocalMux I__5547 (
            .O(N__32866),
            .I(n2445));
    InMux I__5546 (
            .O(N__32853),
            .I(n12946));
    InMux I__5545 (
            .O(N__32850),
            .I(N__32847));
    LocalMux I__5544 (
            .O(N__32847),
            .I(N__32843));
    CascadeMux I__5543 (
            .O(N__32846),
            .I(N__32840));
    Span4Mux_v I__5542 (
            .O(N__32843),
            .I(N__32837));
    InMux I__5541 (
            .O(N__32840),
            .I(N__32834));
    Odrv4 I__5540 (
            .O(N__32837),
            .I(n15765));
    LocalMux I__5539 (
            .O(N__32834),
            .I(n15765));
    InMux I__5538 (
            .O(N__32829),
            .I(N__32825));
    CascadeMux I__5537 (
            .O(N__32828),
            .I(N__32814));
    LocalMux I__5536 (
            .O(N__32825),
            .I(N__32809));
    CascadeMux I__5535 (
            .O(N__32824),
            .I(N__32802));
    CascadeMux I__5534 (
            .O(N__32823),
            .I(N__32799));
    CascadeMux I__5533 (
            .O(N__32822),
            .I(N__32795));
    CascadeMux I__5532 (
            .O(N__32821),
            .I(N__32789));
    CascadeMux I__5531 (
            .O(N__32820),
            .I(N__32786));
    CascadeMux I__5530 (
            .O(N__32819),
            .I(N__32783));
    InMux I__5529 (
            .O(N__32818),
            .I(N__32779));
    InMux I__5528 (
            .O(N__32817),
            .I(N__32772));
    InMux I__5527 (
            .O(N__32814),
            .I(N__32772));
    InMux I__5526 (
            .O(N__32813),
            .I(N__32772));
    CascadeMux I__5525 (
            .O(N__32812),
            .I(N__32769));
    Span12Mux_h I__5524 (
            .O(N__32809),
            .I(N__32765));
    InMux I__5523 (
            .O(N__32808),
            .I(N__32762));
    InMux I__5522 (
            .O(N__32807),
            .I(N__32753));
    InMux I__5521 (
            .O(N__32806),
            .I(N__32753));
    InMux I__5520 (
            .O(N__32805),
            .I(N__32753));
    InMux I__5519 (
            .O(N__32802),
            .I(N__32753));
    InMux I__5518 (
            .O(N__32799),
            .I(N__32742));
    InMux I__5517 (
            .O(N__32798),
            .I(N__32742));
    InMux I__5516 (
            .O(N__32795),
            .I(N__32742));
    InMux I__5515 (
            .O(N__32794),
            .I(N__32742));
    InMux I__5514 (
            .O(N__32793),
            .I(N__32742));
    InMux I__5513 (
            .O(N__32792),
            .I(N__32731));
    InMux I__5512 (
            .O(N__32789),
            .I(N__32731));
    InMux I__5511 (
            .O(N__32786),
            .I(N__32731));
    InMux I__5510 (
            .O(N__32783),
            .I(N__32731));
    InMux I__5509 (
            .O(N__32782),
            .I(N__32731));
    LocalMux I__5508 (
            .O(N__32779),
            .I(N__32726));
    LocalMux I__5507 (
            .O(N__32772),
            .I(N__32726));
    InMux I__5506 (
            .O(N__32769),
            .I(N__32721));
    InMux I__5505 (
            .O(N__32768),
            .I(N__32721));
    Odrv12 I__5504 (
            .O(N__32765),
            .I(n2346));
    LocalMux I__5503 (
            .O(N__32762),
            .I(n2346));
    LocalMux I__5502 (
            .O(N__32753),
            .I(n2346));
    LocalMux I__5501 (
            .O(N__32742),
            .I(n2346));
    LocalMux I__5500 (
            .O(N__32731),
            .I(n2346));
    Odrv4 I__5499 (
            .O(N__32726),
            .I(n2346));
    LocalMux I__5498 (
            .O(N__32721),
            .I(n2346));
    InMux I__5497 (
            .O(N__32706),
            .I(n12947));
    InMux I__5496 (
            .O(N__32703),
            .I(N__32699));
    CascadeMux I__5495 (
            .O(N__32702),
            .I(N__32696));
    LocalMux I__5494 (
            .O(N__32699),
            .I(N__32693));
    InMux I__5493 (
            .O(N__32696),
            .I(N__32690));
    Odrv4 I__5492 (
            .O(N__32693),
            .I(n15739));
    LocalMux I__5491 (
            .O(N__32690),
            .I(n15739));
    CascadeMux I__5490 (
            .O(N__32685),
            .I(N__32677));
    CascadeMux I__5489 (
            .O(N__32684),
            .I(N__32673));
    InMux I__5488 (
            .O(N__32683),
            .I(N__32668));
    CascadeMux I__5487 (
            .O(N__32682),
            .I(N__32665));
    CascadeMux I__5486 (
            .O(N__32681),
            .I(N__32661));
    CascadeMux I__5485 (
            .O(N__32680),
            .I(N__32657));
    InMux I__5484 (
            .O(N__32677),
            .I(N__32647));
    InMux I__5483 (
            .O(N__32676),
            .I(N__32647));
    InMux I__5482 (
            .O(N__32673),
            .I(N__32644));
    InMux I__5481 (
            .O(N__32672),
            .I(N__32641));
    CascadeMux I__5480 (
            .O(N__32671),
            .I(N__32638));
    LocalMux I__5479 (
            .O(N__32668),
            .I(N__32632));
    InMux I__5478 (
            .O(N__32665),
            .I(N__32627));
    InMux I__5477 (
            .O(N__32664),
            .I(N__32627));
    InMux I__5476 (
            .O(N__32661),
            .I(N__32618));
    InMux I__5475 (
            .O(N__32660),
            .I(N__32618));
    InMux I__5474 (
            .O(N__32657),
            .I(N__32618));
    InMux I__5473 (
            .O(N__32656),
            .I(N__32618));
    CascadeMux I__5472 (
            .O(N__32655),
            .I(N__32615));
    InMux I__5471 (
            .O(N__32654),
            .I(N__32608));
    InMux I__5470 (
            .O(N__32653),
            .I(N__32608));
    InMux I__5469 (
            .O(N__32652),
            .I(N__32605));
    LocalMux I__5468 (
            .O(N__32647),
            .I(N__32602));
    LocalMux I__5467 (
            .O(N__32644),
            .I(N__32597));
    LocalMux I__5466 (
            .O(N__32641),
            .I(N__32597));
    InMux I__5465 (
            .O(N__32638),
            .I(N__32594));
    InMux I__5464 (
            .O(N__32637),
            .I(N__32589));
    InMux I__5463 (
            .O(N__32636),
            .I(N__32589));
    InMux I__5462 (
            .O(N__32635),
            .I(N__32586));
    Span4Mux_v I__5461 (
            .O(N__32632),
            .I(N__32581));
    LocalMux I__5460 (
            .O(N__32627),
            .I(N__32581));
    LocalMux I__5459 (
            .O(N__32618),
            .I(N__32578));
    InMux I__5458 (
            .O(N__32615),
            .I(N__32573));
    InMux I__5457 (
            .O(N__32614),
            .I(N__32573));
    InMux I__5456 (
            .O(N__32613),
            .I(N__32570));
    LocalMux I__5455 (
            .O(N__32608),
            .I(N__32567));
    LocalMux I__5454 (
            .O(N__32605),
            .I(N__32562));
    Span4Mux_h I__5453 (
            .O(N__32602),
            .I(N__32562));
    Span4Mux_v I__5452 (
            .O(N__32597),
            .I(N__32555));
    LocalMux I__5451 (
            .O(N__32594),
            .I(N__32555));
    LocalMux I__5450 (
            .O(N__32589),
            .I(N__32555));
    LocalMux I__5449 (
            .O(N__32586),
            .I(n2247));
    Odrv4 I__5448 (
            .O(N__32581),
            .I(n2247));
    Odrv4 I__5447 (
            .O(N__32578),
            .I(n2247));
    LocalMux I__5446 (
            .O(N__32573),
            .I(n2247));
    LocalMux I__5445 (
            .O(N__32570),
            .I(n2247));
    Odrv4 I__5444 (
            .O(N__32567),
            .I(n2247));
    Odrv4 I__5443 (
            .O(N__32562),
            .I(n2247));
    Odrv4 I__5442 (
            .O(N__32555),
            .I(n2247));
    InMux I__5441 (
            .O(N__32538),
            .I(n12948));
    InMux I__5440 (
            .O(N__32535),
            .I(N__32532));
    LocalMux I__5439 (
            .O(N__32532),
            .I(N__32529));
    Odrv4 I__5438 (
            .O(N__32529),
            .I(n2284));
    CascadeMux I__5437 (
            .O(N__32526),
            .I(N__32523));
    InMux I__5436 (
            .O(N__32523),
            .I(N__32519));
    InMux I__5435 (
            .O(N__32522),
            .I(N__32516));
    LocalMux I__5434 (
            .O(N__32519),
            .I(n2217));
    LocalMux I__5433 (
            .O(N__32516),
            .I(n2217));
    CascadeMux I__5432 (
            .O(N__32511),
            .I(N__32508));
    InMux I__5431 (
            .O(N__32508),
            .I(N__32504));
    CascadeMux I__5430 (
            .O(N__32507),
            .I(N__32501));
    LocalMux I__5429 (
            .O(N__32504),
            .I(N__32497));
    InMux I__5428 (
            .O(N__32501),
            .I(N__32494));
    InMux I__5427 (
            .O(N__32500),
            .I(N__32491));
    Span4Mux_v I__5426 (
            .O(N__32497),
            .I(N__32488));
    LocalMux I__5425 (
            .O(N__32494),
            .I(N__32485));
    LocalMux I__5424 (
            .O(N__32491),
            .I(N__32482));
    Span4Mux_h I__5423 (
            .O(N__32488),
            .I(N__32479));
    Span4Mux_v I__5422 (
            .O(N__32485),
            .I(N__32474));
    Span4Mux_v I__5421 (
            .O(N__32482),
            .I(N__32474));
    Odrv4 I__5420 (
            .O(N__32479),
            .I(n2316));
    Odrv4 I__5419 (
            .O(N__32474),
            .I(n2316));
    InMux I__5418 (
            .O(N__32469),
            .I(N__32466));
    LocalMux I__5417 (
            .O(N__32466),
            .I(N__32463));
    Odrv12 I__5416 (
            .O(N__32463),
            .I(n2100));
    CascadeMux I__5415 (
            .O(N__32460),
            .I(N__32457));
    InMux I__5414 (
            .O(N__32457),
            .I(N__32454));
    LocalMux I__5413 (
            .O(N__32454),
            .I(N__32450));
    InMux I__5412 (
            .O(N__32453),
            .I(N__32446));
    Span12Mux_v I__5411 (
            .O(N__32450),
            .I(N__32443));
    InMux I__5410 (
            .O(N__32449),
            .I(N__32440));
    LocalMux I__5409 (
            .O(N__32446),
            .I(n2132));
    Odrv12 I__5408 (
            .O(N__32443),
            .I(n2132));
    LocalMux I__5407 (
            .O(N__32440),
            .I(n2132));
    InMux I__5406 (
            .O(N__32433),
            .I(N__32429));
    InMux I__5405 (
            .O(N__32432),
            .I(N__32426));
    LocalMux I__5404 (
            .O(N__32429),
            .I(N__32420));
    LocalMux I__5403 (
            .O(N__32426),
            .I(N__32420));
    InMux I__5402 (
            .O(N__32425),
            .I(N__32417));
    Span4Mux_v I__5401 (
            .O(N__32420),
            .I(N__32414));
    LocalMux I__5400 (
            .O(N__32417),
            .I(N__32411));
    Span4Mux_h I__5399 (
            .O(N__32414),
            .I(N__32408));
    Span12Mux_s6_h I__5398 (
            .O(N__32411),
            .I(N__32405));
    Span4Mux_v I__5397 (
            .O(N__32408),
            .I(N__32402));
    Odrv12 I__5396 (
            .O(N__32405),
            .I(n315));
    Odrv4 I__5395 (
            .O(N__32402),
            .I(n315));
    InMux I__5394 (
            .O(N__32397),
            .I(N__32394));
    LocalMux I__5393 (
            .O(N__32394),
            .I(n15484));
    CascadeMux I__5392 (
            .O(N__32391),
            .I(N__32387));
    InMux I__5391 (
            .O(N__32390),
            .I(N__32384));
    InMux I__5390 (
            .O(N__32387),
            .I(N__32381));
    LocalMux I__5389 (
            .O(N__32384),
            .I(n12034));
    LocalMux I__5388 (
            .O(N__32381),
            .I(n12034));
    InMux I__5387 (
            .O(N__32376),
            .I(bfn_7_23_0_));
    InMux I__5386 (
            .O(N__32373),
            .I(n12938));
    InMux I__5385 (
            .O(N__32370),
            .I(N__32367));
    LocalMux I__5384 (
            .O(N__32367),
            .I(N__32363));
    CascadeMux I__5383 (
            .O(N__32366),
            .I(N__32360));
    Span4Mux_v I__5382 (
            .O(N__32363),
            .I(N__32357));
    InMux I__5381 (
            .O(N__32360),
            .I(N__32354));
    Odrv4 I__5380 (
            .O(N__32357),
            .I(n15445));
    LocalMux I__5379 (
            .O(N__32354),
            .I(n15445));
    InMux I__5378 (
            .O(N__32349),
            .I(n12939));
    InMux I__5377 (
            .O(N__32346),
            .I(N__32343));
    LocalMux I__5376 (
            .O(N__32343),
            .I(N__32340));
    Span4Mux_v I__5375 (
            .O(N__32340),
            .I(N__32337));
    Span4Mux_v I__5374 (
            .O(N__32337),
            .I(N__32333));
    CascadeMux I__5373 (
            .O(N__32336),
            .I(N__32330));
    Span4Mux_h I__5372 (
            .O(N__32333),
            .I(N__32327));
    InMux I__5371 (
            .O(N__32330),
            .I(N__32324));
    Odrv4 I__5370 (
            .O(N__32327),
            .I(n15412));
    LocalMux I__5369 (
            .O(N__32324),
            .I(n15412));
    InMux I__5368 (
            .O(N__32319),
            .I(n12940));
    InMux I__5367 (
            .O(N__32316),
            .I(N__32313));
    LocalMux I__5366 (
            .O(N__32313),
            .I(N__32310));
    Span4Mux_v I__5365 (
            .O(N__32310),
            .I(N__32307));
    Span4Mux_v I__5364 (
            .O(N__32307),
            .I(N__32303));
    CascadeMux I__5363 (
            .O(N__32306),
            .I(N__32300));
    Span4Mux_h I__5362 (
            .O(N__32303),
            .I(N__32297));
    InMux I__5361 (
            .O(N__32300),
            .I(N__32294));
    Odrv4 I__5360 (
            .O(N__32297),
            .I(n15378));
    LocalMux I__5359 (
            .O(N__32294),
            .I(n15378));
    CascadeMux I__5358 (
            .O(N__32289),
            .I(N__32286));
    InMux I__5357 (
            .O(N__32286),
            .I(N__32282));
    InMux I__5356 (
            .O(N__32285),
            .I(N__32279));
    LocalMux I__5355 (
            .O(N__32282),
            .I(N__32276));
    LocalMux I__5354 (
            .O(N__32279),
            .I(N__32273));
    Span4Mux_v I__5353 (
            .O(N__32276),
            .I(N__32270));
    Odrv4 I__5352 (
            .O(N__32273),
            .I(n2127));
    Odrv4 I__5351 (
            .O(N__32270),
            .I(n2127));
    CascadeMux I__5350 (
            .O(N__32265),
            .I(N__32262));
    InMux I__5349 (
            .O(N__32262),
            .I(N__32259));
    LocalMux I__5348 (
            .O(N__32259),
            .I(N__32256));
    Span4Mux_v I__5347 (
            .O(N__32256),
            .I(N__32253));
    Odrv4 I__5346 (
            .O(N__32253),
            .I(n2194));
    InMux I__5345 (
            .O(N__32250),
            .I(N__32246));
    CascadeMux I__5344 (
            .O(N__32249),
            .I(N__32243));
    LocalMux I__5343 (
            .O(N__32246),
            .I(N__32240));
    InMux I__5342 (
            .O(N__32243),
            .I(N__32237));
    Span4Mux_v I__5341 (
            .O(N__32240),
            .I(N__32231));
    LocalMux I__5340 (
            .O(N__32237),
            .I(N__32231));
    InMux I__5339 (
            .O(N__32236),
            .I(N__32228));
    Odrv4 I__5338 (
            .O(N__32231),
            .I(n2226));
    LocalMux I__5337 (
            .O(N__32228),
            .I(n2226));
    InMux I__5336 (
            .O(N__32223),
            .I(N__32220));
    LocalMux I__5335 (
            .O(N__32220),
            .I(N__32217));
    Odrv12 I__5334 (
            .O(N__32217),
            .I(n2101));
    CascadeMux I__5333 (
            .O(N__32214),
            .I(N__32211));
    InMux I__5332 (
            .O(N__32211),
            .I(N__32208));
    LocalMux I__5331 (
            .O(N__32208),
            .I(N__32204));
    InMux I__5330 (
            .O(N__32207),
            .I(N__32201));
    Span4Mux_h I__5329 (
            .O(N__32204),
            .I(N__32198));
    LocalMux I__5328 (
            .O(N__32201),
            .I(n2133));
    Odrv4 I__5327 (
            .O(N__32198),
            .I(n2133));
    CascadeMux I__5326 (
            .O(N__32193),
            .I(n2133_cascade_));
    InMux I__5325 (
            .O(N__32190),
            .I(N__32187));
    LocalMux I__5324 (
            .O(N__32187),
            .I(n11892));
    InMux I__5323 (
            .O(N__32184),
            .I(N__32179));
    InMux I__5322 (
            .O(N__32183),
            .I(N__32174));
    InMux I__5321 (
            .O(N__32182),
            .I(N__32174));
    LocalMux I__5320 (
            .O(N__32179),
            .I(N__32171));
    LocalMux I__5319 (
            .O(N__32174),
            .I(N__32168));
    Span4Mux_v I__5318 (
            .O(N__32171),
            .I(N__32165));
    Span4Mux_h I__5317 (
            .O(N__32168),
            .I(N__32162));
    Odrv4 I__5316 (
            .O(N__32165),
            .I(n307));
    Odrv4 I__5315 (
            .O(N__32162),
            .I(n307));
    InMux I__5314 (
            .O(N__32157),
            .I(N__32154));
    LocalMux I__5313 (
            .O(N__32154),
            .I(N__32151));
    Span4Mux_v I__5312 (
            .O(N__32151),
            .I(N__32148));
    Odrv4 I__5311 (
            .O(N__32148),
            .I(n2201));
    CascadeMux I__5310 (
            .O(N__32145),
            .I(N__32142));
    InMux I__5309 (
            .O(N__32142),
            .I(N__32139));
    LocalMux I__5308 (
            .O(N__32139),
            .I(N__32135));
    InMux I__5307 (
            .O(N__32138),
            .I(N__32132));
    Span4Mux_h I__5306 (
            .O(N__32135),
            .I(N__32129));
    LocalMux I__5305 (
            .O(N__32132),
            .I(n2233));
    Odrv4 I__5304 (
            .O(N__32129),
            .I(n2233));
    InMux I__5303 (
            .O(N__32124),
            .I(N__32120));
    CascadeMux I__5302 (
            .O(N__32123),
            .I(N__32117));
    LocalMux I__5301 (
            .O(N__32120),
            .I(N__32113));
    InMux I__5300 (
            .O(N__32117),
            .I(N__32110));
    InMux I__5299 (
            .O(N__32116),
            .I(N__32107));
    Odrv12 I__5298 (
            .O(N__32113),
            .I(n2231));
    LocalMux I__5297 (
            .O(N__32110),
            .I(n2231));
    LocalMux I__5296 (
            .O(N__32107),
            .I(n2231));
    CascadeMux I__5295 (
            .O(N__32100),
            .I(n2233_cascade_));
    CascadeMux I__5294 (
            .O(N__32097),
            .I(N__32093));
    InMux I__5293 (
            .O(N__32096),
            .I(N__32089));
    InMux I__5292 (
            .O(N__32093),
            .I(N__32086));
    InMux I__5291 (
            .O(N__32092),
            .I(N__32083));
    LocalMux I__5290 (
            .O(N__32089),
            .I(n2232));
    LocalMux I__5289 (
            .O(N__32086),
            .I(n2232));
    LocalMux I__5288 (
            .O(N__32083),
            .I(n2232));
    InMux I__5287 (
            .O(N__32076),
            .I(N__32073));
    LocalMux I__5286 (
            .O(N__32073),
            .I(n11950));
    InMux I__5285 (
            .O(N__32070),
            .I(N__32067));
    LocalMux I__5284 (
            .O(N__32067),
            .I(N__32064));
    Odrv4 I__5283 (
            .O(N__32064),
            .I(n2086));
    InMux I__5282 (
            .O(N__32061),
            .I(N__32058));
    LocalMux I__5281 (
            .O(N__32058),
            .I(N__32054));
    InMux I__5280 (
            .O(N__32057),
            .I(N__32050));
    Span4Mux_h I__5279 (
            .O(N__32054),
            .I(N__32047));
    InMux I__5278 (
            .O(N__32053),
            .I(N__32044));
    LocalMux I__5277 (
            .O(N__32050),
            .I(n2118));
    Odrv4 I__5276 (
            .O(N__32047),
            .I(n2118));
    LocalMux I__5275 (
            .O(N__32044),
            .I(n2118));
    InMux I__5274 (
            .O(N__32037),
            .I(N__32033));
    InMux I__5273 (
            .O(N__32036),
            .I(N__32030));
    LocalMux I__5272 (
            .O(N__32033),
            .I(N__32027));
    LocalMux I__5271 (
            .O(N__32030),
            .I(N__32024));
    Span4Mux_v I__5270 (
            .O(N__32027),
            .I(N__32020));
    Span12Mux_s6_h I__5269 (
            .O(N__32024),
            .I(N__32017));
    InMux I__5268 (
            .O(N__32023),
            .I(N__32014));
    Odrv4 I__5267 (
            .O(N__32020),
            .I(n308));
    Odrv12 I__5266 (
            .O(N__32017),
            .I(n308));
    LocalMux I__5265 (
            .O(N__32014),
            .I(n308));
    InMux I__5264 (
            .O(N__32007),
            .I(N__32004));
    LocalMux I__5263 (
            .O(N__32004),
            .I(N__32001));
    Odrv4 I__5262 (
            .O(N__32001),
            .I(n2098));
    CascadeMux I__5261 (
            .O(N__31998),
            .I(N__31995));
    InMux I__5260 (
            .O(N__31995),
            .I(N__31992));
    LocalMux I__5259 (
            .O(N__31992),
            .I(N__31988));
    InMux I__5258 (
            .O(N__31991),
            .I(N__31985));
    Span4Mux_h I__5257 (
            .O(N__31988),
            .I(N__31982));
    LocalMux I__5256 (
            .O(N__31985),
            .I(n2130));
    Odrv4 I__5255 (
            .O(N__31982),
            .I(n2130));
    CascadeMux I__5254 (
            .O(N__31977),
            .I(N__31974));
    InMux I__5253 (
            .O(N__31974),
            .I(N__31971));
    LocalMux I__5252 (
            .O(N__31971),
            .I(N__31966));
    CascadeMux I__5251 (
            .O(N__31970),
            .I(N__31963));
    InMux I__5250 (
            .O(N__31969),
            .I(N__31960));
    Span4Mux_v I__5249 (
            .O(N__31966),
            .I(N__31957));
    InMux I__5248 (
            .O(N__31963),
            .I(N__31954));
    LocalMux I__5247 (
            .O(N__31960),
            .I(N__31951));
    Odrv4 I__5246 (
            .O(N__31957),
            .I(n2131));
    LocalMux I__5245 (
            .O(N__31954),
            .I(n2131));
    Odrv4 I__5244 (
            .O(N__31951),
            .I(n2131));
    CascadeMux I__5243 (
            .O(N__31944),
            .I(N__31941));
    InMux I__5242 (
            .O(N__31941),
            .I(N__31937));
    InMux I__5241 (
            .O(N__31940),
            .I(N__31933));
    LocalMux I__5240 (
            .O(N__31937),
            .I(N__31930));
    CascadeMux I__5239 (
            .O(N__31936),
            .I(N__31927));
    LocalMux I__5238 (
            .O(N__31933),
            .I(N__31924));
    Span4Mux_v I__5237 (
            .O(N__31930),
            .I(N__31921));
    InMux I__5236 (
            .O(N__31927),
            .I(N__31918));
    Span4Mux_v I__5235 (
            .O(N__31924),
            .I(N__31915));
    Odrv4 I__5234 (
            .O(N__31921),
            .I(n2129));
    LocalMux I__5233 (
            .O(N__31918),
            .I(n2129));
    Odrv4 I__5232 (
            .O(N__31915),
            .I(n2129));
    CascadeMux I__5231 (
            .O(N__31908),
            .I(n2130_cascade_));
    InMux I__5230 (
            .O(N__31905),
            .I(N__31900));
    InMux I__5229 (
            .O(N__31904),
            .I(N__31897));
    InMux I__5228 (
            .O(N__31903),
            .I(N__31894));
    LocalMux I__5227 (
            .O(N__31900),
            .I(n2119));
    LocalMux I__5226 (
            .O(N__31897),
            .I(n2119));
    LocalMux I__5225 (
            .O(N__31894),
            .I(n2119));
    CascadeMux I__5224 (
            .O(N__31887),
            .I(n13775_cascade_));
    InMux I__5223 (
            .O(N__31884),
            .I(N__31881));
    LocalMux I__5222 (
            .O(N__31881),
            .I(n14398));
    InMux I__5221 (
            .O(N__31878),
            .I(N__31875));
    LocalMux I__5220 (
            .O(N__31875),
            .I(N__31872));
    Odrv4 I__5219 (
            .O(N__31872),
            .I(n2090));
    CascadeMux I__5218 (
            .O(N__31869),
            .I(N__31866));
    InMux I__5217 (
            .O(N__31866),
            .I(N__31863));
    LocalMux I__5216 (
            .O(N__31863),
            .I(N__31859));
    InMux I__5215 (
            .O(N__31862),
            .I(N__31856));
    Span4Mux_h I__5214 (
            .O(N__31859),
            .I(N__31853));
    LocalMux I__5213 (
            .O(N__31856),
            .I(n2122));
    Odrv4 I__5212 (
            .O(N__31853),
            .I(n2122));
    CascadeMux I__5211 (
            .O(N__31848),
            .I(N__31844));
    InMux I__5210 (
            .O(N__31847),
            .I(N__31840));
    InMux I__5209 (
            .O(N__31844),
            .I(N__31837));
    InMux I__5208 (
            .O(N__31843),
            .I(N__31834));
    LocalMux I__5207 (
            .O(N__31840),
            .I(n2125));
    LocalMux I__5206 (
            .O(N__31837),
            .I(n2125));
    LocalMux I__5205 (
            .O(N__31834),
            .I(n2125));
    CascadeMux I__5204 (
            .O(N__31827),
            .I(n2122_cascade_));
    CascadeMux I__5203 (
            .O(N__31824),
            .I(N__31819));
    CascadeMux I__5202 (
            .O(N__31823),
            .I(N__31816));
    InMux I__5201 (
            .O(N__31822),
            .I(N__31813));
    InMux I__5200 (
            .O(N__31819),
            .I(N__31810));
    InMux I__5199 (
            .O(N__31816),
            .I(N__31807));
    LocalMux I__5198 (
            .O(N__31813),
            .I(N__31804));
    LocalMux I__5197 (
            .O(N__31810),
            .I(n2128));
    LocalMux I__5196 (
            .O(N__31807),
            .I(n2128));
    Odrv4 I__5195 (
            .O(N__31804),
            .I(n2128));
    InMux I__5194 (
            .O(N__31797),
            .I(N__31794));
    LocalMux I__5193 (
            .O(N__31794),
            .I(N__31789));
    InMux I__5192 (
            .O(N__31793),
            .I(N__31786));
    InMux I__5191 (
            .O(N__31792),
            .I(N__31783));
    Odrv4 I__5190 (
            .O(N__31789),
            .I(n2120));
    LocalMux I__5189 (
            .O(N__31786),
            .I(n2120));
    LocalMux I__5188 (
            .O(N__31783),
            .I(n2120));
    CascadeMux I__5187 (
            .O(N__31776),
            .I(n14386_cascade_));
    InMux I__5186 (
            .O(N__31773),
            .I(N__31770));
    LocalMux I__5185 (
            .O(N__31770),
            .I(n14384));
    InMux I__5184 (
            .O(N__31767),
            .I(N__31764));
    LocalMux I__5183 (
            .O(N__31764),
            .I(n14392));
    InMux I__5182 (
            .O(N__31761),
            .I(N__31758));
    LocalMux I__5181 (
            .O(N__31758),
            .I(N__31755));
    Odrv4 I__5180 (
            .O(N__31755),
            .I(n2089));
    InMux I__5179 (
            .O(N__31752),
            .I(N__31748));
    CascadeMux I__5178 (
            .O(N__31751),
            .I(N__31745));
    LocalMux I__5177 (
            .O(N__31748),
            .I(N__31742));
    InMux I__5176 (
            .O(N__31745),
            .I(N__31738));
    Span4Mux_h I__5175 (
            .O(N__31742),
            .I(N__31735));
    InMux I__5174 (
            .O(N__31741),
            .I(N__31732));
    LocalMux I__5173 (
            .O(N__31738),
            .I(n2121));
    Odrv4 I__5172 (
            .O(N__31735),
            .I(n2121));
    LocalMux I__5171 (
            .O(N__31732),
            .I(n2121));
    InMux I__5170 (
            .O(N__31725),
            .I(n12639));
    CascadeMux I__5169 (
            .O(N__31722),
            .I(N__31719));
    InMux I__5168 (
            .O(N__31719),
            .I(N__31716));
    LocalMux I__5167 (
            .O(N__31716),
            .I(n2085));
    InMux I__5166 (
            .O(N__31713),
            .I(bfn_7_19_0_));
    InMux I__5165 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__5164 (
            .O(N__31707),
            .I(n2084));
    InMux I__5163 (
            .O(N__31704),
            .I(n12641));
    InMux I__5162 (
            .O(N__31701),
            .I(n12642));
    CascadeMux I__5161 (
            .O(N__31698),
            .I(N__31695));
    InMux I__5160 (
            .O(N__31695),
            .I(N__31692));
    LocalMux I__5159 (
            .O(N__31692),
            .I(N__31688));
    InMux I__5158 (
            .O(N__31691),
            .I(N__31685));
    Odrv4 I__5157 (
            .O(N__31688),
            .I(n2115));
    LocalMux I__5156 (
            .O(N__31685),
            .I(n2115));
    InMux I__5155 (
            .O(N__31680),
            .I(N__31677));
    LocalMux I__5154 (
            .O(N__31677),
            .I(N__31674));
    Odrv4 I__5153 (
            .O(N__31674),
            .I(n2095));
    InMux I__5152 (
            .O(N__31671),
            .I(N__31667));
    CascadeMux I__5151 (
            .O(N__31670),
            .I(N__31664));
    LocalMux I__5150 (
            .O(N__31667),
            .I(N__31660));
    InMux I__5149 (
            .O(N__31664),
            .I(N__31657));
    InMux I__5148 (
            .O(N__31663),
            .I(N__31654));
    Odrv4 I__5147 (
            .O(N__31660),
            .I(n2123));
    LocalMux I__5146 (
            .O(N__31657),
            .I(n2123));
    LocalMux I__5145 (
            .O(N__31654),
            .I(n2123));
    CascadeMux I__5144 (
            .O(N__31647),
            .I(n2127_cascade_));
    CascadeMux I__5143 (
            .O(N__31644),
            .I(N__31641));
    InMux I__5142 (
            .O(N__31641),
            .I(N__31637));
    InMux I__5141 (
            .O(N__31640),
            .I(N__31634));
    LocalMux I__5140 (
            .O(N__31637),
            .I(n2126));
    LocalMux I__5139 (
            .O(N__31634),
            .I(n2126));
    CascadeMux I__5138 (
            .O(N__31629),
            .I(N__31624));
    InMux I__5137 (
            .O(N__31628),
            .I(N__31621));
    InMux I__5136 (
            .O(N__31627),
            .I(N__31618));
    InMux I__5135 (
            .O(N__31624),
            .I(N__31615));
    LocalMux I__5134 (
            .O(N__31621),
            .I(n2018));
    LocalMux I__5133 (
            .O(N__31618),
            .I(n2018));
    LocalMux I__5132 (
            .O(N__31615),
            .I(n2018));
    CascadeMux I__5131 (
            .O(N__31608),
            .I(N__31605));
    InMux I__5130 (
            .O(N__31605),
            .I(N__31602));
    LocalMux I__5129 (
            .O(N__31602),
            .I(n2092));
    CascadeMux I__5128 (
            .O(N__31599),
            .I(N__31596));
    InMux I__5127 (
            .O(N__31596),
            .I(N__31592));
    InMux I__5126 (
            .O(N__31595),
            .I(N__31589));
    LocalMux I__5125 (
            .O(N__31592),
            .I(N__31586));
    LocalMux I__5124 (
            .O(N__31589),
            .I(N__31580));
    Span4Mux_h I__5123 (
            .O(N__31586),
            .I(N__31580));
    InMux I__5122 (
            .O(N__31585),
            .I(N__31577));
    Odrv4 I__5121 (
            .O(N__31580),
            .I(n2124));
    LocalMux I__5120 (
            .O(N__31577),
            .I(n2124));
    InMux I__5119 (
            .O(N__31572),
            .I(n12630));
    InMux I__5118 (
            .O(N__31569),
            .I(N__31566));
    LocalMux I__5117 (
            .O(N__31566),
            .I(n2094));
    InMux I__5116 (
            .O(N__31563),
            .I(n12631));
    InMux I__5115 (
            .O(N__31560),
            .I(N__31557));
    LocalMux I__5114 (
            .O(N__31557),
            .I(n2093));
    InMux I__5113 (
            .O(N__31554),
            .I(bfn_7_18_0_));
    InMux I__5112 (
            .O(N__31551),
            .I(n12633));
    InMux I__5111 (
            .O(N__31548),
            .I(N__31545));
    LocalMux I__5110 (
            .O(N__31545),
            .I(n2091));
    InMux I__5109 (
            .O(N__31542),
            .I(n12634));
    InMux I__5108 (
            .O(N__31539),
            .I(n12635));
    InMux I__5107 (
            .O(N__31536),
            .I(n12636));
    InMux I__5106 (
            .O(N__31533),
            .I(N__31530));
    LocalMux I__5105 (
            .O(N__31530),
            .I(n2088));
    InMux I__5104 (
            .O(N__31527),
            .I(n12637));
    InMux I__5103 (
            .O(N__31524),
            .I(N__31521));
    LocalMux I__5102 (
            .O(N__31521),
            .I(n2087));
    InMux I__5101 (
            .O(N__31518),
            .I(n12638));
    InMux I__5100 (
            .O(N__31515),
            .I(N__31512));
    LocalMux I__5099 (
            .O(N__31512),
            .I(n14258));
    CascadeMux I__5098 (
            .O(N__31509),
            .I(n14260_cascade_));
    InMux I__5097 (
            .O(N__31506),
            .I(N__31503));
    LocalMux I__5096 (
            .O(N__31503),
            .I(n14262));
    InMux I__5095 (
            .O(N__31500),
            .I(N__31497));
    LocalMux I__5094 (
            .O(N__31497),
            .I(N__31493));
    CascadeMux I__5093 (
            .O(N__31496),
            .I(N__31490));
    Span4Mux_h I__5092 (
            .O(N__31493),
            .I(N__31486));
    InMux I__5091 (
            .O(N__31490),
            .I(N__31483));
    InMux I__5090 (
            .O(N__31489),
            .I(N__31480));
    Odrv4 I__5089 (
            .O(N__31486),
            .I(n3021));
    LocalMux I__5088 (
            .O(N__31483),
            .I(n3021));
    LocalMux I__5087 (
            .O(N__31480),
            .I(n3021));
    CascadeMux I__5086 (
            .O(N__31473),
            .I(N__31470));
    InMux I__5085 (
            .O(N__31470),
            .I(N__31467));
    LocalMux I__5084 (
            .O(N__31467),
            .I(N__31464));
    Span4Mux_s2_v I__5083 (
            .O(N__31464),
            .I(N__31461));
    Odrv4 I__5082 (
            .O(N__31461),
            .I(n3088));
    CascadeMux I__5081 (
            .O(N__31458),
            .I(N__31454));
    CascadeMux I__5080 (
            .O(N__31457),
            .I(N__31451));
    InMux I__5079 (
            .O(N__31454),
            .I(N__31448));
    InMux I__5078 (
            .O(N__31451),
            .I(N__31445));
    LocalMux I__5077 (
            .O(N__31448),
            .I(N__31442));
    LocalMux I__5076 (
            .O(N__31445),
            .I(N__31436));
    Span12Mux_s5_h I__5075 (
            .O(N__31442),
            .I(N__31436));
    InMux I__5074 (
            .O(N__31441),
            .I(N__31433));
    Odrv12 I__5073 (
            .O(N__31436),
            .I(n3120));
    LocalMux I__5072 (
            .O(N__31433),
            .I(n3120));
    InMux I__5071 (
            .O(N__31428),
            .I(bfn_7_17_0_));
    InMux I__5070 (
            .O(N__31425),
            .I(n12625));
    InMux I__5069 (
            .O(N__31422),
            .I(N__31419));
    LocalMux I__5068 (
            .O(N__31419),
            .I(n2099));
    InMux I__5067 (
            .O(N__31416),
            .I(n12626));
    InMux I__5066 (
            .O(N__31413),
            .I(n12627));
    InMux I__5065 (
            .O(N__31410),
            .I(N__31407));
    LocalMux I__5064 (
            .O(N__31407),
            .I(n2097));
    InMux I__5063 (
            .O(N__31404),
            .I(n12628));
    InMux I__5062 (
            .O(N__31401),
            .I(N__31398));
    LocalMux I__5061 (
            .O(N__31398),
            .I(n2096));
    InMux I__5060 (
            .O(N__31395),
            .I(n12629));
    CascadeMux I__5059 (
            .O(N__31392),
            .I(n14250_cascade_));
    InMux I__5058 (
            .O(N__31389),
            .I(N__31386));
    LocalMux I__5057 (
            .O(N__31386),
            .I(N__31381));
    InMux I__5056 (
            .O(N__31385),
            .I(N__31378));
    InMux I__5055 (
            .O(N__31384),
            .I(N__31375));
    Span4Mux_h I__5054 (
            .O(N__31381),
            .I(N__31370));
    LocalMux I__5053 (
            .O(N__31378),
            .I(N__31370));
    LocalMux I__5052 (
            .O(N__31375),
            .I(N__31367));
    Odrv4 I__5051 (
            .O(N__31370),
            .I(n3026));
    Odrv4 I__5050 (
            .O(N__31367),
            .I(n3026));
    CascadeMux I__5049 (
            .O(N__31362),
            .I(N__31359));
    InMux I__5048 (
            .O(N__31359),
            .I(N__31356));
    LocalMux I__5047 (
            .O(N__31356),
            .I(N__31353));
    Span4Mux_s2_v I__5046 (
            .O(N__31353),
            .I(N__31350));
    Odrv4 I__5045 (
            .O(N__31350),
            .I(n3093));
    CascadeMux I__5044 (
            .O(N__31347),
            .I(N__31344));
    InMux I__5043 (
            .O(N__31344),
            .I(N__31341));
    LocalMux I__5042 (
            .O(N__31341),
            .I(N__31338));
    Span4Mux_v I__5041 (
            .O(N__31338),
            .I(N__31335));
    Odrv4 I__5040 (
            .O(N__31335),
            .I(n59));
    InMux I__5039 (
            .O(N__31332),
            .I(N__31329));
    LocalMux I__5038 (
            .O(N__31329),
            .I(n14252));
    InMux I__5037 (
            .O(N__31326),
            .I(N__31323));
    LocalMux I__5036 (
            .O(N__31323),
            .I(n5_adj_703));
    CascadeMux I__5035 (
            .O(N__31320),
            .I(n14254_cascade_));
    InMux I__5034 (
            .O(N__31317),
            .I(N__31314));
    LocalMux I__5033 (
            .O(N__31314),
            .I(N__31311));
    Odrv4 I__5032 (
            .O(N__31311),
            .I(n11926));
    CascadeMux I__5031 (
            .O(N__31308),
            .I(n14256_cascade_));
    InMux I__5030 (
            .O(N__31305),
            .I(N__31302));
    LocalMux I__5029 (
            .O(N__31302),
            .I(n7_adj_708));
    CascadeMux I__5028 (
            .O(N__31299),
            .I(n14264_cascade_));
    InMux I__5027 (
            .O(N__31296),
            .I(N__31293));
    LocalMux I__5026 (
            .O(N__31293),
            .I(N__31290));
    Span4Mux_v I__5025 (
            .O(N__31290),
            .I(N__31287));
    Odrv4 I__5024 (
            .O(N__31287),
            .I(n14266));
    InMux I__5023 (
            .O(N__31284),
            .I(N__31281));
    LocalMux I__5022 (
            .O(N__31281),
            .I(N__31278));
    Odrv12 I__5021 (
            .O(N__31278),
            .I(n3101));
    InMux I__5020 (
            .O(N__31275),
            .I(N__31272));
    LocalMux I__5019 (
            .O(N__31272),
            .I(N__31269));
    Span4Mux_v I__5018 (
            .O(N__31269),
            .I(N__31266));
    Odrv4 I__5017 (
            .O(N__31266),
            .I(n3200));
    CascadeMux I__5016 (
            .O(N__31263),
            .I(n3133_cascade_));
    CascadeMux I__5015 (
            .O(N__31260),
            .I(n3232_cascade_));
    CascadeMux I__5014 (
            .O(N__31257),
            .I(n25_adj_712_cascade_));
    InMux I__5013 (
            .O(N__31254),
            .I(N__31251));
    LocalMux I__5012 (
            .O(N__31251),
            .I(n37_adj_715));
    InMux I__5011 (
            .O(N__31248),
            .I(N__31245));
    LocalMux I__5010 (
            .O(N__31245),
            .I(n14234));
    CascadeMux I__5009 (
            .O(N__31242),
            .I(n14238_cascade_));
    InMux I__5008 (
            .O(N__31239),
            .I(N__31236));
    LocalMux I__5007 (
            .O(N__31236),
            .I(N__31233));
    Odrv12 I__5006 (
            .O(N__31233),
            .I(n14248));
    InMux I__5005 (
            .O(N__31230),
            .I(N__31227));
    LocalMux I__5004 (
            .O(N__31227),
            .I(N__31224));
    Span4Mux_v I__5003 (
            .O(N__31224),
            .I(N__31221));
    Span4Mux_h I__5002 (
            .O(N__31221),
            .I(N__31218));
    Odrv4 I__5001 (
            .O(N__31218),
            .I(n3201));
    InMux I__5000 (
            .O(N__31215),
            .I(N__31212));
    LocalMux I__4999 (
            .O(N__31212),
            .I(N__31209));
    Odrv4 I__4998 (
            .O(N__31209),
            .I(n11861));
    CascadeMux I__4997 (
            .O(N__31206),
            .I(n3233_cascade_));
    InMux I__4996 (
            .O(N__31203),
            .I(N__31196));
    InMux I__4995 (
            .O(N__31202),
            .I(N__31196));
    InMux I__4994 (
            .O(N__31201),
            .I(N__31193));
    LocalMux I__4993 (
            .O(N__31196),
            .I(N__31190));
    LocalMux I__4992 (
            .O(N__31193),
            .I(N__31187));
    Span4Mux_v I__4991 (
            .O(N__31190),
            .I(N__31184));
    Odrv12 I__4990 (
            .O(N__31187),
            .I(n3111));
    Odrv4 I__4989 (
            .O(N__31184),
            .I(n3111));
    CascadeMux I__4988 (
            .O(N__31179),
            .I(N__31176));
    InMux I__4987 (
            .O(N__31176),
            .I(N__31173));
    LocalMux I__4986 (
            .O(N__31173),
            .I(n3178));
    InMux I__4985 (
            .O(N__31170),
            .I(N__31166));
    CascadeMux I__4984 (
            .O(N__31169),
            .I(N__31163));
    LocalMux I__4983 (
            .O(N__31166),
            .I(N__31160));
    InMux I__4982 (
            .O(N__31163),
            .I(N__31157));
    Odrv4 I__4981 (
            .O(N__31160),
            .I(n3023));
    LocalMux I__4980 (
            .O(N__31157),
            .I(n3023));
    InMux I__4979 (
            .O(N__31152),
            .I(N__31149));
    LocalMux I__4978 (
            .O(N__31149),
            .I(N__31146));
    Span4Mux_h I__4977 (
            .O(N__31146),
            .I(N__31143));
    Odrv4 I__4976 (
            .O(N__31143),
            .I(n3090));
    InMux I__4975 (
            .O(N__31140),
            .I(N__31135));
    InMux I__4974 (
            .O(N__31139),
            .I(N__31132));
    InMux I__4973 (
            .O(N__31138),
            .I(N__31129));
    LocalMux I__4972 (
            .O(N__31135),
            .I(N__31126));
    LocalMux I__4971 (
            .O(N__31132),
            .I(N__31121));
    LocalMux I__4970 (
            .O(N__31129),
            .I(N__31121));
    Span4Mux_s1_v I__4969 (
            .O(N__31126),
            .I(N__31118));
    Odrv4 I__4968 (
            .O(N__31121),
            .I(n3122));
    Odrv4 I__4967 (
            .O(N__31118),
            .I(n3122));
    InMux I__4966 (
            .O(N__31113),
            .I(N__31110));
    LocalMux I__4965 (
            .O(N__31110),
            .I(N__31107));
    Odrv4 I__4964 (
            .O(N__31107),
            .I(n3181));
    CascadeMux I__4963 (
            .O(N__31104),
            .I(N__31101));
    InMux I__4962 (
            .O(N__31101),
            .I(N__31098));
    LocalMux I__4961 (
            .O(N__31098),
            .I(N__31095));
    Span4Mux_v I__4960 (
            .O(N__31095),
            .I(N__31092));
    Odrv4 I__4959 (
            .O(N__31092),
            .I(n3199));
    InMux I__4958 (
            .O(N__31089),
            .I(N__31086));
    LocalMux I__4957 (
            .O(N__31086),
            .I(N__31083));
    Span4Mux_v I__4956 (
            .O(N__31083),
            .I(N__31080));
    Odrv4 I__4955 (
            .O(N__31080),
            .I(n3198));
    InMux I__4954 (
            .O(N__31077),
            .I(N__31073));
    InMux I__4953 (
            .O(N__31076),
            .I(N__31069));
    LocalMux I__4952 (
            .O(N__31073),
            .I(N__31066));
    InMux I__4951 (
            .O(N__31072),
            .I(N__31063));
    LocalMux I__4950 (
            .O(N__31069),
            .I(N__31060));
    Span4Mux_v I__4949 (
            .O(N__31066),
            .I(N__31055));
    LocalMux I__4948 (
            .O(N__31063),
            .I(N__31055));
    Odrv4 I__4947 (
            .O(N__31060),
            .I(n3115));
    Odrv4 I__4946 (
            .O(N__31055),
            .I(n3115));
    InMux I__4945 (
            .O(N__31050),
            .I(N__31047));
    LocalMux I__4944 (
            .O(N__31047),
            .I(N__31043));
    InMux I__4943 (
            .O(N__31046),
            .I(N__31039));
    Span4Mux_h I__4942 (
            .O(N__31043),
            .I(N__31036));
    InMux I__4941 (
            .O(N__31042),
            .I(N__31033));
    LocalMux I__4940 (
            .O(N__31039),
            .I(n3114));
    Odrv4 I__4939 (
            .O(N__31036),
            .I(n3114));
    LocalMux I__4938 (
            .O(N__31033),
            .I(n3114));
    InMux I__4937 (
            .O(N__31026),
            .I(N__31023));
    LocalMux I__4936 (
            .O(N__31023),
            .I(N__31020));
    Odrv4 I__4935 (
            .O(N__31020),
            .I(n14204));
    InMux I__4934 (
            .O(N__31017),
            .I(N__31014));
    LocalMux I__4933 (
            .O(N__31014),
            .I(n14210));
    InMux I__4932 (
            .O(N__31011),
            .I(N__31008));
    LocalMux I__4931 (
            .O(N__31008),
            .I(n3175));
    CascadeMux I__4930 (
            .O(N__31005),
            .I(N__31001));
    InMux I__4929 (
            .O(N__31004),
            .I(N__30998));
    InMux I__4928 (
            .O(N__31001),
            .I(N__30995));
    LocalMux I__4927 (
            .O(N__30998),
            .I(N__30992));
    LocalMux I__4926 (
            .O(N__30995),
            .I(N__30989));
    Span4Mux_h I__4925 (
            .O(N__30992),
            .I(N__30985));
    Span4Mux_v I__4924 (
            .O(N__30989),
            .I(N__30982));
    InMux I__4923 (
            .O(N__30988),
            .I(N__30979));
    Odrv4 I__4922 (
            .O(N__30985),
            .I(n3121));
    Odrv4 I__4921 (
            .O(N__30982),
            .I(n3121));
    LocalMux I__4920 (
            .O(N__30979),
            .I(n3121));
    CascadeMux I__4919 (
            .O(N__30972),
            .I(N__30969));
    InMux I__4918 (
            .O(N__30969),
            .I(N__30966));
    LocalMux I__4917 (
            .O(N__30966),
            .I(n3188));
    InMux I__4916 (
            .O(N__30963),
            .I(N__30960));
    LocalMux I__4915 (
            .O(N__30960),
            .I(n3191));
    InMux I__4914 (
            .O(N__30957),
            .I(N__30954));
    LocalMux I__4913 (
            .O(N__30954),
            .I(N__30950));
    InMux I__4912 (
            .O(N__30953),
            .I(N__30947));
    Span4Mux_v I__4911 (
            .O(N__30950),
            .I(N__30943));
    LocalMux I__4910 (
            .O(N__30947),
            .I(N__30940));
    InMux I__4909 (
            .O(N__30946),
            .I(N__30937));
    Odrv4 I__4908 (
            .O(N__30943),
            .I(n3124));
    Odrv12 I__4907 (
            .O(N__30940),
            .I(n3124));
    LocalMux I__4906 (
            .O(N__30937),
            .I(n3124));
    CascadeMux I__4905 (
            .O(N__30930),
            .I(N__30927));
    InMux I__4904 (
            .O(N__30927),
            .I(N__30924));
    LocalMux I__4903 (
            .O(N__30924),
            .I(n3179));
    InMux I__4902 (
            .O(N__30921),
            .I(N__30916));
    CascadeMux I__4901 (
            .O(N__30920),
            .I(N__30913));
    InMux I__4900 (
            .O(N__30919),
            .I(N__30910));
    LocalMux I__4899 (
            .O(N__30916),
            .I(N__30907));
    InMux I__4898 (
            .O(N__30913),
            .I(N__30904));
    LocalMux I__4897 (
            .O(N__30910),
            .I(n3113));
    Odrv4 I__4896 (
            .O(N__30907),
            .I(n3113));
    LocalMux I__4895 (
            .O(N__30904),
            .I(n3113));
    InMux I__4894 (
            .O(N__30897),
            .I(N__30894));
    LocalMux I__4893 (
            .O(N__30894),
            .I(N__30889));
    InMux I__4892 (
            .O(N__30893),
            .I(N__30886));
    InMux I__4891 (
            .O(N__30892),
            .I(N__30883));
    Odrv4 I__4890 (
            .O(N__30889),
            .I(n3108));
    LocalMux I__4889 (
            .O(N__30886),
            .I(n3108));
    LocalMux I__4888 (
            .O(N__30883),
            .I(n3108));
    CascadeMux I__4887 (
            .O(N__30876),
            .I(n14216_cascade_));
    InMux I__4886 (
            .O(N__30873),
            .I(N__30869));
    InMux I__4885 (
            .O(N__30872),
            .I(N__30866));
    LocalMux I__4884 (
            .O(N__30869),
            .I(N__30861));
    LocalMux I__4883 (
            .O(N__30866),
            .I(N__30861));
    Span4Mux_h I__4882 (
            .O(N__30861),
            .I(N__30858));
    Odrv4 I__4881 (
            .O(N__30858),
            .I(n3105));
    CascadeMux I__4880 (
            .O(N__30855),
            .I(n14222_cascade_));
    InMux I__4879 (
            .O(N__30852),
            .I(N__30849));
    LocalMux I__4878 (
            .O(N__30849),
            .I(N__30844));
    InMux I__4877 (
            .O(N__30848),
            .I(N__30841));
    InMux I__4876 (
            .O(N__30847),
            .I(N__30838));
    Span4Mux_v I__4875 (
            .O(N__30844),
            .I(N__30835));
    LocalMux I__4874 (
            .O(N__30841),
            .I(N__30830));
    LocalMux I__4873 (
            .O(N__30838),
            .I(N__30830));
    Span4Mux_v I__4872 (
            .O(N__30835),
            .I(N__30827));
    Span4Mux_h I__4871 (
            .O(N__30830),
            .I(N__30824));
    Odrv4 I__4870 (
            .O(N__30827),
            .I(n3106));
    Odrv4 I__4869 (
            .O(N__30824),
            .I(n3106));
    CascadeMux I__4868 (
            .O(N__30819),
            .I(n3138_cascade_));
    InMux I__4867 (
            .O(N__30816),
            .I(N__30811));
    InMux I__4866 (
            .O(N__30815),
            .I(N__30806));
    InMux I__4865 (
            .O(N__30814),
            .I(N__30806));
    LocalMux I__4864 (
            .O(N__30811),
            .I(N__30801));
    LocalMux I__4863 (
            .O(N__30806),
            .I(N__30801));
    Span4Mux_h I__4862 (
            .O(N__30801),
            .I(N__30798));
    Odrv4 I__4861 (
            .O(N__30798),
            .I(n3107));
    InMux I__4860 (
            .O(N__30795),
            .I(N__30792));
    LocalMux I__4859 (
            .O(N__30792),
            .I(n3174));
    CascadeMux I__4858 (
            .O(N__30789),
            .I(n3214_cascade_));
    CascadeMux I__4857 (
            .O(N__30786),
            .I(N__30783));
    InMux I__4856 (
            .O(N__30783),
            .I(N__30780));
    LocalMux I__4855 (
            .O(N__30780),
            .I(n3190));
    CascadeMux I__4854 (
            .O(N__30777),
            .I(n3222_cascade_));
    InMux I__4853 (
            .O(N__30774),
            .I(N__30771));
    LocalMux I__4852 (
            .O(N__30771),
            .I(n27_adj_713));
    InMux I__4851 (
            .O(N__30768),
            .I(N__30765));
    LocalMux I__4850 (
            .O(N__30765),
            .I(n3183));
    CascadeMux I__4849 (
            .O(N__30762),
            .I(N__30759));
    InMux I__4848 (
            .O(N__30759),
            .I(N__30756));
    LocalMux I__4847 (
            .O(N__30756),
            .I(N__30752));
    InMux I__4846 (
            .O(N__30755),
            .I(N__30749));
    Span4Mux_v I__4845 (
            .O(N__30752),
            .I(N__30745));
    LocalMux I__4844 (
            .O(N__30749),
            .I(N__30742));
    InMux I__4843 (
            .O(N__30748),
            .I(N__30739));
    Odrv4 I__4842 (
            .O(N__30745),
            .I(n3116));
    Odrv12 I__4841 (
            .O(N__30742),
            .I(n3116));
    LocalMux I__4840 (
            .O(N__30739),
            .I(n3116));
    InMux I__4839 (
            .O(N__30732),
            .I(N__30729));
    LocalMux I__4838 (
            .O(N__30729),
            .I(n14794));
    InMux I__4837 (
            .O(N__30726),
            .I(N__30723));
    LocalMux I__4836 (
            .O(N__30723),
            .I(n14800));
    InMux I__4835 (
            .O(N__30720),
            .I(N__30717));
    LocalMux I__4834 (
            .O(N__30717),
            .I(N__30714));
    Odrv12 I__4833 (
            .O(N__30714),
            .I(n2891));
    CascadeMux I__4832 (
            .O(N__30711),
            .I(N__30707));
    CascadeMux I__4831 (
            .O(N__30710),
            .I(N__30704));
    InMux I__4830 (
            .O(N__30707),
            .I(N__30701));
    InMux I__4829 (
            .O(N__30704),
            .I(N__30698));
    LocalMux I__4828 (
            .O(N__30701),
            .I(N__30694));
    LocalMux I__4827 (
            .O(N__30698),
            .I(N__30691));
    CascadeMux I__4826 (
            .O(N__30697),
            .I(N__30688));
    Span4Mux_v I__4825 (
            .O(N__30694),
            .I(N__30685));
    Span4Mux_v I__4824 (
            .O(N__30691),
            .I(N__30682));
    InMux I__4823 (
            .O(N__30688),
            .I(N__30679));
    Odrv4 I__4822 (
            .O(N__30685),
            .I(n2824));
    Odrv4 I__4821 (
            .O(N__30682),
            .I(n2824));
    LocalMux I__4820 (
            .O(N__30679),
            .I(n2824));
    InMux I__4819 (
            .O(N__30672),
            .I(N__30668));
    InMux I__4818 (
            .O(N__30671),
            .I(N__30665));
    LocalMux I__4817 (
            .O(N__30668),
            .I(N__30661));
    LocalMux I__4816 (
            .O(N__30665),
            .I(N__30658));
    InMux I__4815 (
            .O(N__30664),
            .I(N__30655));
    Span4Mux_s3_v I__4814 (
            .O(N__30661),
            .I(N__30652));
    Span12Mux_s5_v I__4813 (
            .O(N__30658),
            .I(N__30649));
    LocalMux I__4812 (
            .O(N__30655),
            .I(N__30646));
    Odrv4 I__4811 (
            .O(N__30652),
            .I(n2923));
    Odrv12 I__4810 (
            .O(N__30649),
            .I(n2923));
    Odrv4 I__4809 (
            .O(N__30646),
            .I(n2923));
    InMux I__4808 (
            .O(N__30639),
            .I(N__30636));
    LocalMux I__4807 (
            .O(N__30636),
            .I(n3187));
    InMux I__4806 (
            .O(N__30633),
            .I(N__30630));
    LocalMux I__4805 (
            .O(N__30630),
            .I(n3189));
    CascadeMux I__4804 (
            .O(N__30627),
            .I(n3221_cascade_));
    CascadeMux I__4803 (
            .O(N__30624),
            .I(n14268_cascade_));
    CascadeMux I__4802 (
            .O(N__30621),
            .I(n14806_cascade_));
    CascadeMux I__4801 (
            .O(N__30618),
            .I(n3237_cascade_));
    InMux I__4800 (
            .O(N__30615),
            .I(N__30612));
    LocalMux I__4799 (
            .O(N__30612),
            .I(n14228));
    InMux I__4798 (
            .O(N__30609),
            .I(N__30606));
    LocalMux I__4797 (
            .O(N__30606),
            .I(n14270));
    InMux I__4796 (
            .O(N__30603),
            .I(N__30600));
    LocalMux I__4795 (
            .O(N__30600),
            .I(n14272));
    InMux I__4794 (
            .O(N__30597),
            .I(N__30594));
    LocalMux I__4793 (
            .O(N__30594),
            .I(N__30591));
    Odrv4 I__4792 (
            .O(N__30591),
            .I(n3173));
    CascadeMux I__4791 (
            .O(N__30588),
            .I(N__30585));
    InMux I__4790 (
            .O(N__30585),
            .I(N__30582));
    LocalMux I__4789 (
            .O(N__30582),
            .I(n3182));
    InMux I__4788 (
            .O(N__30579),
            .I(N__30575));
    InMux I__4787 (
            .O(N__30578),
            .I(N__30572));
    LocalMux I__4786 (
            .O(N__30575),
            .I(N__30569));
    LocalMux I__4785 (
            .O(N__30572),
            .I(N__30566));
    Span4Mux_h I__4784 (
            .O(N__30569),
            .I(N__30562));
    Span4Mux_v I__4783 (
            .O(N__30566),
            .I(N__30559));
    InMux I__4782 (
            .O(N__30565),
            .I(N__30556));
    Span4Mux_v I__4781 (
            .O(N__30562),
            .I(N__30553));
    Span4Mux_v I__4780 (
            .O(N__30559),
            .I(N__30548));
    LocalMux I__4779 (
            .O(N__30556),
            .I(N__30548));
    Odrv4 I__4778 (
            .O(N__30553),
            .I(n309));
    Odrv4 I__4777 (
            .O(N__30548),
            .I(n309));
    CascadeMux I__4776 (
            .O(N__30543),
            .I(n17_adj_710_cascade_));
    CascadeMux I__4775 (
            .O(N__30540),
            .I(n19_adj_711_cascade_));
    InMux I__4774 (
            .O(N__30537),
            .I(N__30534));
    LocalMux I__4773 (
            .O(N__30534),
            .I(n14236));
    CascadeMux I__4772 (
            .O(N__30531),
            .I(n14230_cascade_));
    InMux I__4771 (
            .O(N__30528),
            .I(N__30525));
    LocalMux I__4770 (
            .O(N__30525),
            .I(n61));
    CascadeMux I__4769 (
            .O(N__30522),
            .I(N__30519));
    InMux I__4768 (
            .O(N__30519),
            .I(N__30516));
    LocalMux I__4767 (
            .O(N__30516),
            .I(N__30513));
    Span4Mux_v I__4766 (
            .O(N__30513),
            .I(N__30510));
    Odrv4 I__4765 (
            .O(N__30510),
            .I(n2190));
    InMux I__4764 (
            .O(N__30507),
            .I(N__30503));
    CascadeMux I__4763 (
            .O(N__30506),
            .I(N__30500));
    LocalMux I__4762 (
            .O(N__30503),
            .I(N__30496));
    InMux I__4761 (
            .O(N__30500),
            .I(N__30493));
    CascadeMux I__4760 (
            .O(N__30499),
            .I(N__30490));
    Span4Mux_v I__4759 (
            .O(N__30496),
            .I(N__30487));
    LocalMux I__4758 (
            .O(N__30493),
            .I(N__30484));
    InMux I__4757 (
            .O(N__30490),
            .I(N__30481));
    Odrv4 I__4756 (
            .O(N__30487),
            .I(n2228));
    Odrv4 I__4755 (
            .O(N__30484),
            .I(n2228));
    LocalMux I__4754 (
            .O(N__30481),
            .I(n2228));
    CascadeMux I__4753 (
            .O(N__30474),
            .I(N__30471));
    InMux I__4752 (
            .O(N__30471),
            .I(N__30468));
    LocalMux I__4751 (
            .O(N__30468),
            .I(N__30464));
    InMux I__4750 (
            .O(N__30467),
            .I(N__30461));
    Sp12to4 I__4749 (
            .O(N__30464),
            .I(N__30456));
    LocalMux I__4748 (
            .O(N__30461),
            .I(N__30456));
    Odrv12 I__4747 (
            .O(N__30456),
            .I(n2224));
    CascadeMux I__4746 (
            .O(N__30453),
            .I(N__30448));
    InMux I__4745 (
            .O(N__30452),
            .I(N__30445));
    InMux I__4744 (
            .O(N__30451),
            .I(N__30442));
    InMux I__4743 (
            .O(N__30448),
            .I(N__30439));
    LocalMux I__4742 (
            .O(N__30445),
            .I(N__30436));
    LocalMux I__4741 (
            .O(N__30442),
            .I(n2227));
    LocalMux I__4740 (
            .O(N__30439),
            .I(n2227));
    Odrv4 I__4739 (
            .O(N__30436),
            .I(n2227));
    CascadeMux I__4738 (
            .O(N__30429),
            .I(n14578_cascade_));
    CascadeMux I__4737 (
            .O(N__30426),
            .I(N__30423));
    InMux I__4736 (
            .O(N__30423),
            .I(N__30419));
    InMux I__4735 (
            .O(N__30422),
            .I(N__30416));
    LocalMux I__4734 (
            .O(N__30419),
            .I(N__30413));
    LocalMux I__4733 (
            .O(N__30416),
            .I(N__30410));
    Odrv4 I__4732 (
            .O(N__30413),
            .I(n2225));
    Odrv12 I__4731 (
            .O(N__30410),
            .I(n2225));
    CascadeMux I__4730 (
            .O(N__30405),
            .I(N__30400));
    InMux I__4729 (
            .O(N__30404),
            .I(N__30397));
    InMux I__4728 (
            .O(N__30403),
            .I(N__30394));
    InMux I__4727 (
            .O(N__30400),
            .I(N__30391));
    LocalMux I__4726 (
            .O(N__30397),
            .I(N__30388));
    LocalMux I__4725 (
            .O(N__30394),
            .I(n2223));
    LocalMux I__4724 (
            .O(N__30391),
            .I(n2223));
    Odrv4 I__4723 (
            .O(N__30388),
            .I(n2223));
    CascadeMux I__4722 (
            .O(N__30381),
            .I(N__30377));
    InMux I__4721 (
            .O(N__30380),
            .I(N__30373));
    InMux I__4720 (
            .O(N__30377),
            .I(N__30370));
    InMux I__4719 (
            .O(N__30376),
            .I(N__30367));
    LocalMux I__4718 (
            .O(N__30373),
            .I(n2222));
    LocalMux I__4717 (
            .O(N__30370),
            .I(n2222));
    LocalMux I__4716 (
            .O(N__30367),
            .I(n2222));
    CascadeMux I__4715 (
            .O(N__30360),
            .I(n14582_cascade_));
    CascadeMux I__4714 (
            .O(N__30357),
            .I(N__30354));
    InMux I__4713 (
            .O(N__30354),
            .I(N__30349));
    CascadeMux I__4712 (
            .O(N__30353),
            .I(N__30346));
    InMux I__4711 (
            .O(N__30352),
            .I(N__30343));
    LocalMux I__4710 (
            .O(N__30349),
            .I(N__30340));
    InMux I__4709 (
            .O(N__30346),
            .I(N__30337));
    LocalMux I__4708 (
            .O(N__30343),
            .I(N__30334));
    Odrv4 I__4707 (
            .O(N__30340),
            .I(n2221));
    LocalMux I__4706 (
            .O(N__30337),
            .I(n2221));
    Odrv4 I__4705 (
            .O(N__30334),
            .I(n2221));
    InMux I__4704 (
            .O(N__30327),
            .I(N__30324));
    LocalMux I__4703 (
            .O(N__30324),
            .I(N__30321));
    Span4Mux_h I__4702 (
            .O(N__30321),
            .I(N__30316));
    InMux I__4701 (
            .O(N__30320),
            .I(N__30313));
    InMux I__4700 (
            .O(N__30319),
            .I(N__30310));
    Odrv4 I__4699 (
            .O(N__30316),
            .I(n2220));
    LocalMux I__4698 (
            .O(N__30313),
            .I(n2220));
    LocalMux I__4697 (
            .O(N__30310),
            .I(n2220));
    CascadeMux I__4696 (
            .O(N__30303),
            .I(n14588_cascade_));
    InMux I__4695 (
            .O(N__30300),
            .I(N__30297));
    LocalMux I__4694 (
            .O(N__30297),
            .I(N__30294));
    Odrv4 I__4693 (
            .O(N__30294),
            .I(n14812));
    InMux I__4692 (
            .O(N__30291),
            .I(N__30288));
    LocalMux I__4691 (
            .O(N__30288),
            .I(n14592));
    InMux I__4690 (
            .O(N__30285),
            .I(N__30282));
    LocalMux I__4689 (
            .O(N__30282),
            .I(N__30279));
    Odrv4 I__4688 (
            .O(N__30279),
            .I(n2187));
    CascadeMux I__4687 (
            .O(N__30276),
            .I(N__30273));
    InMux I__4686 (
            .O(N__30273),
            .I(N__30270));
    LocalMux I__4685 (
            .O(N__30270),
            .I(N__30267));
    Span4Mux_v I__4684 (
            .O(N__30267),
            .I(N__30264));
    Odrv4 I__4683 (
            .O(N__30264),
            .I(n2199));
    CascadeMux I__4682 (
            .O(N__30261),
            .I(N__30258));
    InMux I__4681 (
            .O(N__30258),
            .I(N__30255));
    LocalMux I__4680 (
            .O(N__30255),
            .I(n2285));
    CascadeMux I__4679 (
            .O(N__30252),
            .I(N__30248));
    CascadeMux I__4678 (
            .O(N__30251),
            .I(N__30244));
    InMux I__4677 (
            .O(N__30248),
            .I(N__30241));
    InMux I__4676 (
            .O(N__30247),
            .I(N__30238));
    InMux I__4675 (
            .O(N__30244),
            .I(N__30235));
    LocalMux I__4674 (
            .O(N__30241),
            .I(N__30232));
    LocalMux I__4673 (
            .O(N__30238),
            .I(N__30227));
    LocalMux I__4672 (
            .O(N__30235),
            .I(N__30227));
    Span4Mux_v I__4671 (
            .O(N__30232),
            .I(N__30224));
    Span4Mux_v I__4670 (
            .O(N__30227),
            .I(N__30221));
    Odrv4 I__4669 (
            .O(N__30224),
            .I(n2317));
    Odrv4 I__4668 (
            .O(N__30221),
            .I(n2317));
    CascadeMux I__4667 (
            .O(N__30216),
            .I(N__30213));
    InMux I__4666 (
            .O(N__30213),
            .I(N__30210));
    LocalMux I__4665 (
            .O(N__30210),
            .I(N__30207));
    Span4Mux_v I__4664 (
            .O(N__30207),
            .I(N__30204));
    Odrv4 I__4663 (
            .O(N__30204),
            .I(n2200));
    InMux I__4662 (
            .O(N__30201),
            .I(N__30198));
    LocalMux I__4661 (
            .O(N__30198),
            .I(N__30195));
    Odrv4 I__4660 (
            .O(N__30195),
            .I(n2191));
    CascadeMux I__4659 (
            .O(N__30192),
            .I(N__30189));
    InMux I__4658 (
            .O(N__30189),
            .I(N__30186));
    LocalMux I__4657 (
            .O(N__30186),
            .I(N__30183));
    Span4Mux_v I__4656 (
            .O(N__30183),
            .I(N__30180));
    Odrv4 I__4655 (
            .O(N__30180),
            .I(n2185));
    CascadeMux I__4654 (
            .O(N__30177),
            .I(N__30174));
    InMux I__4653 (
            .O(N__30174),
            .I(N__30169));
    InMux I__4652 (
            .O(N__30173),
            .I(N__30164));
    InMux I__4651 (
            .O(N__30172),
            .I(N__30164));
    LocalMux I__4650 (
            .O(N__30169),
            .I(N__30161));
    LocalMux I__4649 (
            .O(N__30164),
            .I(N__30158));
    Odrv4 I__4648 (
            .O(N__30161),
            .I(n2218));
    Odrv4 I__4647 (
            .O(N__30158),
            .I(n2218));
    InMux I__4646 (
            .O(N__30153),
            .I(N__30150));
    LocalMux I__4645 (
            .O(N__30150),
            .I(N__30147));
    Span4Mux_v I__4644 (
            .O(N__30147),
            .I(N__30142));
    InMux I__4643 (
            .O(N__30146),
            .I(N__30139));
    InMux I__4642 (
            .O(N__30145),
            .I(N__30136));
    Odrv4 I__4641 (
            .O(N__30142),
            .I(n2219));
    LocalMux I__4640 (
            .O(N__30139),
            .I(n2219));
    LocalMux I__4639 (
            .O(N__30136),
            .I(n2219));
    CascadeMux I__4638 (
            .O(N__30129),
            .I(n2217_cascade_));
    InMux I__4637 (
            .O(N__30126),
            .I(N__30123));
    LocalMux I__4636 (
            .O(N__30123),
            .I(n14598));
    InMux I__4635 (
            .O(N__30120),
            .I(N__30117));
    LocalMux I__4634 (
            .O(N__30117),
            .I(N__30114));
    Odrv4 I__4633 (
            .O(N__30114),
            .I(n2188));
    CascadeMux I__4632 (
            .O(N__30111),
            .I(N__30108));
    InMux I__4631 (
            .O(N__30108),
            .I(N__30105));
    LocalMux I__4630 (
            .O(N__30105),
            .I(N__30102));
    Odrv4 I__4629 (
            .O(N__30102),
            .I(n2300));
    CascadeMux I__4628 (
            .O(N__30099),
            .I(N__30095));
    InMux I__4627 (
            .O(N__30098),
            .I(N__30092));
    InMux I__4626 (
            .O(N__30095),
            .I(N__30089));
    LocalMux I__4625 (
            .O(N__30092),
            .I(N__30086));
    LocalMux I__4624 (
            .O(N__30089),
            .I(N__30083));
    Span4Mux_h I__4623 (
            .O(N__30086),
            .I(N__30078));
    Span4Mux_v I__4622 (
            .O(N__30083),
            .I(N__30078));
    Span4Mux_v I__4621 (
            .O(N__30078),
            .I(N__30074));
    InMux I__4620 (
            .O(N__30077),
            .I(N__30071));
    Odrv4 I__4619 (
            .O(N__30074),
            .I(n2332));
    LocalMux I__4618 (
            .O(N__30071),
            .I(n2332));
    CascadeMux I__4617 (
            .O(N__30066),
            .I(N__30063));
    InMux I__4616 (
            .O(N__30063),
            .I(N__30060));
    LocalMux I__4615 (
            .O(N__30060),
            .I(n2290));
    CascadeMux I__4614 (
            .O(N__30057),
            .I(N__30053));
    InMux I__4613 (
            .O(N__30056),
            .I(N__30050));
    InMux I__4612 (
            .O(N__30053),
            .I(N__30047));
    LocalMux I__4611 (
            .O(N__30050),
            .I(N__30041));
    LocalMux I__4610 (
            .O(N__30047),
            .I(N__30041));
    InMux I__4609 (
            .O(N__30046),
            .I(N__30038));
    Span4Mux_v I__4608 (
            .O(N__30041),
            .I(N__30033));
    LocalMux I__4607 (
            .O(N__30038),
            .I(N__30033));
    Odrv4 I__4606 (
            .O(N__30033),
            .I(n2322));
    InMux I__4605 (
            .O(N__30030),
            .I(N__30026));
    InMux I__4604 (
            .O(N__30029),
            .I(N__30023));
    LocalMux I__4603 (
            .O(N__30026),
            .I(n2116));
    LocalMux I__4602 (
            .O(N__30023),
            .I(n2116));
    CascadeMux I__4601 (
            .O(N__30018),
            .I(n2117_cascade_));
    CascadeMux I__4600 (
            .O(N__30015),
            .I(n2148_cascade_));
    InMux I__4599 (
            .O(N__30012),
            .I(N__30009));
    LocalMux I__4598 (
            .O(N__30009),
            .I(N__30006));
    Odrv4 I__4597 (
            .O(N__30006),
            .I(n2197));
    InMux I__4596 (
            .O(N__30003),
            .I(N__29998));
    CascadeMux I__4595 (
            .O(N__30002),
            .I(N__29995));
    InMux I__4594 (
            .O(N__30001),
            .I(N__29992));
    LocalMux I__4593 (
            .O(N__29998),
            .I(N__29989));
    InMux I__4592 (
            .O(N__29995),
            .I(N__29986));
    LocalMux I__4591 (
            .O(N__29992),
            .I(N__29983));
    Odrv12 I__4590 (
            .O(N__29989),
            .I(n2229));
    LocalMux I__4589 (
            .O(N__29986),
            .I(n2229));
    Odrv4 I__4588 (
            .O(N__29983),
            .I(n2229));
    CascadeMux I__4587 (
            .O(N__29976),
            .I(N__29973));
    InMux I__4586 (
            .O(N__29973),
            .I(N__29970));
    LocalMux I__4585 (
            .O(N__29970),
            .I(N__29967));
    Odrv4 I__4584 (
            .O(N__29967),
            .I(n2189));
    InMux I__4583 (
            .O(N__29964),
            .I(N__29961));
    LocalMux I__4582 (
            .O(N__29961),
            .I(n2184));
    InMux I__4581 (
            .O(N__29958),
            .I(N__29954));
    InMux I__4580 (
            .O(N__29957),
            .I(N__29951));
    LocalMux I__4579 (
            .O(N__29954),
            .I(N__29948));
    LocalMux I__4578 (
            .O(N__29951),
            .I(N__29945));
    Odrv4 I__4577 (
            .O(N__29948),
            .I(n2117));
    Odrv4 I__4576 (
            .O(N__29945),
            .I(n2117));
    InMux I__4575 (
            .O(N__29940),
            .I(N__29936));
    InMux I__4574 (
            .O(N__29939),
            .I(N__29933));
    LocalMux I__4573 (
            .O(N__29936),
            .I(N__29930));
    LocalMux I__4572 (
            .O(N__29933),
            .I(n2216));
    Odrv4 I__4571 (
            .O(N__29930),
            .I(n2216));
    InMux I__4570 (
            .O(N__29925),
            .I(N__29920));
    InMux I__4569 (
            .O(N__29924),
            .I(N__29917));
    InMux I__4568 (
            .O(N__29923),
            .I(N__29914));
    LocalMux I__4567 (
            .O(N__29920),
            .I(N__29911));
    LocalMux I__4566 (
            .O(N__29917),
            .I(N__29906));
    LocalMux I__4565 (
            .O(N__29914),
            .I(N__29906));
    Odrv4 I__4564 (
            .O(N__29911),
            .I(n2215));
    Odrv4 I__4563 (
            .O(N__29906),
            .I(n2215));
    InMux I__4562 (
            .O(N__29901),
            .I(N__29898));
    LocalMux I__4561 (
            .O(N__29898),
            .I(N__29894));
    InMux I__4560 (
            .O(N__29897),
            .I(N__29891));
    Odrv4 I__4559 (
            .O(N__29894),
            .I(n2214));
    LocalMux I__4558 (
            .O(N__29891),
            .I(n2214));
    CascadeMux I__4557 (
            .O(N__29886),
            .I(n2216_cascade_));
    InMux I__4556 (
            .O(N__29883),
            .I(N__29880));
    LocalMux I__4555 (
            .O(N__29880),
            .I(n2298));
    CascadeMux I__4554 (
            .O(N__29877),
            .I(n2247_cascade_));
    CascadeMux I__4553 (
            .O(N__29874),
            .I(N__29869));
    InMux I__4552 (
            .O(N__29873),
            .I(N__29866));
    InMux I__4551 (
            .O(N__29872),
            .I(N__29863));
    InMux I__4550 (
            .O(N__29869),
            .I(N__29860));
    LocalMux I__4549 (
            .O(N__29866),
            .I(N__29857));
    LocalMux I__4548 (
            .O(N__29863),
            .I(N__29854));
    LocalMux I__4547 (
            .O(N__29860),
            .I(N__29851));
    Span4Mux_v I__4546 (
            .O(N__29857),
            .I(N__29848));
    Span4Mux_h I__4545 (
            .O(N__29854),
            .I(N__29843));
    Span4Mux_v I__4544 (
            .O(N__29851),
            .I(N__29843));
    Odrv4 I__4543 (
            .O(N__29848),
            .I(n2330));
    Odrv4 I__4542 (
            .O(N__29843),
            .I(n2330));
    InMux I__4541 (
            .O(N__29838),
            .I(N__29835));
    LocalMux I__4540 (
            .O(N__29835),
            .I(n2193));
    CascadeMux I__4539 (
            .O(N__29832),
            .I(n2126_cascade_));
    InMux I__4538 (
            .O(N__29829),
            .I(N__29826));
    LocalMux I__4537 (
            .O(N__29826),
            .I(N__29823));
    Odrv4 I__4536 (
            .O(N__29823),
            .I(n2292));
    CascadeMux I__4535 (
            .O(N__29820),
            .I(n2225_cascade_));
    CascadeMux I__4534 (
            .O(N__29817),
            .I(N__29812));
    CascadeMux I__4533 (
            .O(N__29816),
            .I(N__29809));
    InMux I__4532 (
            .O(N__29815),
            .I(N__29806));
    InMux I__4531 (
            .O(N__29812),
            .I(N__29803));
    InMux I__4530 (
            .O(N__29809),
            .I(N__29800));
    LocalMux I__4529 (
            .O(N__29806),
            .I(N__29797));
    LocalMux I__4528 (
            .O(N__29803),
            .I(N__29794));
    LocalMux I__4527 (
            .O(N__29800),
            .I(N__29791));
    Span4Mux_h I__4526 (
            .O(N__29797),
            .I(N__29788));
    Odrv4 I__4525 (
            .O(N__29794),
            .I(n2324));
    Odrv4 I__4524 (
            .O(N__29791),
            .I(n2324));
    Odrv4 I__4523 (
            .O(N__29788),
            .I(n2324));
    CascadeMux I__4522 (
            .O(N__29781),
            .I(n2116_cascade_));
    InMux I__4521 (
            .O(N__29778),
            .I(N__29775));
    LocalMux I__4520 (
            .O(N__29775),
            .I(N__29772));
    Odrv4 I__4519 (
            .O(N__29772),
            .I(n2183));
    CascadeMux I__4518 (
            .O(N__29769),
            .I(n2049_cascade_));
    CascadeMux I__4517 (
            .O(N__29766),
            .I(N__29763));
    InMux I__4516 (
            .O(N__29763),
            .I(N__29760));
    LocalMux I__4515 (
            .O(N__29760),
            .I(n2186));
    InMux I__4514 (
            .O(N__29757),
            .I(N__29754));
    LocalMux I__4513 (
            .O(N__29754),
            .I(N__29749));
    InMux I__4512 (
            .O(N__29753),
            .I(N__29746));
    InMux I__4511 (
            .O(N__29752),
            .I(N__29743));
    Odrv4 I__4510 (
            .O(N__29749),
            .I(n3010));
    LocalMux I__4509 (
            .O(N__29746),
            .I(n3010));
    LocalMux I__4508 (
            .O(N__29743),
            .I(n3010));
    CascadeMux I__4507 (
            .O(N__29736),
            .I(N__29733));
    InMux I__4506 (
            .O(N__29733),
            .I(N__29730));
    LocalMux I__4505 (
            .O(N__29730),
            .I(N__29727));
    Odrv4 I__4504 (
            .O(N__29727),
            .I(n3077));
    CascadeMux I__4503 (
            .O(N__29724),
            .I(N__29721));
    InMux I__4502 (
            .O(N__29721),
            .I(N__29718));
    LocalMux I__4501 (
            .O(N__29718),
            .I(n2192));
    InMux I__4500 (
            .O(N__29715),
            .I(N__29712));
    LocalMux I__4499 (
            .O(N__29712),
            .I(N__29709));
    Odrv4 I__4498 (
            .O(N__29709),
            .I(n2291));
    CascadeMux I__4497 (
            .O(N__29706),
            .I(n2224_cascade_));
    InMux I__4496 (
            .O(N__29703),
            .I(N__29698));
    CascadeMux I__4495 (
            .O(N__29702),
            .I(N__29695));
    InMux I__4494 (
            .O(N__29701),
            .I(N__29692));
    LocalMux I__4493 (
            .O(N__29698),
            .I(N__29689));
    InMux I__4492 (
            .O(N__29695),
            .I(N__29686));
    LocalMux I__4491 (
            .O(N__29692),
            .I(N__29683));
    Span4Mux_s2_h I__4490 (
            .O(N__29689),
            .I(N__29676));
    LocalMux I__4489 (
            .O(N__29686),
            .I(N__29676));
    Span4Mux_v I__4488 (
            .O(N__29683),
            .I(N__29676));
    Odrv4 I__4487 (
            .O(N__29676),
            .I(n2323));
    InMux I__4486 (
            .O(N__29673),
            .I(N__29670));
    LocalMux I__4485 (
            .O(N__29670),
            .I(N__29667));
    Span4Mux_h I__4484 (
            .O(N__29667),
            .I(N__29662));
    InMux I__4483 (
            .O(N__29666),
            .I(N__29659));
    InMux I__4482 (
            .O(N__29665),
            .I(N__29656));
    Odrv4 I__4481 (
            .O(N__29662),
            .I(n3009));
    LocalMux I__4480 (
            .O(N__29659),
            .I(n3009));
    LocalMux I__4479 (
            .O(N__29656),
            .I(n3009));
    InMux I__4478 (
            .O(N__29649),
            .I(N__29645));
    InMux I__4477 (
            .O(N__29648),
            .I(N__29642));
    LocalMux I__4476 (
            .O(N__29645),
            .I(n3007));
    LocalMux I__4475 (
            .O(N__29642),
            .I(n3007));
    CascadeMux I__4474 (
            .O(N__29637),
            .I(N__29634));
    InMux I__4473 (
            .O(N__29634),
            .I(N__29630));
    InMux I__4472 (
            .O(N__29633),
            .I(N__29627));
    LocalMux I__4471 (
            .O(N__29630),
            .I(N__29624));
    LocalMux I__4470 (
            .O(N__29627),
            .I(N__29620));
    Span4Mux_h I__4469 (
            .O(N__29624),
            .I(N__29617));
    InMux I__4468 (
            .O(N__29623),
            .I(N__29614));
    Span4Mux_h I__4467 (
            .O(N__29620),
            .I(N__29611));
    Odrv4 I__4466 (
            .O(N__29617),
            .I(n3008));
    LocalMux I__4465 (
            .O(N__29614),
            .I(n3008));
    Odrv4 I__4464 (
            .O(N__29611),
            .I(n3008));
    CascadeMux I__4463 (
            .O(N__29604),
            .I(n14754_cascade_));
    InMux I__4462 (
            .O(N__29601),
            .I(N__29598));
    LocalMux I__4461 (
            .O(N__29598),
            .I(N__29594));
    InMux I__4460 (
            .O(N__29597),
            .I(N__29591));
    Span4Mux_h I__4459 (
            .O(N__29594),
            .I(N__29588));
    LocalMux I__4458 (
            .O(N__29591),
            .I(n3006));
    Odrv4 I__4457 (
            .O(N__29588),
            .I(n3006));
    InMux I__4456 (
            .O(N__29583),
            .I(N__29580));
    LocalMux I__4455 (
            .O(N__29580),
            .I(N__29577));
    Odrv4 I__4454 (
            .O(N__29577),
            .I(n3079));
    CascadeMux I__4453 (
            .O(N__29574),
            .I(n3039_cascade_));
    CascadeMux I__4452 (
            .O(N__29571),
            .I(N__29566));
    InMux I__4451 (
            .O(N__29570),
            .I(N__29563));
    InMux I__4450 (
            .O(N__29569),
            .I(N__29558));
    InMux I__4449 (
            .O(N__29566),
            .I(N__29558));
    LocalMux I__4448 (
            .O(N__29563),
            .I(n3012));
    LocalMux I__4447 (
            .O(N__29558),
            .I(n3012));
    CascadeMux I__4446 (
            .O(N__29553),
            .I(n14194_cascade_));
    InMux I__4445 (
            .O(N__29550),
            .I(N__29547));
    LocalMux I__4444 (
            .O(N__29547),
            .I(n14196));
    InMux I__4443 (
            .O(N__29544),
            .I(N__29541));
    LocalMux I__4442 (
            .O(N__29541),
            .I(N__29537));
    InMux I__4441 (
            .O(N__29540),
            .I(N__29534));
    Odrv4 I__4440 (
            .O(N__29537),
            .I(n3018));
    LocalMux I__4439 (
            .O(N__29534),
            .I(n3018));
    InMux I__4438 (
            .O(N__29529),
            .I(N__29526));
    LocalMux I__4437 (
            .O(N__29526),
            .I(N__29523));
    Span4Mux_s1_v I__4436 (
            .O(N__29523),
            .I(N__29520));
    Odrv4 I__4435 (
            .O(N__29520),
            .I(n3085));
    CascadeMux I__4434 (
            .O(N__29517),
            .I(n3117_cascade_));
    InMux I__4433 (
            .O(N__29514),
            .I(N__29511));
    LocalMux I__4432 (
            .O(N__29511),
            .I(n14198));
    InMux I__4431 (
            .O(N__29508),
            .I(N__29505));
    LocalMux I__4430 (
            .O(N__29505),
            .I(N__29500));
    InMux I__4429 (
            .O(N__29504),
            .I(N__29497));
    InMux I__4428 (
            .O(N__29503),
            .I(N__29494));
    Odrv4 I__4427 (
            .O(N__29500),
            .I(n3017));
    LocalMux I__4426 (
            .O(N__29497),
            .I(n3017));
    LocalMux I__4425 (
            .O(N__29494),
            .I(n3017));
    InMux I__4424 (
            .O(N__29487),
            .I(N__29484));
    LocalMux I__4423 (
            .O(N__29484),
            .I(N__29481));
    Span4Mux_s1_v I__4422 (
            .O(N__29481),
            .I(N__29478));
    Odrv4 I__4421 (
            .O(N__29478),
            .I(n3084));
    CascadeMux I__4420 (
            .O(N__29475),
            .I(N__29471));
    InMux I__4419 (
            .O(N__29474),
            .I(N__29468));
    InMux I__4418 (
            .O(N__29471),
            .I(N__29465));
    LocalMux I__4417 (
            .O(N__29468),
            .I(N__29462));
    LocalMux I__4416 (
            .O(N__29465),
            .I(N__29459));
    Span4Mux_s2_v I__4415 (
            .O(N__29462),
            .I(N__29454));
    Span4Mux_h I__4414 (
            .O(N__29459),
            .I(N__29454));
    Odrv4 I__4413 (
            .O(N__29454),
            .I(n3025));
    CascadeMux I__4412 (
            .O(N__29451),
            .I(N__29448));
    InMux I__4411 (
            .O(N__29448),
            .I(N__29445));
    LocalMux I__4410 (
            .O(N__29445),
            .I(N__29442));
    Span4Mux_s2_v I__4409 (
            .O(N__29442),
            .I(N__29439));
    Odrv4 I__4408 (
            .O(N__29439),
            .I(n3092));
    InMux I__4407 (
            .O(N__29436),
            .I(N__29433));
    LocalMux I__4406 (
            .O(N__29433),
            .I(N__29430));
    Span4Mux_h I__4405 (
            .O(N__29430),
            .I(N__29427));
    Odrv4 I__4404 (
            .O(N__29427),
            .I(n2999));
    CascadeMux I__4403 (
            .O(N__29424),
            .I(N__29421));
    InMux I__4402 (
            .O(N__29421),
            .I(N__29418));
    LocalMux I__4401 (
            .O(N__29418),
            .I(N__29414));
    CascadeMux I__4400 (
            .O(N__29417),
            .I(N__29411));
    Span4Mux_h I__4399 (
            .O(N__29414),
            .I(N__29408));
    InMux I__4398 (
            .O(N__29411),
            .I(N__29405));
    Odrv4 I__4397 (
            .O(N__29408),
            .I(n2932));
    LocalMux I__4396 (
            .O(N__29405),
            .I(n2932));
    CascadeMux I__4395 (
            .O(N__29400),
            .I(N__29397));
    InMux I__4394 (
            .O(N__29397),
            .I(N__29393));
    CascadeMux I__4393 (
            .O(N__29396),
            .I(N__29390));
    LocalMux I__4392 (
            .O(N__29393),
            .I(N__29387));
    InMux I__4391 (
            .O(N__29390),
            .I(N__29384));
    Span4Mux_v I__4390 (
            .O(N__29387),
            .I(N__29381));
    LocalMux I__4389 (
            .O(N__29384),
            .I(n3031));
    Odrv4 I__4388 (
            .O(N__29381),
            .I(n3031));
    InMux I__4387 (
            .O(N__29376),
            .I(N__29373));
    LocalMux I__4386 (
            .O(N__29373),
            .I(N__29370));
    Span4Mux_s3_v I__4385 (
            .O(N__29370),
            .I(N__29367));
    Odrv4 I__4384 (
            .O(N__29367),
            .I(n3098));
    CascadeMux I__4383 (
            .O(N__29364),
            .I(n3031_cascade_));
    InMux I__4382 (
            .O(N__29361),
            .I(N__29357));
    InMux I__4381 (
            .O(N__29360),
            .I(N__29353));
    LocalMux I__4380 (
            .O(N__29357),
            .I(N__29350));
    InMux I__4379 (
            .O(N__29356),
            .I(N__29347));
    LocalMux I__4378 (
            .O(N__29353),
            .I(N__29344));
    Span4Mux_h I__4377 (
            .O(N__29350),
            .I(N__29341));
    LocalMux I__4376 (
            .O(N__29347),
            .I(N__29338));
    Span4Mux_v I__4375 (
            .O(N__29344),
            .I(N__29335));
    Odrv4 I__4374 (
            .O(N__29341),
            .I(n2916));
    Odrv12 I__4373 (
            .O(N__29338),
            .I(n2916));
    Odrv4 I__4372 (
            .O(N__29335),
            .I(n2916));
    CascadeMux I__4371 (
            .O(N__29328),
            .I(N__29325));
    InMux I__4370 (
            .O(N__29325),
            .I(N__29322));
    LocalMux I__4369 (
            .O(N__29322),
            .I(N__29319));
    Span4Mux_h I__4368 (
            .O(N__29319),
            .I(N__29316));
    Odrv4 I__4367 (
            .O(N__29316),
            .I(n2983));
    InMux I__4366 (
            .O(N__29313),
            .I(N__29310));
    LocalMux I__4365 (
            .O(N__29310),
            .I(N__29307));
    Span4Mux_s2_v I__4364 (
            .O(N__29307),
            .I(N__29303));
    InMux I__4363 (
            .O(N__29306),
            .I(N__29300));
    Odrv4 I__4362 (
            .O(N__29303),
            .I(n3015));
    LocalMux I__4361 (
            .O(N__29300),
            .I(n3015));
    InMux I__4360 (
            .O(N__29295),
            .I(N__29292));
    LocalMux I__4359 (
            .O(N__29292),
            .I(N__29289));
    Span4Mux_h I__4358 (
            .O(N__29289),
            .I(N__29286));
    Odrv4 I__4357 (
            .O(N__29286),
            .I(n3082));
    CascadeMux I__4356 (
            .O(N__29283),
            .I(n3015_cascade_));
    InMux I__4355 (
            .O(N__29280),
            .I(N__29277));
    LocalMux I__4354 (
            .O(N__29277),
            .I(N__29274));
    Span4Mux_s2_v I__4353 (
            .O(N__29274),
            .I(N__29271));
    Odrv4 I__4352 (
            .O(N__29271),
            .I(n3089));
    CascadeMux I__4351 (
            .O(N__29268),
            .I(N__29265));
    InMux I__4350 (
            .O(N__29265),
            .I(N__29261));
    InMux I__4349 (
            .O(N__29264),
            .I(N__29258));
    LocalMux I__4348 (
            .O(N__29261),
            .I(N__29255));
    LocalMux I__4347 (
            .O(N__29258),
            .I(N__29252));
    Odrv4 I__4346 (
            .O(N__29255),
            .I(n3022));
    Odrv4 I__4345 (
            .O(N__29252),
            .I(n3022));
    InMux I__4344 (
            .O(N__29247),
            .I(N__29244));
    LocalMux I__4343 (
            .O(N__29244),
            .I(N__29241));
    Span4Mux_h I__4342 (
            .O(N__29241),
            .I(N__29238));
    Odrv4 I__4341 (
            .O(N__29238),
            .I(n3095));
    CascadeMux I__4340 (
            .O(N__29235),
            .I(N__29230));
    InMux I__4339 (
            .O(N__29234),
            .I(N__29227));
    InMux I__4338 (
            .O(N__29233),
            .I(N__29224));
    InMux I__4337 (
            .O(N__29230),
            .I(N__29221));
    LocalMux I__4336 (
            .O(N__29227),
            .I(N__29216));
    LocalMux I__4335 (
            .O(N__29224),
            .I(N__29216));
    LocalMux I__4334 (
            .O(N__29221),
            .I(n3028));
    Odrv4 I__4333 (
            .O(N__29216),
            .I(n3028));
    CascadeMux I__4332 (
            .O(N__29211),
            .I(n3127_cascade_));
    InMux I__4331 (
            .O(N__29208),
            .I(N__29203));
    InMux I__4330 (
            .O(N__29207),
            .I(N__29200));
    InMux I__4329 (
            .O(N__29206),
            .I(N__29197));
    LocalMux I__4328 (
            .O(N__29203),
            .I(n3011));
    LocalMux I__4327 (
            .O(N__29200),
            .I(n3011));
    LocalMux I__4326 (
            .O(N__29197),
            .I(n3011));
    InMux I__4325 (
            .O(N__29190),
            .I(N__29187));
    LocalMux I__4324 (
            .O(N__29187),
            .I(n14744));
    InMux I__4323 (
            .O(N__29184),
            .I(N__29181));
    LocalMux I__4322 (
            .O(N__29181),
            .I(n14816));
    CascadeMux I__4321 (
            .O(N__29178),
            .I(n14750_cascade_));
    InMux I__4320 (
            .O(N__29175),
            .I(N__29172));
    LocalMux I__4319 (
            .O(N__29172),
            .I(N__29167));
    InMux I__4318 (
            .O(N__29171),
            .I(N__29164));
    InMux I__4317 (
            .O(N__29170),
            .I(N__29161));
    Odrv4 I__4316 (
            .O(N__29167),
            .I(n3014));
    LocalMux I__4315 (
            .O(N__29164),
            .I(n3014));
    LocalMux I__4314 (
            .O(N__29161),
            .I(n3014));
    CascadeMux I__4313 (
            .O(N__29154),
            .I(N__29151));
    InMux I__4312 (
            .O(N__29151),
            .I(N__29148));
    LocalMux I__4311 (
            .O(N__29148),
            .I(N__29145));
    Span4Mux_v I__4310 (
            .O(N__29145),
            .I(N__29142));
    Odrv4 I__4309 (
            .O(N__29142),
            .I(n3081));
    InMux I__4308 (
            .O(N__29139),
            .I(N__29136));
    LocalMux I__4307 (
            .O(N__29136),
            .I(N__29133));
    Odrv4 I__4306 (
            .O(N__29133),
            .I(n3100));
    CascadeMux I__4305 (
            .O(N__29130),
            .I(N__29127));
    InMux I__4304 (
            .O(N__29127),
            .I(N__29124));
    LocalMux I__4303 (
            .O(N__29124),
            .I(N__29121));
    Odrv4 I__4302 (
            .O(N__29121),
            .I(n3001));
    CascadeMux I__4301 (
            .O(N__29118),
            .I(N__29115));
    InMux I__4300 (
            .O(N__29115),
            .I(N__29111));
    InMux I__4299 (
            .O(N__29114),
            .I(N__29108));
    LocalMux I__4298 (
            .O(N__29111),
            .I(N__29105));
    LocalMux I__4297 (
            .O(N__29108),
            .I(n3033));
    Odrv4 I__4296 (
            .O(N__29105),
            .I(n3033));
    CascadeMux I__4295 (
            .O(N__29100),
            .I(n3033_cascade_));
    CascadeMux I__4294 (
            .O(N__29097),
            .I(N__29094));
    InMux I__4293 (
            .O(N__29094),
            .I(N__29089));
    InMux I__4292 (
            .O(N__29093),
            .I(N__29084));
    InMux I__4291 (
            .O(N__29092),
            .I(N__29084));
    LocalMux I__4290 (
            .O(N__29089),
            .I(N__29079));
    LocalMux I__4289 (
            .O(N__29084),
            .I(N__29079));
    Span4Mux_h I__4288 (
            .O(N__29079),
            .I(N__29076));
    Odrv4 I__4287 (
            .O(N__29076),
            .I(n3032));
    CascadeMux I__4286 (
            .O(N__29073),
            .I(N__29070));
    InMux I__4285 (
            .O(N__29070),
            .I(N__29067));
    LocalMux I__4284 (
            .O(N__29067),
            .I(N__29064));
    Odrv4 I__4283 (
            .O(N__29064),
            .I(n2990));
    CascadeMux I__4282 (
            .O(N__29061),
            .I(n3022_cascade_));
    InMux I__4281 (
            .O(N__29058),
            .I(N__29055));
    LocalMux I__4280 (
            .O(N__29055),
            .I(n14732));
    CascadeMux I__4279 (
            .O(N__29052),
            .I(N__29049));
    InMux I__4278 (
            .O(N__29049),
            .I(N__29045));
    InMux I__4277 (
            .O(N__29048),
            .I(N__29042));
    LocalMux I__4276 (
            .O(N__29045),
            .I(n3030));
    LocalMux I__4275 (
            .O(N__29042),
            .I(n3030));
    CascadeMux I__4274 (
            .O(N__29037),
            .I(N__29034));
    InMux I__4273 (
            .O(N__29034),
            .I(N__29030));
    InMux I__4272 (
            .O(N__29033),
            .I(N__29027));
    LocalMux I__4271 (
            .O(N__29030),
            .I(n3029));
    LocalMux I__4270 (
            .O(N__29027),
            .I(n3029));
    InMux I__4269 (
            .O(N__29022),
            .I(N__29019));
    LocalMux I__4268 (
            .O(N__29019),
            .I(n11932));
    CascadeMux I__4267 (
            .O(N__29016),
            .I(n13859_cascade_));
    InMux I__4266 (
            .O(N__29013),
            .I(N__29010));
    LocalMux I__4265 (
            .O(N__29010),
            .I(n14738));
    InMux I__4264 (
            .O(N__29007),
            .I(n12904));
    InMux I__4263 (
            .O(N__29004),
            .I(n12905));
    InMux I__4262 (
            .O(N__29001),
            .I(n12906));
    CascadeMux I__4261 (
            .O(N__28998),
            .I(N__28995));
    InMux I__4260 (
            .O(N__28995),
            .I(N__28992));
    LocalMux I__4259 (
            .O(N__28992),
            .I(N__28989));
    Odrv4 I__4258 (
            .O(N__28989),
            .I(n3180));
    CascadeMux I__4257 (
            .O(N__28986),
            .I(N__28982));
    InMux I__4256 (
            .O(N__28985),
            .I(N__28979));
    InMux I__4255 (
            .O(N__28982),
            .I(N__28976));
    LocalMux I__4254 (
            .O(N__28979),
            .I(N__28972));
    LocalMux I__4253 (
            .O(N__28976),
            .I(N__28969));
    InMux I__4252 (
            .O(N__28975),
            .I(N__28966));
    Odrv4 I__4251 (
            .O(N__28972),
            .I(n2925));
    Odrv4 I__4250 (
            .O(N__28969),
            .I(n2925));
    LocalMux I__4249 (
            .O(N__28966),
            .I(n2925));
    CascadeMux I__4248 (
            .O(N__28959),
            .I(N__28956));
    InMux I__4247 (
            .O(N__28956),
            .I(N__28953));
    LocalMux I__4246 (
            .O(N__28953),
            .I(N__28950));
    Span4Mux_h I__4245 (
            .O(N__28950),
            .I(N__28947));
    Odrv4 I__4244 (
            .O(N__28947),
            .I(n2992));
    CascadeMux I__4243 (
            .O(N__28944),
            .I(N__28941));
    InMux I__4242 (
            .O(N__28941),
            .I(N__28938));
    LocalMux I__4241 (
            .O(N__28938),
            .I(N__28935));
    Odrv4 I__4240 (
            .O(N__28935),
            .I(n3099));
    CascadeMux I__4239 (
            .O(N__28932),
            .I(N__28929));
    InMux I__4238 (
            .O(N__28929),
            .I(N__28926));
    LocalMux I__4237 (
            .O(N__28926),
            .I(N__28923));
    Span4Mux_v I__4236 (
            .O(N__28923),
            .I(N__28920));
    Odrv4 I__4235 (
            .O(N__28920),
            .I(n3076));
    CascadeMux I__4234 (
            .O(N__28917),
            .I(N__28914));
    InMux I__4233 (
            .O(N__28914),
            .I(N__28910));
    InMux I__4232 (
            .O(N__28913),
            .I(N__28907));
    LocalMux I__4231 (
            .O(N__28910),
            .I(N__28904));
    LocalMux I__4230 (
            .O(N__28907),
            .I(N__28901));
    Span4Mux_s3_h I__4229 (
            .O(N__28904),
            .I(N__28898));
    Odrv4 I__4228 (
            .O(N__28901),
            .I(n2926));
    Odrv4 I__4227 (
            .O(N__28898),
            .I(n2926));
    CascadeMux I__4226 (
            .O(N__28893),
            .I(N__28890));
    InMux I__4225 (
            .O(N__28890),
            .I(N__28887));
    LocalMux I__4224 (
            .O(N__28887),
            .I(N__28884));
    Span4Mux_v I__4223 (
            .O(N__28884),
            .I(N__28881));
    Odrv4 I__4222 (
            .O(N__28881),
            .I(n2993));
    InMux I__4221 (
            .O(N__28878),
            .I(N__28874));
    CascadeMux I__4220 (
            .O(N__28877),
            .I(N__28871));
    LocalMux I__4219 (
            .O(N__28874),
            .I(N__28867));
    InMux I__4218 (
            .O(N__28871),
            .I(N__28864));
    InMux I__4217 (
            .O(N__28870),
            .I(N__28861));
    Odrv4 I__4216 (
            .O(N__28867),
            .I(n3027));
    LocalMux I__4215 (
            .O(N__28864),
            .I(n3027));
    LocalMux I__4214 (
            .O(N__28861),
            .I(n3027));
    CascadeMux I__4213 (
            .O(N__28854),
            .I(n3025_cascade_));
    InMux I__4212 (
            .O(N__28851),
            .I(N__28848));
    LocalMux I__4211 (
            .O(N__28848),
            .I(n14736));
    InMux I__4210 (
            .O(N__28845),
            .I(n12895));
    InMux I__4209 (
            .O(N__28842),
            .I(n12896));
    InMux I__4208 (
            .O(N__28839),
            .I(n12897));
    InMux I__4207 (
            .O(N__28836),
            .I(n12898));
    InMux I__4206 (
            .O(N__28833),
            .I(n12899));
    InMux I__4205 (
            .O(N__28830),
            .I(n12900));
    InMux I__4204 (
            .O(N__28827),
            .I(bfn_5_28_0_));
    InMux I__4203 (
            .O(N__28824),
            .I(n12902));
    InMux I__4202 (
            .O(N__28821),
            .I(n12903));
    InMux I__4201 (
            .O(N__28818),
            .I(n12886));
    InMux I__4200 (
            .O(N__28815),
            .I(n12887));
    InMux I__4199 (
            .O(N__28812),
            .I(n12888));
    InMux I__4198 (
            .O(N__28809),
            .I(n12889));
    InMux I__4197 (
            .O(N__28806),
            .I(n12890));
    InMux I__4196 (
            .O(N__28803),
            .I(n12891));
    InMux I__4195 (
            .O(N__28800),
            .I(n12892));
    InMux I__4194 (
            .O(N__28797),
            .I(bfn_5_27_0_));
    InMux I__4193 (
            .O(N__28794),
            .I(n12894));
    InMux I__4192 (
            .O(N__28791),
            .I(bfn_5_25_0_));
    InMux I__4191 (
            .O(N__28788),
            .I(n12878));
    InMux I__4190 (
            .O(N__28785),
            .I(n12879));
    InMux I__4189 (
            .O(N__28782),
            .I(n12880));
    InMux I__4188 (
            .O(N__28779),
            .I(n12881));
    InMux I__4187 (
            .O(N__28776),
            .I(n12882));
    InMux I__4186 (
            .O(N__28773),
            .I(n12883));
    InMux I__4185 (
            .O(N__28770),
            .I(n12884));
    InMux I__4184 (
            .O(N__28767),
            .I(bfn_5_26_0_));
    InMux I__4183 (
            .O(N__28764),
            .I(N__28761));
    LocalMux I__4182 (
            .O(N__28761),
            .I(N__28758));
    Odrv4 I__4181 (
            .O(N__28758),
            .I(n2289));
    CascadeMux I__4180 (
            .O(N__28755),
            .I(N__28751));
    CascadeMux I__4179 (
            .O(N__28754),
            .I(N__28748));
    InMux I__4178 (
            .O(N__28751),
            .I(N__28745));
    InMux I__4177 (
            .O(N__28748),
            .I(N__28741));
    LocalMux I__4176 (
            .O(N__28745),
            .I(N__28738));
    InMux I__4175 (
            .O(N__28744),
            .I(N__28735));
    LocalMux I__4174 (
            .O(N__28741),
            .I(N__28732));
    Span4Mux_v I__4173 (
            .O(N__28738),
            .I(N__28729));
    LocalMux I__4172 (
            .O(N__28735),
            .I(N__28726));
    Span4Mux_v I__4171 (
            .O(N__28732),
            .I(N__28723));
    Span4Mux_v I__4170 (
            .O(N__28729),
            .I(N__28718));
    Span4Mux_v I__4169 (
            .O(N__28726),
            .I(N__28718));
    Odrv4 I__4168 (
            .O(N__28723),
            .I(n2321));
    Odrv4 I__4167 (
            .O(N__28718),
            .I(n2321));
    InMux I__4166 (
            .O(N__28713),
            .I(N__28709));
    InMux I__4165 (
            .O(N__28712),
            .I(N__28706));
    LocalMux I__4164 (
            .O(N__28709),
            .I(N__28702));
    LocalMux I__4163 (
            .O(N__28706),
            .I(N__28699));
    CascadeMux I__4162 (
            .O(N__28705),
            .I(N__28696));
    Span4Mux_h I__4161 (
            .O(N__28702),
            .I(N__28691));
    Span4Mux_v I__4160 (
            .O(N__28699),
            .I(N__28691));
    InMux I__4159 (
            .O(N__28696),
            .I(N__28688));
    Odrv4 I__4158 (
            .O(N__28691),
            .I(n2331));
    LocalMux I__4157 (
            .O(N__28688),
            .I(n2331));
    InMux I__4156 (
            .O(N__28683),
            .I(N__28680));
    LocalMux I__4155 (
            .O(N__28680),
            .I(N__28677));
    Span4Mux_h I__4154 (
            .O(N__28677),
            .I(N__28674));
    Odrv4 I__4153 (
            .O(N__28674),
            .I(n11954));
    InMux I__4152 (
            .O(N__28671),
            .I(N__28666));
    InMux I__4151 (
            .O(N__28670),
            .I(N__28663));
    InMux I__4150 (
            .O(N__28669),
            .I(N__28660));
    LocalMux I__4149 (
            .O(N__28666),
            .I(N__28655));
    LocalMux I__4148 (
            .O(N__28663),
            .I(N__28655));
    LocalMux I__4147 (
            .O(N__28660),
            .I(N__28652));
    Span4Mux_v I__4146 (
            .O(N__28655),
            .I(N__28649));
    Span4Mux_h I__4145 (
            .O(N__28652),
            .I(N__28646));
    Span4Mux_h I__4144 (
            .O(N__28649),
            .I(N__28643));
    Odrv4 I__4143 (
            .O(N__28646),
            .I(n311));
    Odrv4 I__4142 (
            .O(N__28643),
            .I(n311));
    InMux I__4141 (
            .O(N__28638),
            .I(N__28634));
    CascadeMux I__4140 (
            .O(N__28637),
            .I(N__28631));
    LocalMux I__4139 (
            .O(N__28634),
            .I(N__28628));
    InMux I__4138 (
            .O(N__28631),
            .I(N__28625));
    Span4Mux_v I__4137 (
            .O(N__28628),
            .I(N__28622));
    LocalMux I__4136 (
            .O(N__28625),
            .I(N__28619));
    Span4Mux_v I__4135 (
            .O(N__28622),
            .I(N__28613));
    Span4Mux_v I__4134 (
            .O(N__28619),
            .I(N__28613));
    InMux I__4133 (
            .O(N__28618),
            .I(N__28610));
    Odrv4 I__4132 (
            .O(N__28613),
            .I(n2533));
    LocalMux I__4131 (
            .O(N__28610),
            .I(n2533));
    CascadeMux I__4130 (
            .O(N__28605),
            .I(N__28602));
    InMux I__4129 (
            .O(N__28602),
            .I(N__28599));
    LocalMux I__4128 (
            .O(N__28599),
            .I(N__28596));
    Span4Mux_v I__4127 (
            .O(N__28596),
            .I(N__28593));
    Odrv4 I__4126 (
            .O(N__28593),
            .I(n2600));
    InMux I__4125 (
            .O(N__28590),
            .I(N__28587));
    LocalMux I__4124 (
            .O(N__28587),
            .I(N__28583));
    CascadeMux I__4123 (
            .O(N__28586),
            .I(N__28580));
    Span4Mux_h I__4122 (
            .O(N__28583),
            .I(N__28577));
    InMux I__4121 (
            .O(N__28580),
            .I(N__28574));
    Span4Mux_v I__4120 (
            .O(N__28577),
            .I(N__28569));
    LocalMux I__4119 (
            .O(N__28574),
            .I(N__28569));
    Odrv4 I__4118 (
            .O(N__28569),
            .I(n2532));
    CascadeMux I__4117 (
            .O(N__28566),
            .I(N__28563));
    InMux I__4116 (
            .O(N__28563),
            .I(N__28560));
    LocalMux I__4115 (
            .O(N__28560),
            .I(N__28557));
    Span4Mux_v I__4114 (
            .O(N__28557),
            .I(N__28554));
    Odrv4 I__4113 (
            .O(N__28554),
            .I(n2599));
    InMux I__4112 (
            .O(N__28551),
            .I(N__28547));
    InMux I__4111 (
            .O(N__28550),
            .I(N__28544));
    LocalMux I__4110 (
            .O(N__28547),
            .I(N__28541));
    LocalMux I__4109 (
            .O(N__28544),
            .I(n2631));
    Odrv4 I__4108 (
            .O(N__28541),
            .I(n2631));
    InMux I__4107 (
            .O(N__28536),
            .I(N__28531));
    CascadeMux I__4106 (
            .O(N__28535),
            .I(N__28528));
    CascadeMux I__4105 (
            .O(N__28534),
            .I(N__28525));
    LocalMux I__4104 (
            .O(N__28531),
            .I(N__28522));
    InMux I__4103 (
            .O(N__28528),
            .I(N__28519));
    InMux I__4102 (
            .O(N__28525),
            .I(N__28516));
    Span4Mux_v I__4101 (
            .O(N__28522),
            .I(N__28513));
    LocalMux I__4100 (
            .O(N__28519),
            .I(n2633));
    LocalMux I__4099 (
            .O(N__28516),
            .I(n2633));
    Odrv4 I__4098 (
            .O(N__28513),
            .I(n2633));
    CascadeMux I__4097 (
            .O(N__28506),
            .I(n2631_cascade_));
    InMux I__4096 (
            .O(N__28503),
            .I(N__28499));
    InMux I__4095 (
            .O(N__28502),
            .I(N__28495));
    LocalMux I__4094 (
            .O(N__28499),
            .I(N__28492));
    InMux I__4093 (
            .O(N__28498),
            .I(N__28489));
    LocalMux I__4092 (
            .O(N__28495),
            .I(n2632));
    Odrv4 I__4091 (
            .O(N__28492),
            .I(n2632));
    LocalMux I__4090 (
            .O(N__28489),
            .I(n2632));
    InMux I__4089 (
            .O(N__28482),
            .I(N__28479));
    LocalMux I__4088 (
            .O(N__28479),
            .I(N__28476));
    Span4Mux_h I__4087 (
            .O(N__28476),
            .I(N__28473));
    Odrv4 I__4086 (
            .O(N__28473),
            .I(n12044));
    CascadeMux I__4085 (
            .O(N__28470),
            .I(N__28467));
    InMux I__4084 (
            .O(N__28467),
            .I(N__28464));
    LocalMux I__4083 (
            .O(N__28464),
            .I(N__28461));
    Odrv12 I__4082 (
            .O(N__28461),
            .I(n2301));
    CascadeMux I__4081 (
            .O(N__28458),
            .I(N__28455));
    InMux I__4080 (
            .O(N__28455),
            .I(N__28451));
    InMux I__4079 (
            .O(N__28454),
            .I(N__28448));
    LocalMux I__4078 (
            .O(N__28451),
            .I(N__28445));
    LocalMux I__4077 (
            .O(N__28448),
            .I(N__28442));
    Span12Mux_v I__4076 (
            .O(N__28445),
            .I(N__28438));
    Sp12to4 I__4075 (
            .O(N__28442),
            .I(N__28435));
    InMux I__4074 (
            .O(N__28441),
            .I(N__28432));
    Odrv12 I__4073 (
            .O(N__28438),
            .I(n2333));
    Odrv12 I__4072 (
            .O(N__28435),
            .I(n2333));
    LocalMux I__4071 (
            .O(N__28432),
            .I(n2333));
    InMux I__4070 (
            .O(N__28425),
            .I(bfn_5_22_0_));
    InMux I__4069 (
            .O(N__28422),
            .I(n12678));
    InMux I__4068 (
            .O(N__28419),
            .I(N__28416));
    LocalMux I__4067 (
            .O(N__28416),
            .I(N__28413));
    Odrv4 I__4066 (
            .O(N__28413),
            .I(n2283));
    InMux I__4065 (
            .O(N__28410),
            .I(n12679));
    InMux I__4064 (
            .O(N__28407),
            .I(N__28404));
    LocalMux I__4063 (
            .O(N__28404),
            .I(N__28401));
    Span4Mux_h I__4062 (
            .O(N__28401),
            .I(N__28398));
    Odrv4 I__4061 (
            .O(N__28398),
            .I(n2282));
    InMux I__4060 (
            .O(N__28395),
            .I(n12680));
    InMux I__4059 (
            .O(N__28392),
            .I(n12681));
    InMux I__4058 (
            .O(N__28389),
            .I(N__28385));
    InMux I__4057 (
            .O(N__28388),
            .I(N__28382));
    LocalMux I__4056 (
            .O(N__28385),
            .I(N__28379));
    LocalMux I__4055 (
            .O(N__28382),
            .I(N__28376));
    Span4Mux_v I__4054 (
            .O(N__28379),
            .I(N__28373));
    Odrv4 I__4053 (
            .O(N__28376),
            .I(n2313));
    Odrv4 I__4052 (
            .O(N__28373),
            .I(n2313));
    InMux I__4051 (
            .O(N__28368),
            .I(N__28365));
    LocalMux I__4050 (
            .O(N__28365),
            .I(N__28362));
    Odrv4 I__4049 (
            .O(N__28362),
            .I(n2299));
    InMux I__4048 (
            .O(N__28359),
            .I(N__28356));
    LocalMux I__4047 (
            .O(N__28356),
            .I(N__28353));
    Span4Mux_v I__4046 (
            .O(N__28353),
            .I(N__28350));
    Odrv4 I__4045 (
            .O(N__28350),
            .I(n2196));
    InMux I__4044 (
            .O(N__28347),
            .I(N__28344));
    LocalMux I__4043 (
            .O(N__28344),
            .I(N__28341));
    Odrv12 I__4042 (
            .O(N__28341),
            .I(n2198));
    InMux I__4041 (
            .O(N__28338),
            .I(N__28335));
    LocalMux I__4040 (
            .O(N__28335),
            .I(N__28331));
    InMux I__4039 (
            .O(N__28334),
            .I(N__28328));
    Span4Mux_h I__4038 (
            .O(N__28331),
            .I(N__28325));
    LocalMux I__4037 (
            .O(N__28328),
            .I(N__28322));
    Odrv4 I__4036 (
            .O(N__28325),
            .I(n2230));
    Odrv4 I__4035 (
            .O(N__28322),
            .I(n2230));
    CascadeMux I__4034 (
            .O(N__28317),
            .I(n2230_cascade_));
    InMux I__4033 (
            .O(N__28314),
            .I(n12668));
    CascadeMux I__4032 (
            .O(N__28311),
            .I(N__28308));
    InMux I__4031 (
            .O(N__28308),
            .I(N__28305));
    LocalMux I__4030 (
            .O(N__28305),
            .I(N__28302));
    Odrv4 I__4029 (
            .O(N__28302),
            .I(n2293));
    InMux I__4028 (
            .O(N__28299),
            .I(bfn_5_21_0_));
    InMux I__4027 (
            .O(N__28296),
            .I(n12670));
    InMux I__4026 (
            .O(N__28293),
            .I(n12671));
    InMux I__4025 (
            .O(N__28290),
            .I(n12672));
    InMux I__4024 (
            .O(N__28287),
            .I(n12673));
    InMux I__4023 (
            .O(N__28284),
            .I(N__28281));
    LocalMux I__4022 (
            .O(N__28281),
            .I(n2288));
    InMux I__4021 (
            .O(N__28278),
            .I(n12674));
    InMux I__4020 (
            .O(N__28275),
            .I(N__28272));
    LocalMux I__4019 (
            .O(N__28272),
            .I(n2287));
    InMux I__4018 (
            .O(N__28269),
            .I(n12675));
    InMux I__4017 (
            .O(N__28266),
            .I(N__28263));
    LocalMux I__4016 (
            .O(N__28263),
            .I(n2286));
    InMux I__4015 (
            .O(N__28260),
            .I(n12676));
    InMux I__4014 (
            .O(N__28257),
            .I(N__28254));
    LocalMux I__4013 (
            .O(N__28254),
            .I(N__28251));
    Odrv4 I__4012 (
            .O(N__28251),
            .I(n2195));
    InMux I__4011 (
            .O(N__28248),
            .I(bfn_5_20_0_));
    InMux I__4010 (
            .O(N__28245),
            .I(n12662));
    InMux I__4009 (
            .O(N__28242),
            .I(n12663));
    InMux I__4008 (
            .O(N__28239),
            .I(n12664));
    CascadeMux I__4007 (
            .O(N__28236),
            .I(N__28233));
    InMux I__4006 (
            .O(N__28233),
            .I(N__28230));
    LocalMux I__4005 (
            .O(N__28230),
            .I(N__28227));
    Odrv4 I__4004 (
            .O(N__28227),
            .I(n2297));
    InMux I__4003 (
            .O(N__28224),
            .I(n12665));
    InMux I__4002 (
            .O(N__28221),
            .I(N__28218));
    LocalMux I__4001 (
            .O(N__28218),
            .I(N__28215));
    Odrv4 I__4000 (
            .O(N__28215),
            .I(n2296));
    InMux I__3999 (
            .O(N__28212),
            .I(n12666));
    CascadeMux I__3998 (
            .O(N__28209),
            .I(N__28206));
    InMux I__3997 (
            .O(N__28206),
            .I(N__28203));
    LocalMux I__3996 (
            .O(N__28203),
            .I(n2295));
    InMux I__3995 (
            .O(N__28200),
            .I(n12667));
    CascadeMux I__3994 (
            .O(N__28197),
            .I(N__28194));
    InMux I__3993 (
            .O(N__28194),
            .I(N__28191));
    LocalMux I__3992 (
            .O(N__28191),
            .I(n2294));
    InMux I__3991 (
            .O(N__28188),
            .I(n12655));
    InMux I__3990 (
            .O(N__28185),
            .I(n12656));
    InMux I__3989 (
            .O(N__28182),
            .I(n12657));
    InMux I__3988 (
            .O(N__28179),
            .I(bfn_5_19_0_));
    InMux I__3987 (
            .O(N__28176),
            .I(n12659));
    InMux I__3986 (
            .O(N__28173),
            .I(n12660));
    InMux I__3985 (
            .O(N__28170),
            .I(n12661));
    CascadeMux I__3984 (
            .O(N__28167),
            .I(N__28163));
    CascadeMux I__3983 (
            .O(N__28166),
            .I(N__28159));
    InMux I__3982 (
            .O(N__28163),
            .I(N__28154));
    InMux I__3981 (
            .O(N__28162),
            .I(N__28154));
    InMux I__3980 (
            .O(N__28159),
            .I(N__28151));
    LocalMux I__3979 (
            .O(N__28154),
            .I(N__28148));
    LocalMux I__3978 (
            .O(N__28151),
            .I(n2315));
    Odrv4 I__3977 (
            .O(N__28148),
            .I(n2315));
    InMux I__3976 (
            .O(N__28143),
            .I(N__28140));
    LocalMux I__3975 (
            .O(N__28140),
            .I(N__28136));
    CascadeMux I__3974 (
            .O(N__28139),
            .I(N__28133));
    Span4Mux_h I__3973 (
            .O(N__28136),
            .I(N__28129));
    InMux I__3972 (
            .O(N__28133),
            .I(N__28126));
    InMux I__3971 (
            .O(N__28132),
            .I(N__28123));
    Odrv4 I__3970 (
            .O(N__28129),
            .I(n2325));
    LocalMux I__3969 (
            .O(N__28126),
            .I(n2325));
    LocalMux I__3968 (
            .O(N__28123),
            .I(n2325));
    InMux I__3967 (
            .O(N__28116),
            .I(n12645));
    InMux I__3966 (
            .O(N__28113),
            .I(n12646));
    InMux I__3965 (
            .O(N__28110),
            .I(n12647));
    InMux I__3964 (
            .O(N__28107),
            .I(n12648));
    InMux I__3963 (
            .O(N__28104),
            .I(n12649));
    InMux I__3962 (
            .O(N__28101),
            .I(bfn_5_18_0_));
    InMux I__3961 (
            .O(N__28098),
            .I(n12651));
    InMux I__3960 (
            .O(N__28095),
            .I(n12652));
    InMux I__3959 (
            .O(N__28092),
            .I(n12653));
    InMux I__3958 (
            .O(N__28089),
            .I(n12654));
    InMux I__3957 (
            .O(N__28086),
            .I(N__28082));
    InMux I__3956 (
            .O(N__28085),
            .I(N__28079));
    LocalMux I__3955 (
            .O(N__28082),
            .I(N__28076));
    LocalMux I__3954 (
            .O(N__28079),
            .I(N__28070));
    Span4Mux_s3_h I__3953 (
            .O(N__28076),
            .I(N__28070));
    InMux I__3952 (
            .O(N__28075),
            .I(N__28067));
    Span4Mux_v I__3951 (
            .O(N__28070),
            .I(N__28062));
    LocalMux I__3950 (
            .O(N__28067),
            .I(N__28062));
    Span4Mux_v I__3949 (
            .O(N__28062),
            .I(N__28059));
    Odrv4 I__3948 (
            .O(N__28059),
            .I(n2908));
    CascadeMux I__3947 (
            .O(N__28056),
            .I(N__28053));
    InMux I__3946 (
            .O(N__28053),
            .I(N__28050));
    LocalMux I__3945 (
            .O(N__28050),
            .I(N__28047));
    Odrv4 I__3944 (
            .O(N__28047),
            .I(n2975));
    InMux I__3943 (
            .O(N__28044),
            .I(N__28041));
    LocalMux I__3942 (
            .O(N__28041),
            .I(n3074));
    CascadeMux I__3941 (
            .O(N__28038),
            .I(n3007_cascade_));
    InMux I__3940 (
            .O(N__28035),
            .I(N__28032));
    LocalMux I__3939 (
            .O(N__28032),
            .I(N__28028));
    InMux I__3938 (
            .O(N__28031),
            .I(N__28025));
    Span12Mux_s4_v I__3937 (
            .O(N__28028),
            .I(N__28021));
    LocalMux I__3936 (
            .O(N__28025),
            .I(N__28018));
    InMux I__3935 (
            .O(N__28024),
            .I(N__28015));
    Odrv12 I__3934 (
            .O(N__28021),
            .I(n2910));
    Odrv12 I__3933 (
            .O(N__28018),
            .I(n2910));
    LocalMux I__3932 (
            .O(N__28015),
            .I(n2910));
    CascadeMux I__3931 (
            .O(N__28008),
            .I(N__28005));
    InMux I__3930 (
            .O(N__28005),
            .I(N__28002));
    LocalMux I__3929 (
            .O(N__28002),
            .I(N__27999));
    Odrv12 I__3928 (
            .O(N__27999),
            .I(n2977));
    InMux I__3927 (
            .O(N__27996),
            .I(N__27992));
    InMux I__3926 (
            .O(N__27995),
            .I(N__27989));
    LocalMux I__3925 (
            .O(N__27992),
            .I(N__27984));
    LocalMux I__3924 (
            .O(N__27989),
            .I(N__27984));
    Span4Mux_s2_v I__3923 (
            .O(N__27984),
            .I(N__27981));
    Odrv4 I__3922 (
            .O(N__27981),
            .I(\debounce.reg_A_2 ));
    SRMux I__3921 (
            .O(N__27978),
            .I(N__27975));
    LocalMux I__3920 (
            .O(N__27975),
            .I(N__27971));
    SRMux I__3919 (
            .O(N__27974),
            .I(N__27968));
    Span4Mux_v I__3918 (
            .O(N__27971),
            .I(N__27965));
    LocalMux I__3917 (
            .O(N__27968),
            .I(N__27962));
    Span4Mux_s1_h I__3916 (
            .O(N__27965),
            .I(N__27957));
    Span4Mux_s1_h I__3915 (
            .O(N__27962),
            .I(N__27957));
    Odrv4 I__3914 (
            .O(N__27957),
            .I(\debounce.cnt_next_9__N_424 ));
    InMux I__3913 (
            .O(N__27954),
            .I(bfn_5_17_0_));
    InMux I__3912 (
            .O(N__27951),
            .I(n12643));
    InMux I__3911 (
            .O(N__27948),
            .I(n12644));
    InMux I__3910 (
            .O(N__27945),
            .I(N__27942));
    LocalMux I__3909 (
            .O(N__27942),
            .I(N__27939));
    Span4Mux_v I__3908 (
            .O(N__27939),
            .I(N__27936));
    Odrv4 I__3907 (
            .O(N__27936),
            .I(n2985));
    InMux I__3906 (
            .O(N__27933),
            .I(N__27929));
    InMux I__3905 (
            .O(N__27932),
            .I(N__27926));
    LocalMux I__3904 (
            .O(N__27929),
            .I(N__27923));
    LocalMux I__3903 (
            .O(N__27926),
            .I(N__27920));
    Span4Mux_v I__3902 (
            .O(N__27923),
            .I(N__27917));
    Odrv12 I__3901 (
            .O(N__27920),
            .I(n2918));
    Odrv4 I__3900 (
            .O(N__27917),
            .I(n2918));
    InMux I__3899 (
            .O(N__27912),
            .I(N__27908));
    InMux I__3898 (
            .O(N__27911),
            .I(N__27905));
    LocalMux I__3897 (
            .O(N__27908),
            .I(N__27902));
    LocalMux I__3896 (
            .O(N__27905),
            .I(N__27899));
    Odrv4 I__3895 (
            .O(N__27902),
            .I(n2911));
    Odrv4 I__3894 (
            .O(N__27899),
            .I(n2911));
    InMux I__3893 (
            .O(N__27894),
            .I(N__27891));
    LocalMux I__3892 (
            .O(N__27891),
            .I(N__27888));
    Odrv4 I__3891 (
            .O(N__27888),
            .I(n2978));
    CascadeMux I__3890 (
            .O(N__27885),
            .I(N__27881));
    InMux I__3889 (
            .O(N__27884),
            .I(N__27878));
    InMux I__3888 (
            .O(N__27881),
            .I(N__27875));
    LocalMux I__3887 (
            .O(N__27878),
            .I(N__27872));
    LocalMux I__3886 (
            .O(N__27875),
            .I(N__27869));
    Span4Mux_s3_v I__3885 (
            .O(N__27872),
            .I(N__27865));
    Span4Mux_s2_h I__3884 (
            .O(N__27869),
            .I(N__27862));
    InMux I__3883 (
            .O(N__27868),
            .I(N__27859));
    Odrv4 I__3882 (
            .O(N__27865),
            .I(n2825));
    Odrv4 I__3881 (
            .O(N__27862),
            .I(n2825));
    LocalMux I__3880 (
            .O(N__27859),
            .I(n2825));
    CascadeMux I__3879 (
            .O(N__27852),
            .I(N__27849));
    InMux I__3878 (
            .O(N__27849),
            .I(N__27846));
    LocalMux I__3877 (
            .O(N__27846),
            .I(N__27843));
    Span4Mux_v I__3876 (
            .O(N__27843),
            .I(N__27840));
    Odrv4 I__3875 (
            .O(N__27840),
            .I(n2892));
    CascadeMux I__3874 (
            .O(N__27837),
            .I(N__27834));
    InMux I__3873 (
            .O(N__27834),
            .I(N__27830));
    InMux I__3872 (
            .O(N__27833),
            .I(N__27826));
    LocalMux I__3871 (
            .O(N__27830),
            .I(N__27823));
    InMux I__3870 (
            .O(N__27829),
            .I(N__27820));
    LocalMux I__3869 (
            .O(N__27826),
            .I(N__27817));
    Span4Mux_v I__3868 (
            .O(N__27823),
            .I(N__27814));
    LocalMux I__3867 (
            .O(N__27820),
            .I(N__27809));
    Span4Mux_h I__3866 (
            .O(N__27817),
            .I(N__27809));
    Odrv4 I__3865 (
            .O(N__27814),
            .I(n2924));
    Odrv4 I__3864 (
            .O(N__27809),
            .I(n2924));
    CascadeMux I__3863 (
            .O(N__27804),
            .I(N__27801));
    InMux I__3862 (
            .O(N__27801),
            .I(N__27797));
    InMux I__3861 (
            .O(N__27800),
            .I(N__27794));
    LocalMux I__3860 (
            .O(N__27797),
            .I(N__27791));
    LocalMux I__3859 (
            .O(N__27794),
            .I(N__27787));
    Span4Mux_v I__3858 (
            .O(N__27791),
            .I(N__27784));
    InMux I__3857 (
            .O(N__27790),
            .I(N__27781));
    Odrv12 I__3856 (
            .O(N__27787),
            .I(n2913));
    Odrv4 I__3855 (
            .O(N__27784),
            .I(n2913));
    LocalMux I__3854 (
            .O(N__27781),
            .I(n2913));
    CascadeMux I__3853 (
            .O(N__27774),
            .I(N__27771));
    InMux I__3852 (
            .O(N__27771),
            .I(N__27768));
    LocalMux I__3851 (
            .O(N__27768),
            .I(N__27765));
    Odrv12 I__3850 (
            .O(N__27765),
            .I(n2980));
    InMux I__3849 (
            .O(N__27762),
            .I(N__27758));
    InMux I__3848 (
            .O(N__27761),
            .I(N__27755));
    LocalMux I__3847 (
            .O(N__27758),
            .I(N__27752));
    LocalMux I__3846 (
            .O(N__27755),
            .I(N__27746));
    Span4Mux_s3_h I__3845 (
            .O(N__27752),
            .I(N__27746));
    InMux I__3844 (
            .O(N__27751),
            .I(N__27743));
    Span4Mux_v I__3843 (
            .O(N__27746),
            .I(N__27740));
    LocalMux I__3842 (
            .O(N__27743),
            .I(N__27737));
    Odrv4 I__3841 (
            .O(N__27740),
            .I(n2915));
    Odrv12 I__3840 (
            .O(N__27737),
            .I(n2915));
    CascadeMux I__3839 (
            .O(N__27732),
            .I(N__27729));
    InMux I__3838 (
            .O(N__27729),
            .I(N__27726));
    LocalMux I__3837 (
            .O(N__27726),
            .I(N__27723));
    Odrv4 I__3836 (
            .O(N__27723),
            .I(n2982));
    InMux I__3835 (
            .O(N__27720),
            .I(N__27717));
    LocalMux I__3834 (
            .O(N__27717),
            .I(N__27713));
    InMux I__3833 (
            .O(N__27716),
            .I(N__27710));
    Span4Mux_h I__3832 (
            .O(N__27713),
            .I(N__27704));
    LocalMux I__3831 (
            .O(N__27710),
            .I(N__27704));
    InMux I__3830 (
            .O(N__27709),
            .I(N__27701));
    Odrv4 I__3829 (
            .O(N__27704),
            .I(n2912));
    LocalMux I__3828 (
            .O(N__27701),
            .I(n2912));
    InMux I__3827 (
            .O(N__27696),
            .I(N__27693));
    LocalMux I__3826 (
            .O(N__27693),
            .I(N__27690));
    Odrv4 I__3825 (
            .O(N__27690),
            .I(n2979));
    InMux I__3824 (
            .O(N__27687),
            .I(N__27683));
    CascadeMux I__3823 (
            .O(N__27686),
            .I(N__27680));
    LocalMux I__3822 (
            .O(N__27683),
            .I(N__27677));
    InMux I__3821 (
            .O(N__27680),
            .I(N__27674));
    Span4Mux_v I__3820 (
            .O(N__27677),
            .I(N__27670));
    LocalMux I__3819 (
            .O(N__27674),
            .I(N__27667));
    InMux I__3818 (
            .O(N__27673),
            .I(N__27664));
    Odrv4 I__3817 (
            .O(N__27670),
            .I(n2919));
    Odrv4 I__3816 (
            .O(N__27667),
            .I(n2919));
    LocalMux I__3815 (
            .O(N__27664),
            .I(n2919));
    CascadeMux I__3814 (
            .O(N__27657),
            .I(N__27654));
    InMux I__3813 (
            .O(N__27654),
            .I(N__27651));
    LocalMux I__3812 (
            .O(N__27651),
            .I(N__27648));
    Span4Mux_s2_v I__3811 (
            .O(N__27648),
            .I(N__27645));
    Odrv4 I__3810 (
            .O(N__27645),
            .I(n2986));
    InMux I__3809 (
            .O(N__27642),
            .I(N__27637));
    InMux I__3808 (
            .O(N__27641),
            .I(N__27634));
    InMux I__3807 (
            .O(N__27640),
            .I(N__27631));
    LocalMux I__3806 (
            .O(N__27637),
            .I(n3016));
    LocalMux I__3805 (
            .O(N__27634),
            .I(n3016));
    LocalMux I__3804 (
            .O(N__27631),
            .I(n3016));
    CascadeMux I__3803 (
            .O(N__27624),
            .I(n3018_cascade_));
    InMux I__3802 (
            .O(N__27621),
            .I(N__27618));
    LocalMux I__3801 (
            .O(N__27618),
            .I(N__27614));
    InMux I__3800 (
            .O(N__27617),
            .I(N__27611));
    Span4Mux_s1_v I__3799 (
            .O(N__27614),
            .I(N__27607));
    LocalMux I__3798 (
            .O(N__27611),
            .I(N__27604));
    InMux I__3797 (
            .O(N__27610),
            .I(N__27601));
    Odrv4 I__3796 (
            .O(N__27607),
            .I(n2914));
    Odrv4 I__3795 (
            .O(N__27604),
            .I(n2914));
    LocalMux I__3794 (
            .O(N__27601),
            .I(n2914));
    CascadeMux I__3793 (
            .O(N__27594),
            .I(N__27591));
    InMux I__3792 (
            .O(N__27591),
            .I(N__27588));
    LocalMux I__3791 (
            .O(N__27588),
            .I(N__27585));
    Span4Mux_s1_v I__3790 (
            .O(N__27585),
            .I(N__27582));
    Odrv4 I__3789 (
            .O(N__27582),
            .I(n2981));
    CascadeMux I__3788 (
            .O(N__27579),
            .I(N__27576));
    InMux I__3787 (
            .O(N__27576),
            .I(N__27572));
    InMux I__3786 (
            .O(N__27575),
            .I(N__27568));
    LocalMux I__3785 (
            .O(N__27572),
            .I(N__27565));
    InMux I__3784 (
            .O(N__27571),
            .I(N__27562));
    LocalMux I__3783 (
            .O(N__27568),
            .I(n3019));
    Odrv4 I__3782 (
            .O(N__27565),
            .I(n3019));
    LocalMux I__3781 (
            .O(N__27562),
            .I(n3019));
    CascadeMux I__3780 (
            .O(N__27555),
            .I(n3023_cascade_));
    InMux I__3779 (
            .O(N__27552),
            .I(N__27548));
    InMux I__3778 (
            .O(N__27551),
            .I(N__27545));
    LocalMux I__3777 (
            .O(N__27548),
            .I(N__27541));
    LocalMux I__3776 (
            .O(N__27545),
            .I(N__27538));
    InMux I__3775 (
            .O(N__27544),
            .I(N__27535));
    Odrv4 I__3774 (
            .O(N__27541),
            .I(n2922));
    Odrv4 I__3773 (
            .O(N__27538),
            .I(n2922));
    LocalMux I__3772 (
            .O(N__27535),
            .I(n2922));
    CascadeMux I__3771 (
            .O(N__27528),
            .I(N__27525));
    InMux I__3770 (
            .O(N__27525),
            .I(N__27522));
    LocalMux I__3769 (
            .O(N__27522),
            .I(N__27519));
    Span4Mux_h I__3768 (
            .O(N__27519),
            .I(N__27516));
    Odrv4 I__3767 (
            .O(N__27516),
            .I(n2989));
    CascadeMux I__3766 (
            .O(N__27513),
            .I(N__27510));
    InMux I__3765 (
            .O(N__27510),
            .I(N__27507));
    LocalMux I__3764 (
            .O(N__27507),
            .I(n3078));
    InMux I__3763 (
            .O(N__27504),
            .I(N__27501));
    LocalMux I__3762 (
            .O(N__27501),
            .I(N__27498));
    Odrv4 I__3761 (
            .O(N__27498),
            .I(n3075));
    InMux I__3760 (
            .O(N__27495),
            .I(N__27492));
    LocalMux I__3759 (
            .O(N__27492),
            .I(N__27489));
    Span4Mux_v I__3758 (
            .O(N__27489),
            .I(N__27486));
    Odrv4 I__3757 (
            .O(N__27486),
            .I(n2984));
    CascadeMux I__3756 (
            .O(N__27483),
            .I(N__27479));
    InMux I__3755 (
            .O(N__27482),
            .I(N__27476));
    InMux I__3754 (
            .O(N__27479),
            .I(N__27473));
    LocalMux I__3753 (
            .O(N__27476),
            .I(N__27470));
    LocalMux I__3752 (
            .O(N__27473),
            .I(N__27466));
    Span4Mux_v I__3751 (
            .O(N__27470),
            .I(N__27463));
    InMux I__3750 (
            .O(N__27469),
            .I(N__27460));
    Odrv4 I__3749 (
            .O(N__27466),
            .I(n2917));
    Odrv4 I__3748 (
            .O(N__27463),
            .I(n2917));
    LocalMux I__3747 (
            .O(N__27460),
            .I(n2917));
    InMux I__3746 (
            .O(N__27453),
            .I(N__27449));
    CascadeMux I__3745 (
            .O(N__27452),
            .I(N__27446));
    LocalMux I__3744 (
            .O(N__27449),
            .I(N__27442));
    InMux I__3743 (
            .O(N__27446),
            .I(N__27439));
    InMux I__3742 (
            .O(N__27445),
            .I(N__27436));
    Odrv12 I__3741 (
            .O(N__27442),
            .I(n2931));
    LocalMux I__3740 (
            .O(N__27439),
            .I(n2931));
    LocalMux I__3739 (
            .O(N__27436),
            .I(n2931));
    CascadeMux I__3738 (
            .O(N__27429),
            .I(N__27426));
    InMux I__3737 (
            .O(N__27426),
            .I(N__27423));
    LocalMux I__3736 (
            .O(N__27423),
            .I(N__27420));
    Span4Mux_h I__3735 (
            .O(N__27420),
            .I(N__27417));
    Odrv4 I__3734 (
            .O(N__27417),
            .I(n2998));
    InMux I__3733 (
            .O(N__27414),
            .I(N__27411));
    LocalMux I__3732 (
            .O(N__27411),
            .I(n3097));
    CascadeMux I__3731 (
            .O(N__27408),
            .I(n3030_cascade_));
    CascadeMux I__3730 (
            .O(N__27405),
            .I(N__27401));
    InMux I__3729 (
            .O(N__27404),
            .I(N__27397));
    InMux I__3728 (
            .O(N__27401),
            .I(N__27394));
    InMux I__3727 (
            .O(N__27400),
            .I(N__27391));
    LocalMux I__3726 (
            .O(N__27397),
            .I(n3020));
    LocalMux I__3725 (
            .O(N__27394),
            .I(n3020));
    LocalMux I__3724 (
            .O(N__27391),
            .I(n3020));
    InMux I__3723 (
            .O(N__27384),
            .I(N__27381));
    LocalMux I__3722 (
            .O(N__27381),
            .I(n3087));
    CascadeMux I__3721 (
            .O(N__27378),
            .I(N__27375));
    InMux I__3720 (
            .O(N__27375),
            .I(N__27372));
    LocalMux I__3719 (
            .O(N__27372),
            .I(N__27368));
    InMux I__3718 (
            .O(N__27371),
            .I(N__27364));
    Span4Mux_s3_h I__3717 (
            .O(N__27368),
            .I(N__27361));
    InMux I__3716 (
            .O(N__27367),
            .I(N__27358));
    LocalMux I__3715 (
            .O(N__27364),
            .I(n2927));
    Odrv4 I__3714 (
            .O(N__27361),
            .I(n2927));
    LocalMux I__3713 (
            .O(N__27358),
            .I(n2927));
    CascadeMux I__3712 (
            .O(N__27351),
            .I(N__27348));
    InMux I__3711 (
            .O(N__27348),
            .I(N__27345));
    LocalMux I__3710 (
            .O(N__27345),
            .I(N__27342));
    Span4Mux_h I__3709 (
            .O(N__27342),
            .I(N__27339));
    Odrv4 I__3708 (
            .O(N__27339),
            .I(n2994));
    InMux I__3707 (
            .O(N__27336),
            .I(N__27329));
    InMux I__3706 (
            .O(N__27335),
            .I(N__27329));
    InMux I__3705 (
            .O(N__27334),
            .I(N__27326));
    LocalMux I__3704 (
            .O(N__27329),
            .I(N__27323));
    LocalMux I__3703 (
            .O(N__27326),
            .I(N__27320));
    Odrv12 I__3702 (
            .O(N__27323),
            .I(n2909));
    Odrv4 I__3701 (
            .O(N__27320),
            .I(n2909));
    CascadeMux I__3700 (
            .O(N__27315),
            .I(N__27312));
    InMux I__3699 (
            .O(N__27312),
            .I(N__27308));
    InMux I__3698 (
            .O(N__27311),
            .I(N__27305));
    LocalMux I__3697 (
            .O(N__27308),
            .I(N__27302));
    LocalMux I__3696 (
            .O(N__27305),
            .I(N__27299));
    Span4Mux_h I__3695 (
            .O(N__27302),
            .I(N__27296));
    Odrv4 I__3694 (
            .O(N__27299),
            .I(n2907));
    Odrv4 I__3693 (
            .O(N__27296),
            .I(n2907));
    InMux I__3692 (
            .O(N__27291),
            .I(N__27288));
    LocalMux I__3691 (
            .O(N__27288),
            .I(n14372));
    CascadeMux I__3690 (
            .O(N__27285),
            .I(N__27280));
    InMux I__3689 (
            .O(N__27284),
            .I(N__27275));
    InMux I__3688 (
            .O(N__27283),
            .I(N__27275));
    InMux I__3687 (
            .O(N__27280),
            .I(N__27272));
    LocalMux I__3686 (
            .O(N__27275),
            .I(N__27269));
    LocalMux I__3685 (
            .O(N__27272),
            .I(n2929));
    Odrv4 I__3684 (
            .O(N__27269),
            .I(n2929));
    CascadeMux I__3683 (
            .O(N__27264),
            .I(n2940_cascade_));
    InMux I__3682 (
            .O(N__27261),
            .I(N__27258));
    LocalMux I__3681 (
            .O(N__27258),
            .I(N__27255));
    Span4Mux_h I__3680 (
            .O(N__27255),
            .I(N__27252));
    Odrv4 I__3679 (
            .O(N__27252),
            .I(n2996));
    InMux I__3678 (
            .O(N__27249),
            .I(N__27245));
    InMux I__3677 (
            .O(N__27248),
            .I(N__27242));
    LocalMux I__3676 (
            .O(N__27245),
            .I(N__27239));
    LocalMux I__3675 (
            .O(N__27242),
            .I(N__27236));
    Span4Mux_v I__3674 (
            .O(N__27239),
            .I(N__27233));
    Odrv4 I__3673 (
            .O(N__27236),
            .I(n2921));
    Odrv4 I__3672 (
            .O(N__27233),
            .I(n2921));
    InMux I__3671 (
            .O(N__27228),
            .I(N__27225));
    LocalMux I__3670 (
            .O(N__27225),
            .I(N__27222));
    Span4Mux_h I__3669 (
            .O(N__27222),
            .I(N__27219));
    Odrv4 I__3668 (
            .O(N__27219),
            .I(n2988));
    InMux I__3667 (
            .O(N__27216),
            .I(N__27213));
    LocalMux I__3666 (
            .O(N__27213),
            .I(N__27210));
    Odrv4 I__3665 (
            .O(N__27210),
            .I(n3083));
    InMux I__3664 (
            .O(N__27207),
            .I(N__27204));
    LocalMux I__3663 (
            .O(N__27204),
            .I(N__27201));
    Odrv4 I__3662 (
            .O(N__27201),
            .I(n2995));
    CascadeMux I__3661 (
            .O(N__27198),
            .I(N__27194));
    InMux I__3660 (
            .O(N__27197),
            .I(N__27190));
    InMux I__3659 (
            .O(N__27194),
            .I(N__27187));
    InMux I__3658 (
            .O(N__27193),
            .I(N__27184));
    LocalMux I__3657 (
            .O(N__27190),
            .I(n2928));
    LocalMux I__3656 (
            .O(N__27187),
            .I(n2928));
    LocalMux I__3655 (
            .O(N__27184),
            .I(n2928));
    InMux I__3654 (
            .O(N__27177),
            .I(N__27174));
    LocalMux I__3653 (
            .O(N__27174),
            .I(N__27171));
    Odrv4 I__3652 (
            .O(N__27171),
            .I(n2997));
    CascadeMux I__3651 (
            .O(N__27168),
            .I(N__27164));
    CascadeMux I__3650 (
            .O(N__27167),
            .I(N__27161));
    InMux I__3649 (
            .O(N__27164),
            .I(N__27157));
    InMux I__3648 (
            .O(N__27161),
            .I(N__27154));
    InMux I__3647 (
            .O(N__27160),
            .I(N__27151));
    LocalMux I__3646 (
            .O(N__27157),
            .I(n2930));
    LocalMux I__3645 (
            .O(N__27154),
            .I(n2930));
    LocalMux I__3644 (
            .O(N__27151),
            .I(n2930));
    InMux I__3643 (
            .O(N__27144),
            .I(N__27141));
    LocalMux I__3642 (
            .O(N__27141),
            .I(n3096));
    CascadeMux I__3641 (
            .O(N__27138),
            .I(n3029_cascade_));
    CascadeMux I__3640 (
            .O(N__27135),
            .I(N__27132));
    InMux I__3639 (
            .O(N__27132),
            .I(N__27129));
    LocalMux I__3638 (
            .O(N__27129),
            .I(N__27126));
    Span4Mux_h I__3637 (
            .O(N__27126),
            .I(N__27123));
    Odrv4 I__3636 (
            .O(N__27123),
            .I(n2991));
    CascadeMux I__3635 (
            .O(N__27120),
            .I(n2926_cascade_));
    InMux I__3634 (
            .O(N__27117),
            .I(N__27114));
    LocalMux I__3633 (
            .O(N__27114),
            .I(n14346));
    CascadeMux I__3632 (
            .O(N__27111),
            .I(n14336_cascade_));
    CascadeMux I__3631 (
            .O(N__27108),
            .I(n14352_cascade_));
    InMux I__3630 (
            .O(N__27105),
            .I(N__27102));
    LocalMux I__3629 (
            .O(N__27102),
            .I(n14350));
    CascadeMux I__3628 (
            .O(N__27099),
            .I(N__27096));
    InMux I__3627 (
            .O(N__27096),
            .I(N__27092));
    InMux I__3626 (
            .O(N__27095),
            .I(N__27088));
    LocalMux I__3625 (
            .O(N__27092),
            .I(N__27085));
    InMux I__3624 (
            .O(N__27091),
            .I(N__27082));
    LocalMux I__3623 (
            .O(N__27088),
            .I(n2828));
    Odrv4 I__3622 (
            .O(N__27085),
            .I(n2828));
    LocalMux I__3621 (
            .O(N__27082),
            .I(n2828));
    CascadeMux I__3620 (
            .O(N__27075),
            .I(N__27072));
    InMux I__3619 (
            .O(N__27072),
            .I(N__27069));
    LocalMux I__3618 (
            .O(N__27069),
            .I(N__27066));
    Span4Mux_h I__3617 (
            .O(N__27066),
            .I(N__27063));
    Odrv4 I__3616 (
            .O(N__27063),
            .I(n2895));
    InMux I__3615 (
            .O(N__27060),
            .I(N__27057));
    LocalMux I__3614 (
            .O(N__27057),
            .I(N__27054));
    Span4Mux_v I__3613 (
            .O(N__27054),
            .I(N__27051));
    Odrv4 I__3612 (
            .O(N__27051),
            .I(n2885));
    InMux I__3611 (
            .O(N__27048),
            .I(N__27045));
    LocalMux I__3610 (
            .O(N__27045),
            .I(N__27041));
    InMux I__3609 (
            .O(N__27044),
            .I(N__27038));
    Span4Mux_h I__3608 (
            .O(N__27041),
            .I(N__27034));
    LocalMux I__3607 (
            .O(N__27038),
            .I(N__27031));
    InMux I__3606 (
            .O(N__27037),
            .I(N__27028));
    Odrv4 I__3605 (
            .O(N__27034),
            .I(n2818));
    Odrv12 I__3604 (
            .O(N__27031),
            .I(n2818));
    LocalMux I__3603 (
            .O(N__27028),
            .I(n2818));
    InMux I__3602 (
            .O(N__27021),
            .I(N__27018));
    LocalMux I__3601 (
            .O(N__27018),
            .I(N__27015));
    Odrv4 I__3600 (
            .O(N__27015),
            .I(n2881));
    CascadeMux I__3599 (
            .O(N__27012),
            .I(N__27009));
    InMux I__3598 (
            .O(N__27009),
            .I(N__27006));
    LocalMux I__3597 (
            .O(N__27006),
            .I(N__27002));
    InMux I__3596 (
            .O(N__27005),
            .I(N__26999));
    Span4Mux_h I__3595 (
            .O(N__27002),
            .I(N__26993));
    LocalMux I__3594 (
            .O(N__26999),
            .I(N__26993));
    InMux I__3593 (
            .O(N__26998),
            .I(N__26990));
    Odrv4 I__3592 (
            .O(N__26993),
            .I(n2814));
    LocalMux I__3591 (
            .O(N__26990),
            .I(n2814));
    CascadeMux I__3590 (
            .O(N__26985),
            .I(N__26982));
    InMux I__3589 (
            .O(N__26982),
            .I(N__26979));
    LocalMux I__3588 (
            .O(N__26979),
            .I(N__26976));
    Span4Mux_v I__3587 (
            .O(N__26976),
            .I(N__26973));
    Odrv4 I__3586 (
            .O(N__26973),
            .I(n12038));
    InMux I__3585 (
            .O(N__26970),
            .I(N__26967));
    LocalMux I__3584 (
            .O(N__26967),
            .I(n14358));
    CascadeMux I__3583 (
            .O(N__26964),
            .I(n14360_cascade_));
    InMux I__3582 (
            .O(N__26961),
            .I(N__26958));
    LocalMux I__3581 (
            .O(N__26958),
            .I(n14366));
    CascadeMux I__3580 (
            .O(N__26955),
            .I(N__26952));
    InMux I__3579 (
            .O(N__26952),
            .I(N__26949));
    LocalMux I__3578 (
            .O(N__26949),
            .I(N__26946));
    Span4Mux_h I__3577 (
            .O(N__26946),
            .I(N__26943));
    Odrv4 I__3576 (
            .O(N__26943),
            .I(n3094));
    InMux I__3575 (
            .O(N__26940),
            .I(N__26937));
    LocalMux I__3574 (
            .O(N__26937),
            .I(N__26934));
    Span4Mux_v I__3573 (
            .O(N__26934),
            .I(N__26931));
    Odrv4 I__3572 (
            .O(N__26931),
            .I(n2701));
    CascadeMux I__3571 (
            .O(N__26928),
            .I(N__26924));
    InMux I__3570 (
            .O(N__26927),
            .I(N__26921));
    InMux I__3569 (
            .O(N__26924),
            .I(N__26918));
    LocalMux I__3568 (
            .O(N__26921),
            .I(N__26915));
    LocalMux I__3567 (
            .O(N__26918),
            .I(N__26912));
    Span4Mux_s3_h I__3566 (
            .O(N__26915),
            .I(N__26907));
    Span4Mux_s3_h I__3565 (
            .O(N__26912),
            .I(N__26907));
    Odrv4 I__3564 (
            .O(N__26907),
            .I(n2733));
    CascadeMux I__3563 (
            .O(N__26904),
            .I(n2733_cascade_));
    CascadeMux I__3562 (
            .O(N__26901),
            .I(N__26898));
    InMux I__3561 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__3560 (
            .O(N__26895),
            .I(N__26890));
    InMux I__3559 (
            .O(N__26894),
            .I(N__26887));
    CascadeMux I__3558 (
            .O(N__26893),
            .I(N__26884));
    Span4Mux_s3_h I__3557 (
            .O(N__26890),
            .I(N__26879));
    LocalMux I__3556 (
            .O(N__26887),
            .I(N__26879));
    InMux I__3555 (
            .O(N__26884),
            .I(N__26876));
    Span4Mux_v I__3554 (
            .O(N__26879),
            .I(N__26873));
    LocalMux I__3553 (
            .O(N__26876),
            .I(n2732));
    Odrv4 I__3552 (
            .O(N__26873),
            .I(n2732));
    InMux I__3551 (
            .O(N__26868),
            .I(N__26865));
    LocalMux I__3550 (
            .O(N__26865),
            .I(n11936));
    CascadeMux I__3549 (
            .O(N__26862),
            .I(N__26859));
    InMux I__3548 (
            .O(N__26859),
            .I(N__26856));
    LocalMux I__3547 (
            .O(N__26856),
            .I(N__26852));
    InMux I__3546 (
            .O(N__26855),
            .I(N__26849));
    Span4Mux_h I__3545 (
            .O(N__26852),
            .I(N__26846));
    LocalMux I__3544 (
            .O(N__26849),
            .I(n2729));
    Odrv4 I__3543 (
            .O(N__26846),
            .I(n2729));
    CascadeMux I__3542 (
            .O(N__26841),
            .I(N__26838));
    InMux I__3541 (
            .O(N__26838),
            .I(N__26835));
    LocalMux I__3540 (
            .O(N__26835),
            .I(N__26832));
    Span4Mux_h I__3539 (
            .O(N__26832),
            .I(N__26829));
    Odrv4 I__3538 (
            .O(N__26829),
            .I(n2796));
    InMux I__3537 (
            .O(N__26826),
            .I(N__26823));
    LocalMux I__3536 (
            .O(N__26823),
            .I(N__26819));
    InMux I__3535 (
            .O(N__26822),
            .I(N__26815));
    Span4Mux_s2_h I__3534 (
            .O(N__26819),
            .I(N__26812));
    InMux I__3533 (
            .O(N__26818),
            .I(N__26809));
    LocalMux I__3532 (
            .O(N__26815),
            .I(n2819));
    Odrv4 I__3531 (
            .O(N__26812),
            .I(n2819));
    LocalMux I__3530 (
            .O(N__26809),
            .I(n2819));
    CascadeMux I__3529 (
            .O(N__26802),
            .I(N__26799));
    InMux I__3528 (
            .O(N__26799),
            .I(N__26796));
    LocalMux I__3527 (
            .O(N__26796),
            .I(N__26793));
    Odrv12 I__3526 (
            .O(N__26793),
            .I(n2886));
    CascadeMux I__3525 (
            .O(N__26790),
            .I(n2918_cascade_));
    CascadeMux I__3524 (
            .O(N__26787),
            .I(N__26784));
    InMux I__3523 (
            .O(N__26784),
            .I(N__26780));
    InMux I__3522 (
            .O(N__26783),
            .I(N__26776));
    LocalMux I__3521 (
            .O(N__26780),
            .I(N__26773));
    InMux I__3520 (
            .O(N__26779),
            .I(N__26770));
    LocalMux I__3519 (
            .O(N__26776),
            .I(n2827));
    Odrv4 I__3518 (
            .O(N__26773),
            .I(n2827));
    LocalMux I__3517 (
            .O(N__26770),
            .I(n2827));
    CascadeMux I__3516 (
            .O(N__26763),
            .I(N__26760));
    InMux I__3515 (
            .O(N__26760),
            .I(N__26757));
    LocalMux I__3514 (
            .O(N__26757),
            .I(N__26754));
    Span4Mux_h I__3513 (
            .O(N__26754),
            .I(N__26751));
    Odrv4 I__3512 (
            .O(N__26751),
            .I(n2894));
    CascadeMux I__3511 (
            .O(N__26748),
            .I(N__26745));
    InMux I__3510 (
            .O(N__26745),
            .I(N__26742));
    LocalMux I__3509 (
            .O(N__26742),
            .I(N__26739));
    Odrv4 I__3508 (
            .O(N__26739),
            .I(n2688));
    InMux I__3507 (
            .O(N__26736),
            .I(N__26732));
    InMux I__3506 (
            .O(N__26735),
            .I(N__26729));
    LocalMux I__3505 (
            .O(N__26732),
            .I(N__26726));
    LocalMux I__3504 (
            .O(N__26729),
            .I(N__26723));
    Odrv4 I__3503 (
            .O(N__26726),
            .I(n2720));
    Odrv4 I__3502 (
            .O(N__26723),
            .I(n2720));
    CascadeMux I__3501 (
            .O(N__26718),
            .I(N__26714));
    InMux I__3500 (
            .O(N__26717),
            .I(N__26710));
    InMux I__3499 (
            .O(N__26714),
            .I(N__26707));
    InMux I__3498 (
            .O(N__26713),
            .I(N__26704));
    LocalMux I__3497 (
            .O(N__26710),
            .I(n2726));
    LocalMux I__3496 (
            .O(N__26707),
            .I(n2726));
    LocalMux I__3495 (
            .O(N__26704),
            .I(n2726));
    InMux I__3494 (
            .O(N__26697),
            .I(N__26693));
    CascadeMux I__3493 (
            .O(N__26696),
            .I(N__26690));
    LocalMux I__3492 (
            .O(N__26693),
            .I(N__26686));
    InMux I__3491 (
            .O(N__26690),
            .I(N__26683));
    InMux I__3490 (
            .O(N__26689),
            .I(N__26680));
    Odrv12 I__3489 (
            .O(N__26686),
            .I(n2724));
    LocalMux I__3488 (
            .O(N__26683),
            .I(n2724));
    LocalMux I__3487 (
            .O(N__26680),
            .I(n2724));
    CascadeMux I__3486 (
            .O(N__26673),
            .I(n2720_cascade_));
    InMux I__3485 (
            .O(N__26670),
            .I(N__26666));
    CascadeMux I__3484 (
            .O(N__26669),
            .I(N__26663));
    LocalMux I__3483 (
            .O(N__26666),
            .I(N__26659));
    InMux I__3482 (
            .O(N__26663),
            .I(N__26656));
    InMux I__3481 (
            .O(N__26662),
            .I(N__26653));
    Odrv4 I__3480 (
            .O(N__26659),
            .I(n2723));
    LocalMux I__3479 (
            .O(N__26656),
            .I(n2723));
    LocalMux I__3478 (
            .O(N__26653),
            .I(n2723));
    InMux I__3477 (
            .O(N__26646),
            .I(N__26643));
    LocalMux I__3476 (
            .O(N__26643),
            .I(n14136));
    CascadeMux I__3475 (
            .O(N__26640),
            .I(N__26637));
    InMux I__3474 (
            .O(N__26637),
            .I(N__26634));
    LocalMux I__3473 (
            .O(N__26634),
            .I(N__26631));
    Span4Mux_v I__3472 (
            .O(N__26631),
            .I(N__26628));
    Odrv4 I__3471 (
            .O(N__26628),
            .I(n2699));
    InMux I__3470 (
            .O(N__26625),
            .I(N__26622));
    LocalMux I__3469 (
            .O(N__26622),
            .I(N__26619));
    Odrv12 I__3468 (
            .O(N__26619),
            .I(n2698));
    CascadeMux I__3467 (
            .O(N__26616),
            .I(N__26613));
    InMux I__3466 (
            .O(N__26613),
            .I(N__26610));
    LocalMux I__3465 (
            .O(N__26610),
            .I(N__26606));
    InMux I__3464 (
            .O(N__26609),
            .I(N__26602));
    Span4Mux_s2_h I__3463 (
            .O(N__26606),
            .I(N__26599));
    InMux I__3462 (
            .O(N__26605),
            .I(N__26596));
    LocalMux I__3461 (
            .O(N__26602),
            .I(n2820));
    Odrv4 I__3460 (
            .O(N__26599),
            .I(n2820));
    LocalMux I__3459 (
            .O(N__26596),
            .I(n2820));
    CascadeMux I__3458 (
            .O(N__26589),
            .I(n14688_cascade_));
    InMux I__3457 (
            .O(N__26586),
            .I(N__26583));
    LocalMux I__3456 (
            .O(N__26583),
            .I(N__26580));
    Odrv4 I__3455 (
            .O(N__26580),
            .I(n14690));
    InMux I__3454 (
            .O(N__26577),
            .I(N__26574));
    LocalMux I__3453 (
            .O(N__26574),
            .I(N__26571));
    Odrv4 I__3452 (
            .O(N__26571),
            .I(n14696));
    InMux I__3451 (
            .O(N__26568),
            .I(N__26565));
    LocalMux I__3450 (
            .O(N__26565),
            .I(N__26562));
    Span4Mux_v I__3449 (
            .O(N__26562),
            .I(N__26559));
    Span4Mux_h I__3448 (
            .O(N__26559),
            .I(N__26556));
    Span4Mux_v I__3447 (
            .O(N__26556),
            .I(N__26553));
    Odrv4 I__3446 (
            .O(N__26553),
            .I(ENCODER0_B_N));
    InMux I__3445 (
            .O(N__26550),
            .I(N__26547));
    LocalMux I__3444 (
            .O(N__26547),
            .I(N__26544));
    Odrv12 I__3443 (
            .O(N__26544),
            .I(n2697));
    CascadeMux I__3442 (
            .O(N__26541),
            .I(N__26538));
    InMux I__3441 (
            .O(N__26538),
            .I(N__26534));
    CascadeMux I__3440 (
            .O(N__26537),
            .I(N__26531));
    LocalMux I__3439 (
            .O(N__26534),
            .I(N__26527));
    InMux I__3438 (
            .O(N__26531),
            .I(N__26524));
    InMux I__3437 (
            .O(N__26530),
            .I(N__26521));
    Odrv4 I__3436 (
            .O(N__26527),
            .I(n2630));
    LocalMux I__3435 (
            .O(N__26524),
            .I(n2630));
    LocalMux I__3434 (
            .O(N__26521),
            .I(n2630));
    CascadeMux I__3433 (
            .O(N__26514),
            .I(N__26510));
    CascadeMux I__3432 (
            .O(N__26513),
            .I(N__26507));
    InMux I__3431 (
            .O(N__26510),
            .I(N__26504));
    InMux I__3430 (
            .O(N__26507),
            .I(N__26501));
    LocalMux I__3429 (
            .O(N__26504),
            .I(N__26498));
    LocalMux I__3428 (
            .O(N__26501),
            .I(N__26494));
    Span4Mux_s1_h I__3427 (
            .O(N__26498),
            .I(N__26491));
    InMux I__3426 (
            .O(N__26497),
            .I(N__26488));
    Span4Mux_s3_h I__3425 (
            .O(N__26494),
            .I(N__26485));
    Odrv4 I__3424 (
            .O(N__26491),
            .I(n2731));
    LocalMux I__3423 (
            .O(N__26488),
            .I(n2731));
    Odrv4 I__3422 (
            .O(N__26485),
            .I(n2731));
    CascadeMux I__3421 (
            .O(N__26478),
            .I(N__26475));
    InMux I__3420 (
            .O(N__26475),
            .I(N__26471));
    InMux I__3419 (
            .O(N__26474),
            .I(N__26468));
    LocalMux I__3418 (
            .O(N__26471),
            .I(N__26464));
    LocalMux I__3417 (
            .O(N__26468),
            .I(N__26461));
    InMux I__3416 (
            .O(N__26467),
            .I(N__26458));
    Span4Mux_s3_h I__3415 (
            .O(N__26464),
            .I(N__26455));
    Odrv12 I__3414 (
            .O(N__26461),
            .I(n2730));
    LocalMux I__3413 (
            .O(N__26458),
            .I(n2730));
    Odrv4 I__3412 (
            .O(N__26455),
            .I(n2730));
    CascadeMux I__3411 (
            .O(N__26448),
            .I(n2729_cascade_));
    InMux I__3410 (
            .O(N__26445),
            .I(N__26442));
    LocalMux I__3409 (
            .O(N__26442),
            .I(n13796));
    InMux I__3408 (
            .O(N__26439),
            .I(N__26436));
    LocalMux I__3407 (
            .O(N__26436),
            .I(N__26432));
    InMux I__3406 (
            .O(N__26435),
            .I(N__26429));
    Odrv12 I__3405 (
            .O(N__26432),
            .I(n2613));
    LocalMux I__3404 (
            .O(N__26429),
            .I(n2613));
    InMux I__3403 (
            .O(N__26424),
            .I(N__26421));
    LocalMux I__3402 (
            .O(N__26421),
            .I(N__26418));
    Odrv4 I__3401 (
            .O(N__26418),
            .I(n2680));
    InMux I__3400 (
            .O(N__26415),
            .I(n12768));
    InMux I__3399 (
            .O(N__26412),
            .I(N__26409));
    LocalMux I__3398 (
            .O(N__26409),
            .I(N__26405));
    InMux I__3397 (
            .O(N__26408),
            .I(N__26402));
    Span4Mux_h I__3396 (
            .O(N__26405),
            .I(N__26399));
    LocalMux I__3395 (
            .O(N__26402),
            .I(N__26396));
    Odrv4 I__3394 (
            .O(N__26399),
            .I(n2612));
    Odrv4 I__3393 (
            .O(N__26396),
            .I(n2612));
    InMux I__3392 (
            .O(N__26391),
            .I(N__26388));
    LocalMux I__3391 (
            .O(N__26388),
            .I(N__26385));
    Span4Mux_s3_h I__3390 (
            .O(N__26385),
            .I(N__26382));
    Odrv4 I__3389 (
            .O(N__26382),
            .I(n2679));
    InMux I__3388 (
            .O(N__26379),
            .I(n12769));
    InMux I__3387 (
            .O(N__26376),
            .I(N__26372));
    InMux I__3386 (
            .O(N__26375),
            .I(N__26369));
    LocalMux I__3385 (
            .O(N__26372),
            .I(N__26365));
    LocalMux I__3384 (
            .O(N__26369),
            .I(N__26362));
    InMux I__3383 (
            .O(N__26368),
            .I(N__26359));
    Span4Mux_h I__3382 (
            .O(N__26365),
            .I(N__26356));
    Span4Mux_v I__3381 (
            .O(N__26362),
            .I(N__26351));
    LocalMux I__3380 (
            .O(N__26359),
            .I(N__26351));
    Odrv4 I__3379 (
            .O(N__26356),
            .I(n2611));
    Odrv4 I__3378 (
            .O(N__26351),
            .I(n2611));
    CascadeMux I__3377 (
            .O(N__26346),
            .I(N__26343));
    InMux I__3376 (
            .O(N__26343),
            .I(N__26340));
    LocalMux I__3375 (
            .O(N__26340),
            .I(N__26337));
    Span4Mux_h I__3374 (
            .O(N__26337),
            .I(N__26334));
    Odrv4 I__3373 (
            .O(N__26334),
            .I(n2678));
    InMux I__3372 (
            .O(N__26331),
            .I(n12770));
    CascadeMux I__3371 (
            .O(N__26328),
            .I(N__26325));
    InMux I__3370 (
            .O(N__26325),
            .I(N__26322));
    LocalMux I__3369 (
            .O(N__26322),
            .I(N__26318));
    InMux I__3368 (
            .O(N__26321),
            .I(N__26315));
    Span4Mux_h I__3367 (
            .O(N__26318),
            .I(N__26312));
    LocalMux I__3366 (
            .O(N__26315),
            .I(N__26309));
    Span4Mux_s0_h I__3365 (
            .O(N__26312),
            .I(N__26304));
    Span4Mux_h I__3364 (
            .O(N__26309),
            .I(N__26304));
    Odrv4 I__3363 (
            .O(N__26304),
            .I(n2610));
    InMux I__3362 (
            .O(N__26301),
            .I(bfn_4_24_0_));
    InMux I__3361 (
            .O(N__26298),
            .I(N__26292));
    InMux I__3360 (
            .O(N__26297),
            .I(N__26292));
    LocalMux I__3359 (
            .O(N__26292),
            .I(N__26289));
    Span4Mux_s3_h I__3358 (
            .O(N__26289),
            .I(N__26286));
    Odrv4 I__3357 (
            .O(N__26286),
            .I(n2709));
    InMux I__3356 (
            .O(N__26283),
            .I(N__26279));
    InMux I__3355 (
            .O(N__26282),
            .I(N__26276));
    LocalMux I__3354 (
            .O(N__26279),
            .I(N__26273));
    LocalMux I__3353 (
            .O(N__26276),
            .I(N__26270));
    Odrv4 I__3352 (
            .O(N__26273),
            .I(n2816));
    Odrv12 I__3351 (
            .O(N__26270),
            .I(n2816));
    CascadeMux I__3350 (
            .O(N__26265),
            .I(N__26262));
    InMux I__3349 (
            .O(N__26262),
            .I(N__26259));
    LocalMux I__3348 (
            .O(N__26259),
            .I(N__26256));
    Span4Mux_h I__3347 (
            .O(N__26256),
            .I(N__26253));
    Odrv4 I__3346 (
            .O(N__26253),
            .I(n2883));
    InMux I__3345 (
            .O(N__26250),
            .I(N__26246));
    InMux I__3344 (
            .O(N__26249),
            .I(N__26243));
    LocalMux I__3343 (
            .O(N__26246),
            .I(N__26237));
    LocalMux I__3342 (
            .O(N__26243),
            .I(N__26237));
    CascadeMux I__3341 (
            .O(N__26242),
            .I(N__26234));
    Span4Mux_v I__3340 (
            .O(N__26237),
            .I(N__26231));
    InMux I__3339 (
            .O(N__26234),
            .I(N__26228));
    Odrv4 I__3338 (
            .O(N__26231),
            .I(n2621));
    LocalMux I__3337 (
            .O(N__26228),
            .I(n2621));
    InMux I__3336 (
            .O(N__26223),
            .I(n12760));
    InMux I__3335 (
            .O(N__26220),
            .I(N__26216));
    InMux I__3334 (
            .O(N__26219),
            .I(N__26212));
    LocalMux I__3333 (
            .O(N__26216),
            .I(N__26209));
    InMux I__3332 (
            .O(N__26215),
            .I(N__26206));
    LocalMux I__3331 (
            .O(N__26212),
            .I(n2620));
    Odrv4 I__3330 (
            .O(N__26209),
            .I(n2620));
    LocalMux I__3329 (
            .O(N__26206),
            .I(n2620));
    CascadeMux I__3328 (
            .O(N__26199),
            .I(N__26196));
    InMux I__3327 (
            .O(N__26196),
            .I(N__26193));
    LocalMux I__3326 (
            .O(N__26193),
            .I(N__26190));
    Span4Mux_s3_h I__3325 (
            .O(N__26190),
            .I(N__26187));
    Odrv4 I__3324 (
            .O(N__26187),
            .I(n2687));
    InMux I__3323 (
            .O(N__26184),
            .I(n12761));
    InMux I__3322 (
            .O(N__26181),
            .I(N__26178));
    LocalMux I__3321 (
            .O(N__26178),
            .I(N__26174));
    InMux I__3320 (
            .O(N__26177),
            .I(N__26170));
    Span4Mux_v I__3319 (
            .O(N__26174),
            .I(N__26167));
    InMux I__3318 (
            .O(N__26173),
            .I(N__26164));
    LocalMux I__3317 (
            .O(N__26170),
            .I(n2619));
    Odrv4 I__3316 (
            .O(N__26167),
            .I(n2619));
    LocalMux I__3315 (
            .O(N__26164),
            .I(n2619));
    CascadeMux I__3314 (
            .O(N__26157),
            .I(N__26154));
    InMux I__3313 (
            .O(N__26154),
            .I(N__26151));
    LocalMux I__3312 (
            .O(N__26151),
            .I(n2686));
    InMux I__3311 (
            .O(N__26148),
            .I(n12762));
    CascadeMux I__3310 (
            .O(N__26145),
            .I(N__26142));
    InMux I__3309 (
            .O(N__26142),
            .I(N__26139));
    LocalMux I__3308 (
            .O(N__26139),
            .I(N__26135));
    InMux I__3307 (
            .O(N__26138),
            .I(N__26132));
    Span4Mux_v I__3306 (
            .O(N__26135),
            .I(N__26129));
    LocalMux I__3305 (
            .O(N__26132),
            .I(N__26126));
    Span4Mux_s2_h I__3304 (
            .O(N__26129),
            .I(N__26122));
    Span4Mux_v I__3303 (
            .O(N__26126),
            .I(N__26119));
    InMux I__3302 (
            .O(N__26125),
            .I(N__26116));
    Odrv4 I__3301 (
            .O(N__26122),
            .I(n2618));
    Odrv4 I__3300 (
            .O(N__26119),
            .I(n2618));
    LocalMux I__3299 (
            .O(N__26116),
            .I(n2618));
    InMux I__3298 (
            .O(N__26109),
            .I(N__26106));
    LocalMux I__3297 (
            .O(N__26106),
            .I(n2685));
    InMux I__3296 (
            .O(N__26103),
            .I(bfn_4_23_0_));
    CascadeMux I__3295 (
            .O(N__26100),
            .I(N__26096));
    InMux I__3294 (
            .O(N__26099),
            .I(N__26093));
    InMux I__3293 (
            .O(N__26096),
            .I(N__26090));
    LocalMux I__3292 (
            .O(N__26093),
            .I(n2617));
    LocalMux I__3291 (
            .O(N__26090),
            .I(n2617));
    InMux I__3290 (
            .O(N__26085),
            .I(N__26082));
    LocalMux I__3289 (
            .O(N__26082),
            .I(n2684));
    InMux I__3288 (
            .O(N__26079),
            .I(n12764));
    InMux I__3287 (
            .O(N__26076),
            .I(N__26071));
    InMux I__3286 (
            .O(N__26075),
            .I(N__26068));
    InMux I__3285 (
            .O(N__26074),
            .I(N__26065));
    LocalMux I__3284 (
            .O(N__26071),
            .I(N__26060));
    LocalMux I__3283 (
            .O(N__26068),
            .I(N__26060));
    LocalMux I__3282 (
            .O(N__26065),
            .I(n2616));
    Odrv4 I__3281 (
            .O(N__26060),
            .I(n2616));
    InMux I__3280 (
            .O(N__26055),
            .I(N__26052));
    LocalMux I__3279 (
            .O(N__26052),
            .I(N__26049));
    Odrv4 I__3278 (
            .O(N__26049),
            .I(n2683));
    InMux I__3277 (
            .O(N__26046),
            .I(n12765));
    InMux I__3276 (
            .O(N__26043),
            .I(N__26040));
    LocalMux I__3275 (
            .O(N__26040),
            .I(N__26036));
    InMux I__3274 (
            .O(N__26039),
            .I(N__26033));
    Span4Mux_s3_h I__3273 (
            .O(N__26036),
            .I(N__26027));
    LocalMux I__3272 (
            .O(N__26033),
            .I(N__26027));
    InMux I__3271 (
            .O(N__26032),
            .I(N__26024));
    Span4Mux_v I__3270 (
            .O(N__26027),
            .I(N__26021));
    LocalMux I__3269 (
            .O(N__26024),
            .I(N__26018));
    Odrv4 I__3268 (
            .O(N__26021),
            .I(n2615));
    Odrv4 I__3267 (
            .O(N__26018),
            .I(n2615));
    InMux I__3266 (
            .O(N__26013),
            .I(N__26010));
    LocalMux I__3265 (
            .O(N__26010),
            .I(N__26007));
    Span4Mux_s3_h I__3264 (
            .O(N__26007),
            .I(N__26004));
    Odrv4 I__3263 (
            .O(N__26004),
            .I(n2682));
    InMux I__3262 (
            .O(N__26001),
            .I(n12766));
    InMux I__3261 (
            .O(N__25998),
            .I(N__25991));
    InMux I__3260 (
            .O(N__25997),
            .I(N__25991));
    InMux I__3259 (
            .O(N__25996),
            .I(N__25988));
    LocalMux I__3258 (
            .O(N__25991),
            .I(N__25985));
    LocalMux I__3257 (
            .O(N__25988),
            .I(n2614));
    Odrv4 I__3256 (
            .O(N__25985),
            .I(n2614));
    InMux I__3255 (
            .O(N__25980),
            .I(N__25977));
    LocalMux I__3254 (
            .O(N__25977),
            .I(n2681));
    InMux I__3253 (
            .O(N__25974),
            .I(n12767));
    InMux I__3252 (
            .O(N__25971),
            .I(N__25967));
    CascadeMux I__3251 (
            .O(N__25970),
            .I(N__25964));
    LocalMux I__3250 (
            .O(N__25967),
            .I(N__25961));
    InMux I__3249 (
            .O(N__25964),
            .I(N__25958));
    Odrv4 I__3248 (
            .O(N__25961),
            .I(n2629));
    LocalMux I__3247 (
            .O(N__25958),
            .I(n2629));
    InMux I__3246 (
            .O(N__25953),
            .I(N__25950));
    LocalMux I__3245 (
            .O(N__25950),
            .I(N__25947));
    Odrv4 I__3244 (
            .O(N__25947),
            .I(n2696));
    InMux I__3243 (
            .O(N__25944),
            .I(n12752));
    CascadeMux I__3242 (
            .O(N__25941),
            .I(N__25937));
    InMux I__3241 (
            .O(N__25940),
            .I(N__25934));
    InMux I__3240 (
            .O(N__25937),
            .I(N__25931));
    LocalMux I__3239 (
            .O(N__25934),
            .I(N__25928));
    LocalMux I__3238 (
            .O(N__25931),
            .I(N__25925));
    Odrv4 I__3237 (
            .O(N__25928),
            .I(n2628));
    Odrv4 I__3236 (
            .O(N__25925),
            .I(n2628));
    InMux I__3235 (
            .O(N__25920),
            .I(N__25917));
    LocalMux I__3234 (
            .O(N__25917),
            .I(N__25914));
    Odrv4 I__3233 (
            .O(N__25914),
            .I(n2695));
    InMux I__3232 (
            .O(N__25911),
            .I(n12753));
    InMux I__3231 (
            .O(N__25908),
            .I(N__25905));
    LocalMux I__3230 (
            .O(N__25905),
            .I(N__25901));
    CascadeMux I__3229 (
            .O(N__25904),
            .I(N__25898));
    Span4Mux_h I__3228 (
            .O(N__25901),
            .I(N__25895));
    InMux I__3227 (
            .O(N__25898),
            .I(N__25892));
    Span4Mux_v I__3226 (
            .O(N__25895),
            .I(N__25887));
    LocalMux I__3225 (
            .O(N__25892),
            .I(N__25887));
    Odrv4 I__3224 (
            .O(N__25887),
            .I(n2627));
    CascadeMux I__3223 (
            .O(N__25884),
            .I(N__25881));
    InMux I__3222 (
            .O(N__25881),
            .I(N__25878));
    LocalMux I__3221 (
            .O(N__25878),
            .I(N__25875));
    Span4Mux_v I__3220 (
            .O(N__25875),
            .I(N__25872));
    Odrv4 I__3219 (
            .O(N__25872),
            .I(n2694));
    InMux I__3218 (
            .O(N__25869),
            .I(n12754));
    CascadeMux I__3217 (
            .O(N__25866),
            .I(N__25862));
    InMux I__3216 (
            .O(N__25865),
            .I(N__25859));
    InMux I__3215 (
            .O(N__25862),
            .I(N__25855));
    LocalMux I__3214 (
            .O(N__25859),
            .I(N__25852));
    InMux I__3213 (
            .O(N__25858),
            .I(N__25849));
    LocalMux I__3212 (
            .O(N__25855),
            .I(n2626));
    Odrv12 I__3211 (
            .O(N__25852),
            .I(n2626));
    LocalMux I__3210 (
            .O(N__25849),
            .I(n2626));
    InMux I__3209 (
            .O(N__25842),
            .I(N__25839));
    LocalMux I__3208 (
            .O(N__25839),
            .I(n2693));
    InMux I__3207 (
            .O(N__25836),
            .I(bfn_4_22_0_));
    InMux I__3206 (
            .O(N__25833),
            .I(N__25830));
    LocalMux I__3205 (
            .O(N__25830),
            .I(N__25825));
    InMux I__3204 (
            .O(N__25829),
            .I(N__25822));
    InMux I__3203 (
            .O(N__25828),
            .I(N__25819));
    Odrv4 I__3202 (
            .O(N__25825),
            .I(n2625));
    LocalMux I__3201 (
            .O(N__25822),
            .I(n2625));
    LocalMux I__3200 (
            .O(N__25819),
            .I(n2625));
    InMux I__3199 (
            .O(N__25812),
            .I(N__25809));
    LocalMux I__3198 (
            .O(N__25809),
            .I(n2692));
    InMux I__3197 (
            .O(N__25806),
            .I(n12756));
    InMux I__3196 (
            .O(N__25803),
            .I(N__25800));
    LocalMux I__3195 (
            .O(N__25800),
            .I(N__25797));
    Span4Mux_h I__3194 (
            .O(N__25797),
            .I(N__25793));
    InMux I__3193 (
            .O(N__25796),
            .I(N__25790));
    Odrv4 I__3192 (
            .O(N__25793),
            .I(n2624));
    LocalMux I__3191 (
            .O(N__25790),
            .I(n2624));
    CascadeMux I__3190 (
            .O(N__25785),
            .I(N__25782));
    InMux I__3189 (
            .O(N__25782),
            .I(N__25779));
    LocalMux I__3188 (
            .O(N__25779),
            .I(N__25776));
    Odrv4 I__3187 (
            .O(N__25776),
            .I(n2691));
    InMux I__3186 (
            .O(N__25773),
            .I(n12757));
    CascadeMux I__3185 (
            .O(N__25770),
            .I(N__25767));
    InMux I__3184 (
            .O(N__25767),
            .I(N__25764));
    LocalMux I__3183 (
            .O(N__25764),
            .I(N__25759));
    InMux I__3182 (
            .O(N__25763),
            .I(N__25756));
    InMux I__3181 (
            .O(N__25762),
            .I(N__25753));
    Odrv12 I__3180 (
            .O(N__25759),
            .I(n2623));
    LocalMux I__3179 (
            .O(N__25756),
            .I(n2623));
    LocalMux I__3178 (
            .O(N__25753),
            .I(n2623));
    InMux I__3177 (
            .O(N__25746),
            .I(N__25743));
    LocalMux I__3176 (
            .O(N__25743),
            .I(N__25740));
    Odrv4 I__3175 (
            .O(N__25740),
            .I(n2690));
    InMux I__3174 (
            .O(N__25737),
            .I(n12758));
    InMux I__3173 (
            .O(N__25734),
            .I(N__25731));
    LocalMux I__3172 (
            .O(N__25731),
            .I(N__25726));
    InMux I__3171 (
            .O(N__25730),
            .I(N__25723));
    InMux I__3170 (
            .O(N__25729),
            .I(N__25720));
    Odrv12 I__3169 (
            .O(N__25726),
            .I(n2622));
    LocalMux I__3168 (
            .O(N__25723),
            .I(n2622));
    LocalMux I__3167 (
            .O(N__25720),
            .I(n2622));
    InMux I__3166 (
            .O(N__25713),
            .I(N__25710));
    LocalMux I__3165 (
            .O(N__25710),
            .I(N__25707));
    Odrv4 I__3164 (
            .O(N__25707),
            .I(n2689));
    InMux I__3163 (
            .O(N__25704),
            .I(n12759));
    InMux I__3162 (
            .O(N__25701),
            .I(N__25698));
    LocalMux I__3161 (
            .O(N__25698),
            .I(N__25695));
    Span4Mux_h I__3160 (
            .O(N__25695),
            .I(N__25692));
    Odrv4 I__3159 (
            .O(N__25692),
            .I(n2492));
    CascadeMux I__3158 (
            .O(N__25689),
            .I(N__25686));
    InMux I__3157 (
            .O(N__25686),
            .I(N__25682));
    CascadeMux I__3156 (
            .O(N__25685),
            .I(N__25679));
    LocalMux I__3155 (
            .O(N__25682),
            .I(N__25676));
    InMux I__3154 (
            .O(N__25679),
            .I(N__25673));
    Span4Mux_v I__3153 (
            .O(N__25676),
            .I(N__25670));
    LocalMux I__3152 (
            .O(N__25673),
            .I(n2425));
    Odrv4 I__3151 (
            .O(N__25670),
            .I(n2425));
    CascadeMux I__3150 (
            .O(N__25665),
            .I(N__25662));
    InMux I__3149 (
            .O(N__25662),
            .I(N__25659));
    LocalMux I__3148 (
            .O(N__25659),
            .I(N__25656));
    Span4Mux_v I__3147 (
            .O(N__25656),
            .I(N__25651));
    InMux I__3146 (
            .O(N__25655),
            .I(N__25646));
    InMux I__3145 (
            .O(N__25654),
            .I(N__25646));
    Odrv4 I__3144 (
            .O(N__25651),
            .I(n2524));
    LocalMux I__3143 (
            .O(N__25646),
            .I(n2524));
    CascadeMux I__3142 (
            .O(N__25641),
            .I(N__25638));
    InMux I__3141 (
            .O(N__25638),
            .I(N__25633));
    InMux I__3140 (
            .O(N__25637),
            .I(N__25628));
    InMux I__3139 (
            .O(N__25636),
            .I(N__25628));
    LocalMux I__3138 (
            .O(N__25633),
            .I(n2318));
    LocalMux I__3137 (
            .O(N__25628),
            .I(n2318));
    CascadeMux I__3136 (
            .O(N__25623),
            .I(N__25620));
    InMux I__3135 (
            .O(N__25620),
            .I(N__25616));
    InMux I__3134 (
            .O(N__25619),
            .I(N__25612));
    LocalMux I__3133 (
            .O(N__25616),
            .I(N__25609));
    InMux I__3132 (
            .O(N__25615),
            .I(N__25606));
    LocalMux I__3131 (
            .O(N__25612),
            .I(n2320));
    Odrv4 I__3130 (
            .O(N__25609),
            .I(n2320));
    LocalMux I__3129 (
            .O(N__25606),
            .I(n2320));
    CascadeMux I__3128 (
            .O(N__25599),
            .I(N__25596));
    InMux I__3127 (
            .O(N__25596),
            .I(N__25593));
    LocalMux I__3126 (
            .O(N__25593),
            .I(N__25589));
    InMux I__3125 (
            .O(N__25592),
            .I(N__25586));
    Span4Mux_v I__3124 (
            .O(N__25589),
            .I(N__25582));
    LocalMux I__3123 (
            .O(N__25586),
            .I(N__25579));
    InMux I__3122 (
            .O(N__25585),
            .I(N__25576));
    Odrv4 I__3121 (
            .O(N__25582),
            .I(n2319));
    Odrv4 I__3120 (
            .O(N__25579),
            .I(n2319));
    LocalMux I__3119 (
            .O(N__25576),
            .I(n2319));
    InMux I__3118 (
            .O(N__25569),
            .I(bfn_4_21_0_));
    InMux I__3117 (
            .O(N__25566),
            .I(N__25563));
    LocalMux I__3116 (
            .O(N__25563),
            .I(N__25560));
    Odrv4 I__3115 (
            .O(N__25560),
            .I(n2700));
    InMux I__3114 (
            .O(N__25557),
            .I(n12748));
    InMux I__3113 (
            .O(N__25554),
            .I(n12749));
    InMux I__3112 (
            .O(N__25551),
            .I(n12750));
    InMux I__3111 (
            .O(N__25548),
            .I(n12751));
    InMux I__3110 (
            .O(N__25545),
            .I(n12699));
    InMux I__3109 (
            .O(N__25542),
            .I(N__25539));
    LocalMux I__3108 (
            .O(N__25539),
            .I(n2382));
    InMux I__3107 (
            .O(N__25536),
            .I(n12700));
    InMux I__3106 (
            .O(N__25533),
            .I(N__25530));
    LocalMux I__3105 (
            .O(N__25530),
            .I(n2381));
    InMux I__3104 (
            .O(N__25527),
            .I(n12701));
    InMux I__3103 (
            .O(N__25524),
            .I(n12702));
    CascadeMux I__3102 (
            .O(N__25521),
            .I(N__25518));
    InMux I__3101 (
            .O(N__25518),
            .I(N__25515));
    LocalMux I__3100 (
            .O(N__25515),
            .I(N__25511));
    InMux I__3099 (
            .O(N__25514),
            .I(N__25508));
    Odrv4 I__3098 (
            .O(N__25511),
            .I(n2412));
    LocalMux I__3097 (
            .O(N__25508),
            .I(n2412));
    InMux I__3096 (
            .O(N__25503),
            .I(N__25498));
    InMux I__3095 (
            .O(N__25502),
            .I(N__25495));
    InMux I__3094 (
            .O(N__25501),
            .I(N__25492));
    LocalMux I__3093 (
            .O(N__25498),
            .I(n2314_adj_622));
    LocalMux I__3092 (
            .O(N__25495),
            .I(n2314_adj_622));
    LocalMux I__3091 (
            .O(N__25492),
            .I(n2314_adj_622));
    CascadeMux I__3090 (
            .O(N__25485),
            .I(N__25481));
    CascadeMux I__3089 (
            .O(N__25484),
            .I(N__25478));
    InMux I__3088 (
            .O(N__25481),
            .I(N__25475));
    InMux I__3087 (
            .O(N__25478),
            .I(N__25472));
    LocalMux I__3086 (
            .O(N__25475),
            .I(N__25467));
    LocalMux I__3085 (
            .O(N__25472),
            .I(N__25467));
    Odrv4 I__3084 (
            .O(N__25467),
            .I(n2327));
    CascadeMux I__3083 (
            .O(N__25464),
            .I(n2327_cascade_));
    CascadeMux I__3082 (
            .O(N__25461),
            .I(N__25457));
    InMux I__3081 (
            .O(N__25460),
            .I(N__25453));
    InMux I__3080 (
            .O(N__25457),
            .I(N__25450));
    InMux I__3079 (
            .O(N__25456),
            .I(N__25447));
    LocalMux I__3078 (
            .O(N__25453),
            .I(n2326));
    LocalMux I__3077 (
            .O(N__25450),
            .I(n2326));
    LocalMux I__3076 (
            .O(N__25447),
            .I(n2326));
    InMux I__3075 (
            .O(N__25440),
            .I(N__25437));
    LocalMux I__3074 (
            .O(N__25437),
            .I(n14440));
    InMux I__3073 (
            .O(N__25434),
            .I(N__25431));
    LocalMux I__3072 (
            .O(N__25431),
            .I(n2391));
    InMux I__3071 (
            .O(N__25428),
            .I(n12691));
    InMux I__3070 (
            .O(N__25425),
            .I(N__25422));
    LocalMux I__3069 (
            .O(N__25422),
            .I(N__25419));
    Odrv4 I__3068 (
            .O(N__25419),
            .I(n2390));
    InMux I__3067 (
            .O(N__25416),
            .I(n12692));
    InMux I__3066 (
            .O(N__25413),
            .I(N__25410));
    LocalMux I__3065 (
            .O(N__25410),
            .I(n2389));
    InMux I__3064 (
            .O(N__25407),
            .I(n12693));
    InMux I__3063 (
            .O(N__25404),
            .I(N__25401));
    LocalMux I__3062 (
            .O(N__25401),
            .I(n2388));
    InMux I__3061 (
            .O(N__25398),
            .I(n12694));
    InMux I__3060 (
            .O(N__25395),
            .I(N__25392));
    LocalMux I__3059 (
            .O(N__25392),
            .I(n2387));
    InMux I__3058 (
            .O(N__25389),
            .I(n12695));
    InMux I__3057 (
            .O(N__25386),
            .I(N__25383));
    LocalMux I__3056 (
            .O(N__25383),
            .I(N__25380));
    Odrv4 I__3055 (
            .O(N__25380),
            .I(n2386));
    InMux I__3054 (
            .O(N__25377),
            .I(n12696));
    InMux I__3053 (
            .O(N__25374),
            .I(N__25371));
    LocalMux I__3052 (
            .O(N__25371),
            .I(n2385));
    InMux I__3051 (
            .O(N__25368),
            .I(bfn_4_19_0_));
    InMux I__3050 (
            .O(N__25365),
            .I(N__25362));
    LocalMux I__3049 (
            .O(N__25362),
            .I(N__25359));
    Odrv4 I__3048 (
            .O(N__25359),
            .I(n2384));
    InMux I__3047 (
            .O(N__25356),
            .I(n12698));
    InMux I__3046 (
            .O(N__25353),
            .I(N__25350));
    LocalMux I__3045 (
            .O(N__25350),
            .I(n2383));
    InMux I__3044 (
            .O(N__25347),
            .I(N__25344));
    LocalMux I__3043 (
            .O(N__25344),
            .I(N__25341));
    Span4Mux_s3_h I__3042 (
            .O(N__25341),
            .I(N__25338));
    Odrv4 I__3041 (
            .O(N__25338),
            .I(n2399));
    InMux I__3040 (
            .O(N__25335),
            .I(n12683));
    InMux I__3039 (
            .O(N__25332),
            .I(N__25329));
    LocalMux I__3038 (
            .O(N__25329),
            .I(N__25326));
    Span4Mux_s3_h I__3037 (
            .O(N__25326),
            .I(N__25323));
    Odrv4 I__3036 (
            .O(N__25323),
            .I(n2398));
    InMux I__3035 (
            .O(N__25320),
            .I(n12684));
    CascadeMux I__3034 (
            .O(N__25317),
            .I(N__25314));
    InMux I__3033 (
            .O(N__25314),
            .I(N__25311));
    LocalMux I__3032 (
            .O(N__25311),
            .I(n2397));
    InMux I__3031 (
            .O(N__25308),
            .I(n12685));
    CascadeMux I__3030 (
            .O(N__25305),
            .I(N__25301));
    CascadeMux I__3029 (
            .O(N__25304),
            .I(N__25298));
    InMux I__3028 (
            .O(N__25301),
            .I(N__25294));
    InMux I__3027 (
            .O(N__25298),
            .I(N__25291));
    InMux I__3026 (
            .O(N__25297),
            .I(N__25288));
    LocalMux I__3025 (
            .O(N__25294),
            .I(N__25285));
    LocalMux I__3024 (
            .O(N__25291),
            .I(n2329));
    LocalMux I__3023 (
            .O(N__25288),
            .I(n2329));
    Odrv4 I__3022 (
            .O(N__25285),
            .I(n2329));
    InMux I__3021 (
            .O(N__25278),
            .I(N__25275));
    LocalMux I__3020 (
            .O(N__25275),
            .I(N__25272));
    Span4Mux_s3_h I__3019 (
            .O(N__25272),
            .I(N__25269));
    Odrv4 I__3018 (
            .O(N__25269),
            .I(n2396));
    InMux I__3017 (
            .O(N__25266),
            .I(n12686));
    CascadeMux I__3016 (
            .O(N__25263),
            .I(N__25259));
    InMux I__3015 (
            .O(N__25262),
            .I(N__25256));
    InMux I__3014 (
            .O(N__25259),
            .I(N__25253));
    LocalMux I__3013 (
            .O(N__25256),
            .I(N__25248));
    LocalMux I__3012 (
            .O(N__25253),
            .I(N__25248));
    Odrv4 I__3011 (
            .O(N__25248),
            .I(n2328));
    InMux I__3010 (
            .O(N__25245),
            .I(N__25242));
    LocalMux I__3009 (
            .O(N__25242),
            .I(n2395));
    InMux I__3008 (
            .O(N__25239),
            .I(n12687));
    InMux I__3007 (
            .O(N__25236),
            .I(N__25233));
    LocalMux I__3006 (
            .O(N__25233),
            .I(n2394));
    InMux I__3005 (
            .O(N__25230),
            .I(n12688));
    CascadeMux I__3004 (
            .O(N__25227),
            .I(N__25224));
    InMux I__3003 (
            .O(N__25224),
            .I(N__25221));
    LocalMux I__3002 (
            .O(N__25221),
            .I(n2393));
    InMux I__3001 (
            .O(N__25218),
            .I(bfn_4_18_0_));
    CascadeMux I__3000 (
            .O(N__25215),
            .I(N__25212));
    InMux I__2999 (
            .O(N__25212),
            .I(N__25209));
    LocalMux I__2998 (
            .O(N__25209),
            .I(N__25206));
    Odrv4 I__2997 (
            .O(N__25206),
            .I(n2392));
    InMux I__2996 (
            .O(N__25203),
            .I(n12690));
    InMux I__2995 (
            .O(N__25200),
            .I(bfn_3_32_0_));
    InMux I__2994 (
            .O(N__25197),
            .I(n12874));
    InMux I__2993 (
            .O(N__25194),
            .I(n12875));
    InMux I__2992 (
            .O(N__25191),
            .I(n12876));
    InMux I__2991 (
            .O(N__25188),
            .I(n12877));
    InMux I__2990 (
            .O(N__25185),
            .I(N__25182));
    LocalMux I__2989 (
            .O(N__25182),
            .I(N__25178));
    InMux I__2988 (
            .O(N__25181),
            .I(N__25175));
    Span4Mux_s1_v I__2987 (
            .O(N__25178),
            .I(N__25172));
    LocalMux I__2986 (
            .O(N__25175),
            .I(\debounce.cnt_reg_6 ));
    Odrv4 I__2985 (
            .O(N__25172),
            .I(\debounce.cnt_reg_6 ));
    InMux I__2984 (
            .O(N__25167),
            .I(N__25164));
    LocalMux I__2983 (
            .O(N__25164),
            .I(\debounce.n16 ));
    CascadeMux I__2982 (
            .O(N__25161),
            .I(N__25158));
    InMux I__2981 (
            .O(N__25158),
            .I(N__25155));
    LocalMux I__2980 (
            .O(N__25155),
            .I(N__25151));
    InMux I__2979 (
            .O(N__25154),
            .I(N__25148));
    Span4Mux_s1_v I__2978 (
            .O(N__25151),
            .I(N__25145));
    LocalMux I__2977 (
            .O(N__25148),
            .I(\debounce.cnt_reg_3 ));
    Odrv4 I__2976 (
            .O(N__25145),
            .I(\debounce.cnt_reg_3 ));
    InMux I__2975 (
            .O(N__25140),
            .I(N__25137));
    LocalMux I__2974 (
            .O(N__25137),
            .I(\debounce.n17 ));
    InMux I__2973 (
            .O(N__25134),
            .I(N__25131));
    LocalMux I__2972 (
            .O(N__25131),
            .I(N__25128));
    Odrv4 I__2971 (
            .O(N__25128),
            .I(n2401));
    InMux I__2970 (
            .O(N__25125),
            .I(bfn_4_17_0_));
    InMux I__2969 (
            .O(N__25122),
            .I(N__25119));
    LocalMux I__2968 (
            .O(N__25119),
            .I(N__25116));
    Odrv4 I__2967 (
            .O(N__25116),
            .I(n2400));
    InMux I__2966 (
            .O(N__25113),
            .I(n12682));
    CascadeMux I__2965 (
            .O(N__25110),
            .I(N__25107));
    InMux I__2964 (
            .O(N__25107),
            .I(N__25104));
    LocalMux I__2963 (
            .O(N__25104),
            .I(N__25101));
    Odrv4 I__2962 (
            .O(N__25101),
            .I(n3086));
    InMux I__2961 (
            .O(N__25098),
            .I(n12864));
    InMux I__2960 (
            .O(N__25095),
            .I(bfn_3_31_0_));
    InMux I__2959 (
            .O(N__25092),
            .I(n12866));
    InMux I__2958 (
            .O(N__25089),
            .I(n12867));
    InMux I__2957 (
            .O(N__25086),
            .I(n12868));
    InMux I__2956 (
            .O(N__25083),
            .I(n12869));
    InMux I__2955 (
            .O(N__25080),
            .I(n12870));
    InMux I__2954 (
            .O(N__25077),
            .I(n12871));
    InMux I__2953 (
            .O(N__25074),
            .I(n12872));
    InMux I__2952 (
            .O(N__25071),
            .I(n12855));
    InMux I__2951 (
            .O(N__25068),
            .I(n12856));
    InMux I__2950 (
            .O(N__25065),
            .I(bfn_3_30_0_));
    InMux I__2949 (
            .O(N__25062),
            .I(n12858));
    InMux I__2948 (
            .O(N__25059),
            .I(n12859));
    InMux I__2947 (
            .O(N__25056),
            .I(n12860));
    InMux I__2946 (
            .O(N__25053),
            .I(n12861));
    InMux I__2945 (
            .O(N__25050),
            .I(n12862));
    InMux I__2944 (
            .O(N__25047),
            .I(n12863));
    InMux I__2943 (
            .O(N__25044),
            .I(N__25041));
    LocalMux I__2942 (
            .O(N__25041),
            .I(N__25038));
    Span4Mux_h I__2941 (
            .O(N__25038),
            .I(N__25035));
    Odrv4 I__2940 (
            .O(N__25035),
            .I(n2893));
    CascadeMux I__2939 (
            .O(N__25032),
            .I(N__25028));
    CascadeMux I__2938 (
            .O(N__25031),
            .I(N__25025));
    InMux I__2937 (
            .O(N__25028),
            .I(N__25021));
    InMux I__2936 (
            .O(N__25025),
            .I(N__25018));
    InMux I__2935 (
            .O(N__25024),
            .I(N__25015));
    LocalMux I__2934 (
            .O(N__25021),
            .I(n2826));
    LocalMux I__2933 (
            .O(N__25018),
            .I(n2826));
    LocalMux I__2932 (
            .O(N__25015),
            .I(n2826));
    CascadeMux I__2931 (
            .O(N__25008),
            .I(N__25005));
    InMux I__2930 (
            .O(N__25005),
            .I(N__25002));
    LocalMux I__2929 (
            .O(N__25002),
            .I(N__24999));
    Odrv4 I__2928 (
            .O(N__24999),
            .I(n2882));
    InMux I__2927 (
            .O(N__24996),
            .I(N__24993));
    LocalMux I__2926 (
            .O(N__24993),
            .I(N__24989));
    InMux I__2925 (
            .O(N__24992),
            .I(N__24986));
    Span4Mux_h I__2924 (
            .O(N__24989),
            .I(N__24980));
    LocalMux I__2923 (
            .O(N__24986),
            .I(N__24980));
    InMux I__2922 (
            .O(N__24985),
            .I(N__24977));
    Odrv4 I__2921 (
            .O(N__24980),
            .I(n2815));
    LocalMux I__2920 (
            .O(N__24977),
            .I(n2815));
    InMux I__2919 (
            .O(N__24972),
            .I(N__24967));
    InMux I__2918 (
            .O(N__24971),
            .I(N__24964));
    InMux I__2917 (
            .O(N__24970),
            .I(N__24961));
    LocalMux I__2916 (
            .O(N__24967),
            .I(n2813));
    LocalMux I__2915 (
            .O(N__24964),
            .I(n2813));
    LocalMux I__2914 (
            .O(N__24961),
            .I(n2813));
    CascadeMux I__2913 (
            .O(N__24954),
            .I(N__24951));
    InMux I__2912 (
            .O(N__24951),
            .I(N__24948));
    LocalMux I__2911 (
            .O(N__24948),
            .I(N__24945));
    Span4Mux_h I__2910 (
            .O(N__24945),
            .I(N__24942));
    Odrv4 I__2909 (
            .O(N__24942),
            .I(n2880));
    InMux I__2908 (
            .O(N__24939),
            .I(bfn_3_29_0_));
    InMux I__2907 (
            .O(N__24936),
            .I(n12850));
    InMux I__2906 (
            .O(N__24933),
            .I(n12851));
    InMux I__2905 (
            .O(N__24930),
            .I(n12852));
    InMux I__2904 (
            .O(N__24927),
            .I(n12853));
    InMux I__2903 (
            .O(N__24924),
            .I(n12854));
    InMux I__2902 (
            .O(N__24921),
            .I(N__24918));
    LocalMux I__2901 (
            .O(N__24918),
            .I(n2777));
    CascadeMux I__2900 (
            .O(N__24915),
            .I(N__24912));
    InMux I__2899 (
            .O(N__24912),
            .I(N__24907));
    InMux I__2898 (
            .O(N__24911),
            .I(N__24902));
    InMux I__2897 (
            .O(N__24910),
            .I(N__24902));
    LocalMux I__2896 (
            .O(N__24907),
            .I(n2710));
    LocalMux I__2895 (
            .O(N__24902),
            .I(n2710));
    InMux I__2894 (
            .O(N__24897),
            .I(N__24893));
    InMux I__2893 (
            .O(N__24896),
            .I(N__24890));
    LocalMux I__2892 (
            .O(N__24893),
            .I(N__24887));
    LocalMux I__2891 (
            .O(N__24890),
            .I(N__24884));
    Span4Mux_v I__2890 (
            .O(N__24887),
            .I(N__24881));
    Span4Mux_s2_h I__2889 (
            .O(N__24884),
            .I(N__24878));
    Odrv4 I__2888 (
            .O(N__24881),
            .I(n2809));
    Odrv4 I__2887 (
            .O(N__24878),
            .I(n2809));
    InMux I__2886 (
            .O(N__24873),
            .I(N__24868));
    InMux I__2885 (
            .O(N__24872),
            .I(N__24865));
    InMux I__2884 (
            .O(N__24871),
            .I(N__24862));
    LocalMux I__2883 (
            .O(N__24868),
            .I(N__24857));
    LocalMux I__2882 (
            .O(N__24865),
            .I(N__24857));
    LocalMux I__2881 (
            .O(N__24862),
            .I(N__24854));
    Odrv4 I__2880 (
            .O(N__24857),
            .I(n2810));
    Odrv4 I__2879 (
            .O(N__24854),
            .I(n2810));
    InMux I__2878 (
            .O(N__24849),
            .I(N__24846));
    LocalMux I__2877 (
            .O(N__24846),
            .I(N__24843));
    Span4Mux_v I__2876 (
            .O(N__24843),
            .I(N__24839));
    InMux I__2875 (
            .O(N__24842),
            .I(N__24836));
    Odrv4 I__2874 (
            .O(N__24839),
            .I(n2808));
    LocalMux I__2873 (
            .O(N__24836),
            .I(n2808));
    CascadeMux I__2872 (
            .O(N__24831),
            .I(n2809_cascade_));
    InMux I__2871 (
            .O(N__24828),
            .I(N__24825));
    LocalMux I__2870 (
            .O(N__24825),
            .I(n14714));
    CascadeMux I__2869 (
            .O(N__24822),
            .I(N__24819));
    InMux I__2868 (
            .O(N__24819),
            .I(N__24815));
    InMux I__2867 (
            .O(N__24818),
            .I(N__24812));
    LocalMux I__2866 (
            .O(N__24815),
            .I(N__24809));
    LocalMux I__2865 (
            .O(N__24812),
            .I(n2823));
    Odrv4 I__2864 (
            .O(N__24809),
            .I(n2823));
    CascadeMux I__2863 (
            .O(N__24804),
            .I(n2841_cascade_));
    InMux I__2862 (
            .O(N__24801),
            .I(N__24798));
    LocalMux I__2861 (
            .O(N__24798),
            .I(N__24795));
    Odrv4 I__2860 (
            .O(N__24795),
            .I(n2890));
    CascadeMux I__2859 (
            .O(N__24792),
            .I(N__24789));
    InMux I__2858 (
            .O(N__24789),
            .I(N__24785));
    InMux I__2857 (
            .O(N__24788),
            .I(N__24781));
    LocalMux I__2856 (
            .O(N__24785),
            .I(N__24778));
    InMux I__2855 (
            .O(N__24784),
            .I(N__24775));
    LocalMux I__2854 (
            .O(N__24781),
            .I(n2920));
    Odrv4 I__2853 (
            .O(N__24778),
            .I(n2920));
    LocalMux I__2852 (
            .O(N__24775),
            .I(n2920));
    CascadeMux I__2851 (
            .O(N__24768),
            .I(N__24765));
    InMux I__2850 (
            .O(N__24765),
            .I(N__24762));
    LocalMux I__2849 (
            .O(N__24762),
            .I(N__24759));
    Odrv4 I__2848 (
            .O(N__24759),
            .I(n2987));
    InMux I__2847 (
            .O(N__24756),
            .I(N__24753));
    LocalMux I__2846 (
            .O(N__24753),
            .I(N__24750));
    Span4Mux_v I__2845 (
            .O(N__24750),
            .I(N__24747));
    Odrv4 I__2844 (
            .O(N__24747),
            .I(n2898));
    CascadeMux I__2843 (
            .O(N__24744),
            .I(N__24741));
    InMux I__2842 (
            .O(N__24741),
            .I(N__24738));
    LocalMux I__2841 (
            .O(N__24738),
            .I(N__24734));
    CascadeMux I__2840 (
            .O(N__24737),
            .I(N__24731));
    Span4Mux_h I__2839 (
            .O(N__24734),
            .I(N__24727));
    InMux I__2838 (
            .O(N__24731),
            .I(N__24724));
    InMux I__2837 (
            .O(N__24730),
            .I(N__24721));
    Odrv4 I__2836 (
            .O(N__24727),
            .I(n2831));
    LocalMux I__2835 (
            .O(N__24724),
            .I(n2831));
    LocalMux I__2834 (
            .O(N__24721),
            .I(n2831));
    InMux I__2833 (
            .O(N__24714),
            .I(N__24711));
    LocalMux I__2832 (
            .O(N__24711),
            .I(N__24708));
    Odrv4 I__2831 (
            .O(N__24708),
            .I(n2879));
    InMux I__2830 (
            .O(N__24705),
            .I(N__24700));
    InMux I__2829 (
            .O(N__24704),
            .I(N__24697));
    InMux I__2828 (
            .O(N__24703),
            .I(N__24694));
    LocalMux I__2827 (
            .O(N__24700),
            .I(n2812));
    LocalMux I__2826 (
            .O(N__24697),
            .I(n2812));
    LocalMux I__2825 (
            .O(N__24694),
            .I(n2812));
    CascadeMux I__2824 (
            .O(N__24687),
            .I(n2911_cascade_));
    InMux I__2823 (
            .O(N__24684),
            .I(N__24681));
    LocalMux I__2822 (
            .O(N__24681),
            .I(N__24677));
    CascadeMux I__2821 (
            .O(N__24680),
            .I(N__24674));
    Span4Mux_v I__2820 (
            .O(N__24677),
            .I(N__24671));
    InMux I__2819 (
            .O(N__24674),
            .I(N__24668));
    Odrv4 I__2818 (
            .O(N__24671),
            .I(n2829));
    LocalMux I__2817 (
            .O(N__24668),
            .I(n2829));
    InMux I__2816 (
            .O(N__24663),
            .I(N__24660));
    LocalMux I__2815 (
            .O(N__24660),
            .I(N__24657));
    Span4Mux_h I__2814 (
            .O(N__24657),
            .I(N__24654));
    Odrv4 I__2813 (
            .O(N__24654),
            .I(n2896));
    InMux I__2812 (
            .O(N__24651),
            .I(N__24646));
    CascadeMux I__2811 (
            .O(N__24650),
            .I(N__24643));
    InMux I__2810 (
            .O(N__24649),
            .I(N__24640));
    LocalMux I__2809 (
            .O(N__24646),
            .I(N__24637));
    InMux I__2808 (
            .O(N__24643),
            .I(N__24634));
    LocalMux I__2807 (
            .O(N__24640),
            .I(N__24631));
    Odrv4 I__2806 (
            .O(N__24637),
            .I(n2725));
    LocalMux I__2805 (
            .O(N__24634),
            .I(n2725));
    Odrv4 I__2804 (
            .O(N__24631),
            .I(n2725));
    InMux I__2803 (
            .O(N__24624),
            .I(N__24621));
    LocalMux I__2802 (
            .O(N__24621),
            .I(N__24618));
    Span4Mux_h I__2801 (
            .O(N__24618),
            .I(N__24615));
    Odrv4 I__2800 (
            .O(N__24615),
            .I(n2792));
    InMux I__2799 (
            .O(N__24612),
            .I(N__24608));
    InMux I__2798 (
            .O(N__24611),
            .I(N__24605));
    LocalMux I__2797 (
            .O(N__24608),
            .I(n2721));
    LocalMux I__2796 (
            .O(N__24605),
            .I(n2721));
    InMux I__2795 (
            .O(N__24600),
            .I(N__24597));
    LocalMux I__2794 (
            .O(N__24597),
            .I(N__24594));
    Odrv4 I__2793 (
            .O(N__24594),
            .I(n2788));
    CascadeMux I__2792 (
            .O(N__24591),
            .I(N__24588));
    InMux I__2791 (
            .O(N__24588),
            .I(N__24585));
    LocalMux I__2790 (
            .O(N__24585),
            .I(N__24582));
    Odrv4 I__2789 (
            .O(N__24582),
            .I(n2793));
    CascadeMux I__2788 (
            .O(N__24579),
            .I(N__24576));
    InMux I__2787 (
            .O(N__24576),
            .I(N__24573));
    LocalMux I__2786 (
            .O(N__24573),
            .I(N__24570));
    Odrv4 I__2785 (
            .O(N__24570),
            .I(n2889));
    CascadeMux I__2784 (
            .O(N__24567),
            .I(n2921_cascade_));
    CascadeMux I__2783 (
            .O(N__24564),
            .I(N__24561));
    InMux I__2782 (
            .O(N__24561),
            .I(N__24558));
    LocalMux I__2781 (
            .O(N__24558),
            .I(N__24555));
    Odrv4 I__2780 (
            .O(N__24555),
            .I(n2888));
    CascadeMux I__2779 (
            .O(N__24552),
            .I(N__24549));
    InMux I__2778 (
            .O(N__24549),
            .I(N__24546));
    LocalMux I__2777 (
            .O(N__24546),
            .I(N__24543));
    Odrv4 I__2776 (
            .O(N__24543),
            .I(n2791));
    CascadeMux I__2775 (
            .O(N__24540),
            .I(N__24537));
    InMux I__2774 (
            .O(N__24537),
            .I(N__24532));
    InMux I__2773 (
            .O(N__24536),
            .I(N__24527));
    InMux I__2772 (
            .O(N__24535),
            .I(N__24527));
    LocalMux I__2771 (
            .O(N__24532),
            .I(n2822));
    LocalMux I__2770 (
            .O(N__24527),
            .I(n2822));
    CascadeMux I__2769 (
            .O(N__24522),
            .I(n2823_cascade_));
    CascadeMux I__2768 (
            .O(N__24519),
            .I(N__24516));
    InMux I__2767 (
            .O(N__24516),
            .I(N__24511));
    InMux I__2766 (
            .O(N__24515),
            .I(N__24506));
    InMux I__2765 (
            .O(N__24514),
            .I(N__24506));
    LocalMux I__2764 (
            .O(N__24511),
            .I(n2821));
    LocalMux I__2763 (
            .O(N__24506),
            .I(n2821));
    CascadeMux I__2762 (
            .O(N__24501),
            .I(n2721_cascade_));
    InMux I__2761 (
            .O(N__24498),
            .I(N__24495));
    LocalMux I__2760 (
            .O(N__24495),
            .I(N__24490));
    InMux I__2759 (
            .O(N__24494),
            .I(N__24487));
    InMux I__2758 (
            .O(N__24493),
            .I(N__24484));
    Odrv4 I__2757 (
            .O(N__24490),
            .I(n2717));
    LocalMux I__2756 (
            .O(N__24487),
            .I(n2717));
    LocalMux I__2755 (
            .O(N__24484),
            .I(n2717));
    InMux I__2754 (
            .O(N__24477),
            .I(N__24473));
    CascadeMux I__2753 (
            .O(N__24476),
            .I(N__24470));
    LocalMux I__2752 (
            .O(N__24473),
            .I(N__24466));
    InMux I__2751 (
            .O(N__24470),
            .I(N__24463));
    InMux I__2750 (
            .O(N__24469),
            .I(N__24460));
    Span4Mux_s2_h I__2749 (
            .O(N__24466),
            .I(N__24453));
    LocalMux I__2748 (
            .O(N__24463),
            .I(N__24453));
    LocalMux I__2747 (
            .O(N__24460),
            .I(N__24453));
    Odrv4 I__2746 (
            .O(N__24453),
            .I(n2718));
    CascadeMux I__2745 (
            .O(N__24450),
            .I(n14140_cascade_));
    InMux I__2744 (
            .O(N__24447),
            .I(N__24444));
    LocalMux I__2743 (
            .O(N__24444),
            .I(N__24441));
    Span4Mux_h I__2742 (
            .O(N__24441),
            .I(N__24438));
    Odrv4 I__2741 (
            .O(N__24438),
            .I(n14138));
    InMux I__2740 (
            .O(N__24435),
            .I(N__24431));
    CascadeMux I__2739 (
            .O(N__24434),
            .I(N__24428));
    LocalMux I__2738 (
            .O(N__24431),
            .I(N__24424));
    InMux I__2737 (
            .O(N__24428),
            .I(N__24421));
    InMux I__2736 (
            .O(N__24427),
            .I(N__24418));
    Span4Mux_v I__2735 (
            .O(N__24424),
            .I(N__24415));
    LocalMux I__2734 (
            .O(N__24421),
            .I(N__24410));
    LocalMux I__2733 (
            .O(N__24418),
            .I(N__24410));
    Odrv4 I__2732 (
            .O(N__24415),
            .I(n2716));
    Odrv4 I__2731 (
            .O(N__24410),
            .I(n2716));
    InMux I__2730 (
            .O(N__24405),
            .I(N__24402));
    LocalMux I__2729 (
            .O(N__24402),
            .I(N__24397));
    InMux I__2728 (
            .O(N__24401),
            .I(N__24394));
    InMux I__2727 (
            .O(N__24400),
            .I(N__24391));
    Odrv4 I__2726 (
            .O(N__24397),
            .I(n2715));
    LocalMux I__2725 (
            .O(N__24394),
            .I(n2715));
    LocalMux I__2724 (
            .O(N__24391),
            .I(n2715));
    CascadeMux I__2723 (
            .O(N__24384),
            .I(n14146_cascade_));
    InMux I__2722 (
            .O(N__24381),
            .I(N__24378));
    LocalMux I__2721 (
            .O(N__24378),
            .I(n14152));
    CascadeMux I__2720 (
            .O(N__24375),
            .I(N__24371));
    CascadeMux I__2719 (
            .O(N__24374),
            .I(N__24368));
    InMux I__2718 (
            .O(N__24371),
            .I(N__24364));
    InMux I__2717 (
            .O(N__24368),
            .I(N__24361));
    InMux I__2716 (
            .O(N__24367),
            .I(N__24358));
    LocalMux I__2715 (
            .O(N__24364),
            .I(n2722));
    LocalMux I__2714 (
            .O(N__24361),
            .I(n2722));
    LocalMux I__2713 (
            .O(N__24358),
            .I(n2722));
    InMux I__2712 (
            .O(N__24351),
            .I(N__24348));
    LocalMux I__2711 (
            .O(N__24348),
            .I(N__24345));
    Odrv4 I__2710 (
            .O(N__24345),
            .I(n2787));
    InMux I__2709 (
            .O(N__24342),
            .I(N__24339));
    LocalMux I__2708 (
            .O(N__24339),
            .I(N__24336));
    Odrv4 I__2707 (
            .O(N__24336),
            .I(n2795));
    InMux I__2706 (
            .O(N__24333),
            .I(N__24330));
    LocalMux I__2705 (
            .O(N__24330),
            .I(N__24325));
    InMux I__2704 (
            .O(N__24329),
            .I(N__24322));
    InMux I__2703 (
            .O(N__24328),
            .I(N__24319));
    Odrv4 I__2702 (
            .O(N__24325),
            .I(n2728));
    LocalMux I__2701 (
            .O(N__24322),
            .I(n2728));
    LocalMux I__2700 (
            .O(N__24319),
            .I(n2728));
    CascadeMux I__2699 (
            .O(N__24312),
            .I(N__24307));
    InMux I__2698 (
            .O(N__24311),
            .I(N__24304));
    InMux I__2697 (
            .O(N__24310),
            .I(N__24301));
    InMux I__2696 (
            .O(N__24307),
            .I(N__24298));
    LocalMux I__2695 (
            .O(N__24304),
            .I(n2712));
    LocalMux I__2694 (
            .O(N__24301),
            .I(n2712));
    LocalMux I__2693 (
            .O(N__24298),
            .I(n2712));
    InMux I__2692 (
            .O(N__24291),
            .I(N__24288));
    LocalMux I__2691 (
            .O(N__24288),
            .I(N__24284));
    InMux I__2690 (
            .O(N__24287),
            .I(N__24281));
    Span4Mux_v I__2689 (
            .O(N__24284),
            .I(N__24277));
    LocalMux I__2688 (
            .O(N__24281),
            .I(N__24274));
    InMux I__2687 (
            .O(N__24280),
            .I(N__24271));
    Odrv4 I__2686 (
            .O(N__24277),
            .I(n2514));
    Odrv4 I__2685 (
            .O(N__24274),
            .I(n2514));
    LocalMux I__2684 (
            .O(N__24271),
            .I(n2514));
    CascadeMux I__2683 (
            .O(N__24264),
            .I(N__24261));
    InMux I__2682 (
            .O(N__24261),
            .I(N__24258));
    LocalMux I__2681 (
            .O(N__24258),
            .I(N__24255));
    Span4Mux_h I__2680 (
            .O(N__24255),
            .I(N__24252));
    Odrv4 I__2679 (
            .O(N__24252),
            .I(n2581));
    CascadeMux I__2678 (
            .O(N__24249),
            .I(n2613_cascade_));
    InMux I__2677 (
            .O(N__24246),
            .I(N__24243));
    LocalMux I__2676 (
            .O(N__24243),
            .I(n14664));
    CascadeMux I__2675 (
            .O(N__24240),
            .I(n14670_cascade_));
    CascadeMux I__2674 (
            .O(N__24237),
            .I(n2643_cascade_));
    InMux I__2673 (
            .O(N__24234),
            .I(N__24229));
    InMux I__2672 (
            .O(N__24233),
            .I(N__24226));
    InMux I__2671 (
            .O(N__24232),
            .I(N__24223));
    LocalMux I__2670 (
            .O(N__24229),
            .I(N__24218));
    LocalMux I__2669 (
            .O(N__24226),
            .I(N__24218));
    LocalMux I__2668 (
            .O(N__24223),
            .I(n2713));
    Odrv4 I__2667 (
            .O(N__24218),
            .I(n2713));
    InMux I__2666 (
            .O(N__24213),
            .I(N__24210));
    LocalMux I__2665 (
            .O(N__24210),
            .I(N__24206));
    CascadeMux I__2664 (
            .O(N__24209),
            .I(N__24203));
    Span4Mux_v I__2663 (
            .O(N__24206),
            .I(N__24200));
    InMux I__2662 (
            .O(N__24203),
            .I(N__24197));
    Odrv4 I__2661 (
            .O(N__24200),
            .I(n2592));
    LocalMux I__2660 (
            .O(N__24197),
            .I(n2592));
    CascadeMux I__2659 (
            .O(N__24192),
            .I(n14889_cascade_));
    InMux I__2658 (
            .O(N__24189),
            .I(N__24185));
    CascadeMux I__2657 (
            .O(N__24188),
            .I(N__24182));
    LocalMux I__2656 (
            .O(N__24185),
            .I(N__24179));
    InMux I__2655 (
            .O(N__24182),
            .I(N__24175));
    Span4Mux_v I__2654 (
            .O(N__24179),
            .I(N__24171));
    InMux I__2653 (
            .O(N__24178),
            .I(N__24168));
    LocalMux I__2652 (
            .O(N__24175),
            .I(N__24165));
    InMux I__2651 (
            .O(N__24174),
            .I(N__24162));
    Odrv4 I__2650 (
            .O(N__24171),
            .I(n2525));
    LocalMux I__2649 (
            .O(N__24168),
            .I(n2525));
    Odrv4 I__2648 (
            .O(N__24165),
            .I(n2525));
    LocalMux I__2647 (
            .O(N__24162),
            .I(n2525));
    InMux I__2646 (
            .O(N__24153),
            .I(N__24150));
    LocalMux I__2645 (
            .O(N__24150),
            .I(N__24147));
    Odrv4 I__2644 (
            .O(N__24147),
            .I(n2582));
    CascadeMux I__2643 (
            .O(N__24144),
            .I(N__24140));
    CascadeMux I__2642 (
            .O(N__24143),
            .I(N__24137));
    InMux I__2641 (
            .O(N__24140),
            .I(N__24134));
    InMux I__2640 (
            .O(N__24137),
            .I(N__24131));
    LocalMux I__2639 (
            .O(N__24134),
            .I(N__24127));
    LocalMux I__2638 (
            .O(N__24131),
            .I(N__24124));
    InMux I__2637 (
            .O(N__24130),
            .I(N__24121));
    Odrv4 I__2636 (
            .O(N__24127),
            .I(n2515));
    Odrv4 I__2635 (
            .O(N__24124),
            .I(n2515));
    LocalMux I__2634 (
            .O(N__24121),
            .I(n2515));
    InMux I__2633 (
            .O(N__24114),
            .I(N__24110));
    CascadeMux I__2632 (
            .O(N__24113),
            .I(N__24107));
    LocalMux I__2631 (
            .O(N__24110),
            .I(N__24103));
    InMux I__2630 (
            .O(N__24107),
            .I(N__24100));
    CascadeMux I__2629 (
            .O(N__24106),
            .I(N__24097));
    Span4Mux_v I__2628 (
            .O(N__24103),
            .I(N__24094));
    LocalMux I__2627 (
            .O(N__24100),
            .I(N__24091));
    InMux I__2626 (
            .O(N__24097),
            .I(N__24088));
    Odrv4 I__2625 (
            .O(N__24094),
            .I(n2531));
    Odrv4 I__2624 (
            .O(N__24091),
            .I(n2531));
    LocalMux I__2623 (
            .O(N__24088),
            .I(n2531));
    InMux I__2622 (
            .O(N__24081),
            .I(N__24078));
    LocalMux I__2621 (
            .O(N__24078),
            .I(N__24075));
    Span4Mux_v I__2620 (
            .O(N__24075),
            .I(N__24072));
    Odrv4 I__2619 (
            .O(N__24072),
            .I(n2598));
    CascadeMux I__2618 (
            .O(N__24069),
            .I(N__24066));
    InMux I__2617 (
            .O(N__24066),
            .I(N__24063));
    LocalMux I__2616 (
            .O(N__24063),
            .I(N__24058));
    CascadeMux I__2615 (
            .O(N__24062),
            .I(N__24055));
    InMux I__2614 (
            .O(N__24061),
            .I(N__24052));
    Span4Mux_v I__2613 (
            .O(N__24058),
            .I(N__24049));
    InMux I__2612 (
            .O(N__24055),
            .I(N__24046));
    LocalMux I__2611 (
            .O(N__24052),
            .I(N__24043));
    Odrv4 I__2610 (
            .O(N__24049),
            .I(n2727));
    LocalMux I__2609 (
            .O(N__24046),
            .I(n2727));
    Odrv4 I__2608 (
            .O(N__24043),
            .I(n2727));
    InMux I__2607 (
            .O(N__24036),
            .I(N__24033));
    LocalMux I__2606 (
            .O(N__24033),
            .I(N__24030));
    Span4Mux_h I__2605 (
            .O(N__24030),
            .I(N__24027));
    Odrv4 I__2604 (
            .O(N__24027),
            .I(n2585));
    InMux I__2603 (
            .O(N__24024),
            .I(N__24020));
    InMux I__2602 (
            .O(N__24023),
            .I(N__24017));
    LocalMux I__2601 (
            .O(N__24020),
            .I(N__24013));
    LocalMux I__2600 (
            .O(N__24017),
            .I(N__24010));
    InMux I__2599 (
            .O(N__24016),
            .I(N__24007));
    Span4Mux_h I__2598 (
            .O(N__24013),
            .I(N__24004));
    Odrv4 I__2597 (
            .O(N__24010),
            .I(n2518));
    LocalMux I__2596 (
            .O(N__24007),
            .I(n2518));
    Odrv4 I__2595 (
            .O(N__24004),
            .I(n2518));
    InMux I__2594 (
            .O(N__23997),
            .I(N__23994));
    LocalMux I__2593 (
            .O(N__23994),
            .I(n14658));
    CascadeMux I__2592 (
            .O(N__23991),
            .I(n2617_cascade_));
    CascadeMux I__2591 (
            .O(N__23988),
            .I(N__23985));
    InMux I__2590 (
            .O(N__23985),
            .I(N__23982));
    LocalMux I__2589 (
            .O(N__23982),
            .I(n14324));
    CascadeMux I__2588 (
            .O(N__23979),
            .I(N__23976));
    InMux I__2587 (
            .O(N__23976),
            .I(N__23972));
    InMux I__2586 (
            .O(N__23975),
            .I(N__23969));
    LocalMux I__2585 (
            .O(N__23972),
            .I(n2516));
    LocalMux I__2584 (
            .O(N__23969),
            .I(n2516));
    InMux I__2583 (
            .O(N__23964),
            .I(N__23959));
    InMux I__2582 (
            .O(N__23963),
            .I(N__23956));
    InMux I__2581 (
            .O(N__23962),
            .I(N__23953));
    LocalMux I__2580 (
            .O(N__23959),
            .I(N__23950));
    LocalMux I__2579 (
            .O(N__23956),
            .I(N__23945));
    LocalMux I__2578 (
            .O(N__23953),
            .I(N__23945));
    Span4Mux_v I__2577 (
            .O(N__23950),
            .I(N__23942));
    Odrv4 I__2576 (
            .O(N__23945),
            .I(n2512));
    Odrv4 I__2575 (
            .O(N__23942),
            .I(n2512));
    InMux I__2574 (
            .O(N__23937),
            .I(N__23933));
    InMux I__2573 (
            .O(N__23936),
            .I(N__23930));
    LocalMux I__2572 (
            .O(N__23933),
            .I(N__23924));
    LocalMux I__2571 (
            .O(N__23930),
            .I(N__23924));
    InMux I__2570 (
            .O(N__23929),
            .I(N__23921));
    Odrv4 I__2569 (
            .O(N__23924),
            .I(n2513));
    LocalMux I__2568 (
            .O(N__23921),
            .I(n2513));
    CascadeMux I__2567 (
            .O(N__23916),
            .I(n14330_cascade_));
    InMux I__2566 (
            .O(N__23913),
            .I(N__23909));
    InMux I__2565 (
            .O(N__23912),
            .I(N__23906));
    LocalMux I__2564 (
            .O(N__23909),
            .I(N__23903));
    LocalMux I__2563 (
            .O(N__23906),
            .I(N__23900));
    Span4Mux_h I__2562 (
            .O(N__23903),
            .I(N__23897));
    Odrv4 I__2561 (
            .O(N__23900),
            .I(n2511));
    Odrv4 I__2560 (
            .O(N__23897),
            .I(n2511));
    CascadeMux I__2559 (
            .O(N__23892),
            .I(N__23889));
    InMux I__2558 (
            .O(N__23889),
            .I(N__23884));
    InMux I__2557 (
            .O(N__23888),
            .I(N__23879));
    InMux I__2556 (
            .O(N__23887),
            .I(N__23879));
    LocalMux I__2555 (
            .O(N__23884),
            .I(n2523));
    LocalMux I__2554 (
            .O(N__23879),
            .I(n2523));
    CascadeMux I__2553 (
            .O(N__23874),
            .I(n2544_cascade_));
    InMux I__2552 (
            .O(N__23871),
            .I(N__23868));
    LocalMux I__2551 (
            .O(N__23868),
            .I(N__23865));
    Odrv4 I__2550 (
            .O(N__23865),
            .I(n2590));
    CascadeMux I__2549 (
            .O(N__23862),
            .I(N__23859));
    InMux I__2548 (
            .O(N__23859),
            .I(N__23856));
    LocalMux I__2547 (
            .O(N__23856),
            .I(N__23853));
    Odrv12 I__2546 (
            .O(N__23853),
            .I(n2591));
    CascadeMux I__2545 (
            .O(N__23850),
            .I(N__23846));
    InMux I__2544 (
            .O(N__23849),
            .I(N__23843));
    InMux I__2543 (
            .O(N__23846),
            .I(N__23840));
    LocalMux I__2542 (
            .O(N__23843),
            .I(N__23837));
    LocalMux I__2541 (
            .O(N__23840),
            .I(N__23834));
    Span4Mux_v I__2540 (
            .O(N__23837),
            .I(N__23830));
    Span4Mux_v I__2539 (
            .O(N__23834),
            .I(N__23827));
    InMux I__2538 (
            .O(N__23833),
            .I(N__23824));
    Odrv4 I__2537 (
            .O(N__23830),
            .I(n2530));
    Odrv4 I__2536 (
            .O(N__23827),
            .I(n2530));
    LocalMux I__2535 (
            .O(N__23824),
            .I(n2530));
    CascadeMux I__2534 (
            .O(N__23817),
            .I(N__23814));
    InMux I__2533 (
            .O(N__23814),
            .I(N__23811));
    LocalMux I__2532 (
            .O(N__23811),
            .I(N__23808));
    Span4Mux_h I__2531 (
            .O(N__23808),
            .I(N__23805));
    Span4Mux_s0_h I__2530 (
            .O(N__23805),
            .I(N__23802));
    Odrv4 I__2529 (
            .O(N__23802),
            .I(n2597));
    CascadeMux I__2528 (
            .O(N__23799),
            .I(n2629_cascade_));
    InMux I__2527 (
            .O(N__23796),
            .I(N__23793));
    LocalMux I__2526 (
            .O(N__23793),
            .I(n14656));
    InMux I__2525 (
            .O(N__23790),
            .I(N__23787));
    LocalMux I__2524 (
            .O(N__23787),
            .I(N__23784));
    Span4Mux_v I__2523 (
            .O(N__23784),
            .I(N__23781));
    Sp12to4 I__2522 (
            .O(N__23781),
            .I(N__23778));
    Odrv12 I__2521 (
            .O(N__23778),
            .I(n2601));
    InMux I__2520 (
            .O(N__23775),
            .I(N__23772));
    LocalMux I__2519 (
            .O(N__23772),
            .I(N__23769));
    Odrv4 I__2518 (
            .O(N__23769),
            .I(n2584));
    CascadeMux I__2517 (
            .O(N__23766),
            .I(N__23762));
    InMux I__2516 (
            .O(N__23765),
            .I(N__23759));
    InMux I__2515 (
            .O(N__23762),
            .I(N__23756));
    LocalMux I__2514 (
            .O(N__23759),
            .I(N__23752));
    LocalMux I__2513 (
            .O(N__23756),
            .I(N__23749));
    InMux I__2512 (
            .O(N__23755),
            .I(N__23746));
    Odrv4 I__2511 (
            .O(N__23752),
            .I(n2517));
    Odrv4 I__2510 (
            .O(N__23749),
            .I(n2517));
    LocalMux I__2509 (
            .O(N__23746),
            .I(n2517));
    CascadeMux I__2508 (
            .O(N__23739),
            .I(n2328_cascade_));
    CascadeMux I__2507 (
            .O(N__23736),
            .I(n14442_cascade_));
    CascadeMux I__2506 (
            .O(N__23733),
            .I(n14448_cascade_));
    InMux I__2505 (
            .O(N__23730),
            .I(N__23727));
    LocalMux I__2504 (
            .O(N__23727),
            .I(n14450));
    CascadeMux I__2503 (
            .O(N__23724),
            .I(N__23721));
    InMux I__2502 (
            .O(N__23721),
            .I(N__23718));
    LocalMux I__2501 (
            .O(N__23718),
            .I(N__23715));
    Odrv12 I__2500 (
            .O(N__23715),
            .I(n2593));
    InMux I__2499 (
            .O(N__23712),
            .I(N__23708));
    CascadeMux I__2498 (
            .O(N__23711),
            .I(N__23705));
    LocalMux I__2497 (
            .O(N__23708),
            .I(N__23701));
    InMux I__2496 (
            .O(N__23705),
            .I(N__23698));
    InMux I__2495 (
            .O(N__23704),
            .I(N__23695));
    Odrv4 I__2494 (
            .O(N__23701),
            .I(n2422));
    LocalMux I__2493 (
            .O(N__23698),
            .I(n2422));
    LocalMux I__2492 (
            .O(N__23695),
            .I(n2422));
    InMux I__2491 (
            .O(N__23688),
            .I(N__23685));
    LocalMux I__2490 (
            .O(N__23685),
            .I(N__23682));
    Span4Mux_h I__2489 (
            .O(N__23682),
            .I(N__23679));
    Odrv4 I__2488 (
            .O(N__23679),
            .I(n2489));
    CascadeMux I__2487 (
            .O(N__23676),
            .I(N__23673));
    InMux I__2486 (
            .O(N__23673),
            .I(N__23669));
    InMux I__2485 (
            .O(N__23672),
            .I(N__23666));
    LocalMux I__2484 (
            .O(N__23669),
            .I(N__23663));
    LocalMux I__2483 (
            .O(N__23666),
            .I(n2521));
    Odrv12 I__2482 (
            .O(N__23663),
            .I(n2521));
    CascadeMux I__2481 (
            .O(N__23658),
            .I(N__23655));
    InMux I__2480 (
            .O(N__23655),
            .I(N__23650));
    InMux I__2479 (
            .O(N__23654),
            .I(N__23645));
    InMux I__2478 (
            .O(N__23653),
            .I(N__23645));
    LocalMux I__2477 (
            .O(N__23650),
            .I(n2526));
    LocalMux I__2476 (
            .O(N__23645),
            .I(n2526));
    CascadeMux I__2475 (
            .O(N__23640),
            .I(n2521_cascade_));
    InMux I__2474 (
            .O(N__23637),
            .I(N__23634));
    LocalMux I__2473 (
            .O(N__23634),
            .I(n14312));
    CascadeMux I__2472 (
            .O(N__23631),
            .I(N__23628));
    InMux I__2471 (
            .O(N__23628),
            .I(N__23624));
    InMux I__2470 (
            .O(N__23627),
            .I(N__23620));
    LocalMux I__2469 (
            .O(N__23624),
            .I(N__23617));
    InMux I__2468 (
            .O(N__23623),
            .I(N__23614));
    LocalMux I__2467 (
            .O(N__23620),
            .I(n2423));
    Odrv4 I__2466 (
            .O(N__23617),
            .I(n2423));
    LocalMux I__2465 (
            .O(N__23614),
            .I(n2423));
    CascadeMux I__2464 (
            .O(N__23607),
            .I(n2425_cascade_));
    InMux I__2463 (
            .O(N__23604),
            .I(N__23601));
    LocalMux I__2462 (
            .O(N__23601),
            .I(n14632));
    CascadeMux I__2461 (
            .O(N__23598),
            .I(N__23594));
    InMux I__2460 (
            .O(N__23597),
            .I(N__23591));
    InMux I__2459 (
            .O(N__23594),
            .I(N__23588));
    LocalMux I__2458 (
            .O(N__23591),
            .I(N__23585));
    LocalMux I__2457 (
            .O(N__23588),
            .I(N__23582));
    Span4Mux_v I__2456 (
            .O(N__23585),
            .I(N__23578));
    Span4Mux_s3_h I__2455 (
            .O(N__23582),
            .I(N__23575));
    InMux I__2454 (
            .O(N__23581),
            .I(N__23572));
    Odrv4 I__2453 (
            .O(N__23578),
            .I(n2419));
    Odrv4 I__2452 (
            .O(N__23575),
            .I(n2419));
    LocalMux I__2451 (
            .O(N__23572),
            .I(n2419));
    InMux I__2450 (
            .O(N__23565),
            .I(N__23561));
    InMux I__2449 (
            .O(N__23564),
            .I(N__23557));
    LocalMux I__2448 (
            .O(N__23561),
            .I(N__23554));
    InMux I__2447 (
            .O(N__23560),
            .I(N__23551));
    LocalMux I__2446 (
            .O(N__23557),
            .I(n2415));
    Odrv12 I__2445 (
            .O(N__23554),
            .I(n2415));
    LocalMux I__2444 (
            .O(N__23551),
            .I(n2415));
    CascadeMux I__2443 (
            .O(N__23544),
            .I(n14456_cascade_));
    CascadeMux I__2442 (
            .O(N__23541),
            .I(n2346_cascade_));
    CascadeMux I__2441 (
            .O(N__23538),
            .I(N__23534));
    CascadeMux I__2440 (
            .O(N__23537),
            .I(N__23531));
    InMux I__2439 (
            .O(N__23534),
            .I(N__23528));
    InMux I__2438 (
            .O(N__23531),
            .I(N__23525));
    LocalMux I__2437 (
            .O(N__23528),
            .I(N__23521));
    LocalMux I__2436 (
            .O(N__23525),
            .I(N__23518));
    InMux I__2435 (
            .O(N__23524),
            .I(N__23515));
    Odrv4 I__2434 (
            .O(N__23521),
            .I(n2417));
    Odrv4 I__2433 (
            .O(N__23518),
            .I(n2417));
    LocalMux I__2432 (
            .O(N__23515),
            .I(n2417));
    InMux I__2431 (
            .O(N__23508),
            .I(N__23503));
    InMux I__2430 (
            .O(N__23507),
            .I(N__23500));
    InMux I__2429 (
            .O(N__23506),
            .I(N__23497));
    LocalMux I__2428 (
            .O(N__23503),
            .I(N__23494));
    LocalMux I__2427 (
            .O(N__23500),
            .I(N__23491));
    LocalMux I__2426 (
            .O(N__23497),
            .I(n2414));
    Odrv4 I__2425 (
            .O(N__23494),
            .I(n2414));
    Odrv4 I__2424 (
            .O(N__23491),
            .I(n2414));
    CascadeMux I__2423 (
            .O(N__23484),
            .I(N__23481));
    InMux I__2422 (
            .O(N__23481),
            .I(N__23478));
    LocalMux I__2421 (
            .O(N__23478),
            .I(N__23475));
    Odrv4 I__2420 (
            .O(N__23475),
            .I(n13790));
    InMux I__2419 (
            .O(N__23472),
            .I(N__23469));
    LocalMux I__2418 (
            .O(N__23469),
            .I(n14318));
    CascadeMux I__2417 (
            .O(N__23466),
            .I(N__23463));
    InMux I__2416 (
            .O(N__23463),
            .I(N__23460));
    LocalMux I__2415 (
            .O(N__23460),
            .I(N__23456));
    CascadeMux I__2414 (
            .O(N__23459),
            .I(N__23453));
    Span4Mux_v I__2413 (
            .O(N__23456),
            .I(N__23450));
    InMux I__2412 (
            .O(N__23453),
            .I(N__23447));
    Span4Mux_s1_h I__2411 (
            .O(N__23450),
            .I(N__23441));
    LocalMux I__2410 (
            .O(N__23447),
            .I(N__23441));
    InMux I__2409 (
            .O(N__23446),
            .I(N__23438));
    Odrv4 I__2408 (
            .O(N__23441),
            .I(n2529));
    LocalMux I__2407 (
            .O(N__23438),
            .I(n2529));
    InMux I__2406 (
            .O(N__23433),
            .I(N__23430));
    LocalMux I__2405 (
            .O(N__23430),
            .I(n11942));
    CascadeMux I__2404 (
            .O(N__23427),
            .I(N__23424));
    InMux I__2403 (
            .O(N__23424),
            .I(N__23421));
    LocalMux I__2402 (
            .O(N__23421),
            .I(n13816));
    CascadeMux I__2401 (
            .O(N__23418),
            .I(n14622_cascade_));
    InMux I__2400 (
            .O(N__23415),
            .I(N__23412));
    LocalMux I__2399 (
            .O(N__23412),
            .I(n14638));
    CascadeMux I__2398 (
            .O(N__23409),
            .I(N__23406));
    InMux I__2397 (
            .O(N__23406),
            .I(N__23402));
    InMux I__2396 (
            .O(N__23405),
            .I(N__23399));
    LocalMux I__2395 (
            .O(N__23402),
            .I(N__23396));
    LocalMux I__2394 (
            .O(N__23399),
            .I(n2420));
    Odrv4 I__2393 (
            .O(N__23396),
            .I(n2420));
    CascadeMux I__2392 (
            .O(N__23391),
            .I(n2420_cascade_));
    InMux I__2391 (
            .O(N__23388),
            .I(N__23385));
    LocalMux I__2390 (
            .O(N__23385),
            .I(n14612));
    InMux I__2389 (
            .O(N__23382),
            .I(N__23379));
    LocalMux I__2388 (
            .O(N__23379),
            .I(n14616));
    CascadeMux I__2387 (
            .O(N__23376),
            .I(N__23373));
    InMux I__2386 (
            .O(N__23373),
            .I(N__23369));
    InMux I__2385 (
            .O(N__23372),
            .I(N__23365));
    LocalMux I__2384 (
            .O(N__23369),
            .I(N__23362));
    InMux I__2383 (
            .O(N__23368),
            .I(N__23359));
    LocalMux I__2382 (
            .O(N__23365),
            .I(n2426));
    Odrv4 I__2381 (
            .O(N__23362),
            .I(n2426));
    LocalMux I__2380 (
            .O(N__23359),
            .I(n2426));
    CascadeMux I__2379 (
            .O(N__23352),
            .I(N__23348));
    InMux I__2378 (
            .O(N__23351),
            .I(N__23345));
    InMux I__2377 (
            .O(N__23348),
            .I(N__23342));
    LocalMux I__2376 (
            .O(N__23345),
            .I(N__23338));
    LocalMux I__2375 (
            .O(N__23342),
            .I(N__23335));
    InMux I__2374 (
            .O(N__23341),
            .I(N__23332));
    Odrv4 I__2373 (
            .O(N__23338),
            .I(n2421));
    Odrv4 I__2372 (
            .O(N__23335),
            .I(n2421));
    LocalMux I__2371 (
            .O(N__23332),
            .I(n2421));
    InMux I__2370 (
            .O(N__23325),
            .I(N__23321));
    InMux I__2369 (
            .O(N__23324),
            .I(N__23318));
    LocalMux I__2368 (
            .O(N__23321),
            .I(N__23315));
    LocalMux I__2367 (
            .O(N__23318),
            .I(N__23311));
    Span4Mux_s2_h I__2366 (
            .O(N__23315),
            .I(N__23308));
    InMux I__2365 (
            .O(N__23314),
            .I(N__23305));
    Odrv4 I__2364 (
            .O(N__23311),
            .I(n2413));
    Odrv4 I__2363 (
            .O(N__23308),
            .I(n2413));
    LocalMux I__2362 (
            .O(N__23305),
            .I(n2413));
    InMux I__2361 (
            .O(N__23298),
            .I(N__23294));
    InMux I__2360 (
            .O(N__23297),
            .I(N__23291));
    LocalMux I__2359 (
            .O(N__23294),
            .I(\debounce.cnt_reg_9 ));
    LocalMux I__2358 (
            .O(N__23291),
            .I(\debounce.cnt_reg_9 ));
    InMux I__2357 (
            .O(N__23286),
            .I(N__23282));
    InMux I__2356 (
            .O(N__23285),
            .I(N__23279));
    LocalMux I__2355 (
            .O(N__23282),
            .I(\debounce.cnt_reg_8 ));
    LocalMux I__2354 (
            .O(N__23279),
            .I(\debounce.cnt_reg_8 ));
    CascadeMux I__2353 (
            .O(N__23274),
            .I(N__23271));
    InMux I__2352 (
            .O(N__23271),
            .I(N__23268));
    LocalMux I__2351 (
            .O(N__23268),
            .I(N__23264));
    InMux I__2350 (
            .O(N__23267),
            .I(N__23261));
    Span4Mux_s1_v I__2349 (
            .O(N__23264),
            .I(N__23258));
    LocalMux I__2348 (
            .O(N__23261),
            .I(\debounce.cnt_reg_4 ));
    Odrv4 I__2347 (
            .O(N__23258),
            .I(\debounce.cnt_reg_4 ));
    InMux I__2346 (
            .O(N__23253),
            .I(N__23249));
    InMux I__2345 (
            .O(N__23252),
            .I(N__23246));
    LocalMux I__2344 (
            .O(N__23249),
            .I(\debounce.cnt_reg_5 ));
    LocalMux I__2343 (
            .O(N__23246),
            .I(\debounce.cnt_reg_5 ));
    CascadeMux I__2342 (
            .O(N__23241),
            .I(N__23238));
    InMux I__2341 (
            .O(N__23238),
            .I(N__23235));
    LocalMux I__2340 (
            .O(N__23235),
            .I(n2976));
    CascadeMux I__2339 (
            .O(N__23232),
            .I(N__23228));
    InMux I__2338 (
            .O(N__23231),
            .I(N__23225));
    InMux I__2337 (
            .O(N__23228),
            .I(N__23222));
    LocalMux I__2336 (
            .O(N__23225),
            .I(N__23217));
    LocalMux I__2335 (
            .O(N__23222),
            .I(N__23217));
    Odrv4 I__2334 (
            .O(N__23217),
            .I(n2432));
    CascadeMux I__2333 (
            .O(N__23214),
            .I(n2432_cascade_));
    CascadeMux I__2332 (
            .O(N__23211),
            .I(N__23208));
    InMux I__2331 (
            .O(N__23208),
            .I(N__23204));
    InMux I__2330 (
            .O(N__23207),
            .I(N__23201));
    LocalMux I__2329 (
            .O(N__23204),
            .I(n2433));
    LocalMux I__2328 (
            .O(N__23201),
            .I(n2433));
    CascadeMux I__2327 (
            .O(N__23196),
            .I(N__23193));
    InMux I__2326 (
            .O(N__23193),
            .I(N__23188));
    InMux I__2325 (
            .O(N__23192),
            .I(N__23185));
    InMux I__2324 (
            .O(N__23191),
            .I(N__23182));
    LocalMux I__2323 (
            .O(N__23188),
            .I(n2431));
    LocalMux I__2322 (
            .O(N__23185),
            .I(n2431));
    LocalMux I__2321 (
            .O(N__23182),
            .I(n2431));
    CascadeMux I__2320 (
            .O(N__23175),
            .I(N__23171));
    CascadeMux I__2319 (
            .O(N__23174),
            .I(N__23167));
    InMux I__2318 (
            .O(N__23171),
            .I(N__23164));
    InMux I__2317 (
            .O(N__23170),
            .I(N__23161));
    InMux I__2316 (
            .O(N__23167),
            .I(N__23158));
    LocalMux I__2315 (
            .O(N__23164),
            .I(n2430));
    LocalMux I__2314 (
            .O(N__23161),
            .I(n2430));
    LocalMux I__2313 (
            .O(N__23158),
            .I(n2430));
    CascadeMux I__2312 (
            .O(N__23151),
            .I(n11946_cascade_));
    CascadeMux I__2311 (
            .O(N__23148),
            .I(N__23145));
    InMux I__2310 (
            .O(N__23145),
            .I(N__23140));
    InMux I__2309 (
            .O(N__23144),
            .I(N__23137));
    InMux I__2308 (
            .O(N__23143),
            .I(N__23134));
    LocalMux I__2307 (
            .O(N__23140),
            .I(N__23131));
    LocalMux I__2306 (
            .O(N__23137),
            .I(n2429));
    LocalMux I__2305 (
            .O(N__23134),
            .I(n2429));
    Odrv4 I__2304 (
            .O(N__23131),
            .I(n2429));
    CascadeMux I__2303 (
            .O(N__23124),
            .I(N__23120));
    InMux I__2302 (
            .O(N__23123),
            .I(N__23117));
    InMux I__2301 (
            .O(N__23120),
            .I(N__23114));
    LocalMux I__2300 (
            .O(N__23117),
            .I(N__23111));
    LocalMux I__2299 (
            .O(N__23114),
            .I(N__23108));
    Odrv4 I__2298 (
            .O(N__23111),
            .I(n2427));
    Odrv4 I__2297 (
            .O(N__23108),
            .I(n2427));
    InMux I__2296 (
            .O(N__23103),
            .I(N__23099));
    CascadeMux I__2295 (
            .O(N__23102),
            .I(N__23096));
    LocalMux I__2294 (
            .O(N__23099),
            .I(N__23092));
    InMux I__2293 (
            .O(N__23096),
            .I(N__23089));
    InMux I__2292 (
            .O(N__23095),
            .I(N__23086));
    Odrv4 I__2291 (
            .O(N__23092),
            .I(n2424));
    LocalMux I__2290 (
            .O(N__23089),
            .I(n2424));
    LocalMux I__2289 (
            .O(N__23086),
            .I(n2424));
    CascadeMux I__2288 (
            .O(N__23079),
            .I(n2427_cascade_));
    InMux I__2287 (
            .O(N__23076),
            .I(N__23072));
    InMux I__2286 (
            .O(N__23075),
            .I(N__23069));
    LocalMux I__2285 (
            .O(N__23072),
            .I(N__23066));
    LocalMux I__2284 (
            .O(N__23069),
            .I(N__23063));
    Odrv4 I__2283 (
            .O(N__23066),
            .I(n2428));
    Odrv4 I__2282 (
            .O(N__23063),
            .I(n2428));
    InMux I__2281 (
            .O(N__23058),
            .I(n12842));
    InMux I__2280 (
            .O(N__23055),
            .I(n12843));
    InMux I__2279 (
            .O(N__23052),
            .I(n12844));
    InMux I__2278 (
            .O(N__23049),
            .I(n12845));
    InMux I__2277 (
            .O(N__23046),
            .I(bfn_2_32_0_));
    InMux I__2276 (
            .O(N__23043),
            .I(n12847));
    InMux I__2275 (
            .O(N__23040),
            .I(n12848));
    InMux I__2274 (
            .O(N__23037),
            .I(n12849));
    InMux I__2273 (
            .O(N__23034),
            .I(N__23030));
    InMux I__2272 (
            .O(N__23033),
            .I(N__23027));
    LocalMux I__2271 (
            .O(N__23030),
            .I(\debounce.cnt_reg_0 ));
    LocalMux I__2270 (
            .O(N__23027),
            .I(\debounce.cnt_reg_0 ));
    InMux I__2269 (
            .O(N__23022),
            .I(N__23018));
    InMux I__2268 (
            .O(N__23021),
            .I(N__23015));
    LocalMux I__2267 (
            .O(N__23018),
            .I(\debounce.cnt_reg_7 ));
    LocalMux I__2266 (
            .O(N__23015),
            .I(\debounce.cnt_reg_7 ));
    CascadeMux I__2265 (
            .O(N__23010),
            .I(N__23006));
    InMux I__2264 (
            .O(N__23009),
            .I(N__23003));
    InMux I__2263 (
            .O(N__23006),
            .I(N__23000));
    LocalMux I__2262 (
            .O(N__23003),
            .I(\debounce.cnt_reg_1 ));
    LocalMux I__2261 (
            .O(N__23000),
            .I(\debounce.cnt_reg_1 ));
    InMux I__2260 (
            .O(N__22995),
            .I(N__22991));
    InMux I__2259 (
            .O(N__22994),
            .I(N__22988));
    LocalMux I__2258 (
            .O(N__22991),
            .I(\debounce.cnt_reg_2 ));
    LocalMux I__2257 (
            .O(N__22988),
            .I(\debounce.cnt_reg_2 ));
    InMux I__2256 (
            .O(N__22983),
            .I(n12833));
    InMux I__2255 (
            .O(N__22980),
            .I(n12834));
    InMux I__2254 (
            .O(N__22977),
            .I(n12835));
    InMux I__2253 (
            .O(N__22974),
            .I(n12836));
    InMux I__2252 (
            .O(N__22971),
            .I(n12837));
    InMux I__2251 (
            .O(N__22968),
            .I(bfn_2_31_0_));
    InMux I__2250 (
            .O(N__22965),
            .I(n12839));
    InMux I__2249 (
            .O(N__22962),
            .I(n12840));
    InMux I__2248 (
            .O(N__22959),
            .I(n12841));
    InMux I__2247 (
            .O(N__22956),
            .I(n12824));
    InMux I__2246 (
            .O(N__22953),
            .I(n12825));
    InMux I__2245 (
            .O(N__22950),
            .I(n12826));
    InMux I__2244 (
            .O(N__22947),
            .I(n12827));
    InMux I__2243 (
            .O(N__22944),
            .I(n12828));
    InMux I__2242 (
            .O(N__22941),
            .I(n12829));
    InMux I__2241 (
            .O(N__22938),
            .I(bfn_2_30_0_));
    InMux I__2240 (
            .O(N__22935),
            .I(n12831));
    InMux I__2239 (
            .O(N__22932),
            .I(n12832));
    InMux I__2238 (
            .O(N__22929),
            .I(N__22926));
    LocalMux I__2237 (
            .O(N__22926),
            .I(N__22923));
    Odrv4 I__2236 (
            .O(N__22923),
            .I(n2780));
    InMux I__2235 (
            .O(N__22920),
            .I(N__22916));
    InMux I__2234 (
            .O(N__22919),
            .I(N__22913));
    LocalMux I__2233 (
            .O(N__22916),
            .I(N__22909));
    LocalMux I__2232 (
            .O(N__22913),
            .I(N__22906));
    InMux I__2231 (
            .O(N__22912),
            .I(N__22903));
    Odrv4 I__2230 (
            .O(N__22909),
            .I(n2817));
    Odrv4 I__2229 (
            .O(N__22906),
            .I(n2817));
    LocalMux I__2228 (
            .O(N__22903),
            .I(n2817));
    CascadeMux I__2227 (
            .O(N__22896),
            .I(N__22893));
    InMux I__2226 (
            .O(N__22893),
            .I(N__22890));
    LocalMux I__2225 (
            .O(N__22890),
            .I(n2884));
    InMux I__2224 (
            .O(N__22887),
            .I(N__22884));
    LocalMux I__2223 (
            .O(N__22884),
            .I(n2877));
    InMux I__2222 (
            .O(N__22881),
            .I(N__22878));
    LocalMux I__2221 (
            .O(N__22878),
            .I(N__22875));
    Odrv4 I__2220 (
            .O(N__22875),
            .I(n2897));
    CascadeMux I__2219 (
            .O(N__22872),
            .I(N__22869));
    InMux I__2218 (
            .O(N__22869),
            .I(N__22866));
    LocalMux I__2217 (
            .O(N__22866),
            .I(N__22861));
    InMux I__2216 (
            .O(N__22865),
            .I(N__22858));
    InMux I__2215 (
            .O(N__22864),
            .I(N__22855));
    Odrv4 I__2214 (
            .O(N__22861),
            .I(n2830));
    LocalMux I__2213 (
            .O(N__22858),
            .I(n2830));
    LocalMux I__2212 (
            .O(N__22855),
            .I(n2830));
    InMux I__2211 (
            .O(N__22848),
            .I(N__22844));
    InMux I__2210 (
            .O(N__22847),
            .I(N__22841));
    LocalMux I__2209 (
            .O(N__22844),
            .I(n2811));
    LocalMux I__2208 (
            .O(N__22841),
            .I(n2811));
    InMux I__2207 (
            .O(N__22836),
            .I(N__22833));
    LocalMux I__2206 (
            .O(N__22833),
            .I(n2878));
    InMux I__2205 (
            .O(N__22830),
            .I(bfn_2_29_0_));
    CascadeMux I__2204 (
            .O(N__22827),
            .I(N__22824));
    InMux I__2203 (
            .O(N__22824),
            .I(N__22820));
    InMux I__2202 (
            .O(N__22823),
            .I(N__22817));
    LocalMux I__2201 (
            .O(N__22820),
            .I(n2933));
    LocalMux I__2200 (
            .O(N__22817),
            .I(n2933));
    InMux I__2199 (
            .O(N__22812),
            .I(N__22809));
    LocalMux I__2198 (
            .O(N__22809),
            .I(n3000));
    InMux I__2197 (
            .O(N__22806),
            .I(n12823));
    InMux I__2196 (
            .O(N__22803),
            .I(N__22800));
    LocalMux I__2195 (
            .O(N__22800),
            .I(N__22797));
    Odrv4 I__2194 (
            .O(N__22797),
            .I(n2789));
    InMux I__2193 (
            .O(N__22794),
            .I(N__22789));
    InMux I__2192 (
            .O(N__22793),
            .I(N__22784));
    InMux I__2191 (
            .O(N__22792),
            .I(N__22784));
    LocalMux I__2190 (
            .O(N__22789),
            .I(N__22779));
    LocalMux I__2189 (
            .O(N__22784),
            .I(N__22779));
    Odrv12 I__2188 (
            .O(N__22779),
            .I(n2711));
    InMux I__2187 (
            .O(N__22776),
            .I(N__22773));
    LocalMux I__2186 (
            .O(N__22773),
            .I(N__22770));
    Odrv4 I__2185 (
            .O(N__22770),
            .I(n2778));
    InMux I__2184 (
            .O(N__22767),
            .I(N__22764));
    LocalMux I__2183 (
            .O(N__22764),
            .I(N__22761));
    Odrv4 I__2182 (
            .O(N__22761),
            .I(n2781));
    InMux I__2181 (
            .O(N__22758),
            .I(N__22753));
    InMux I__2180 (
            .O(N__22757),
            .I(N__22750));
    InMux I__2179 (
            .O(N__22756),
            .I(N__22747));
    LocalMux I__2178 (
            .O(N__22753),
            .I(n2714));
    LocalMux I__2177 (
            .O(N__22750),
            .I(n2714));
    LocalMux I__2176 (
            .O(N__22747),
            .I(n2714));
    InMux I__2175 (
            .O(N__22740),
            .I(N__22737));
    LocalMux I__2174 (
            .O(N__22737),
            .I(N__22734));
    Odrv12 I__2173 (
            .O(N__22734),
            .I(n2800));
    CascadeMux I__2172 (
            .O(N__22731),
            .I(N__22728));
    InMux I__2171 (
            .O(N__22728),
            .I(N__22724));
    CascadeMux I__2170 (
            .O(N__22727),
            .I(N__22720));
    LocalMux I__2169 (
            .O(N__22724),
            .I(N__22717));
    InMux I__2168 (
            .O(N__22723),
            .I(N__22714));
    InMux I__2167 (
            .O(N__22720),
            .I(N__22711));
    Span4Mux_s3_v I__2166 (
            .O(N__22717),
            .I(N__22706));
    LocalMux I__2165 (
            .O(N__22714),
            .I(N__22706));
    LocalMux I__2164 (
            .O(N__22711),
            .I(n2832));
    Odrv4 I__2163 (
            .O(N__22706),
            .I(n2832));
    InMux I__2162 (
            .O(N__22701),
            .I(N__22698));
    LocalMux I__2161 (
            .O(N__22698),
            .I(N__22695));
    Odrv12 I__2160 (
            .O(N__22695),
            .I(n2794));
    CascadeMux I__2159 (
            .O(N__22692),
            .I(N__22689));
    InMux I__2158 (
            .O(N__22689),
            .I(N__22686));
    LocalMux I__2157 (
            .O(N__22686),
            .I(n2887));
    InMux I__2156 (
            .O(N__22683),
            .I(N__22680));
    LocalMux I__2155 (
            .O(N__22680),
            .I(N__22677));
    Odrv4 I__2154 (
            .O(N__22677),
            .I(n2779));
    CascadeMux I__2153 (
            .O(N__22674),
            .I(n2811_cascade_));
    InMux I__2152 (
            .O(N__22671),
            .I(N__22668));
    LocalMux I__2151 (
            .O(N__22668),
            .I(N__22665));
    Odrv4 I__2150 (
            .O(N__22665),
            .I(n14708));
    InMux I__2149 (
            .O(N__22662),
            .I(n12791));
    InMux I__2148 (
            .O(N__22659),
            .I(n12792));
    InMux I__2147 (
            .O(N__22656),
            .I(n12793));
    InMux I__2146 (
            .O(N__22653),
            .I(n12794));
    InMux I__2145 (
            .O(N__22650),
            .I(bfn_2_26_0_));
    InMux I__2144 (
            .O(N__22647),
            .I(n12796));
    CascadeMux I__2143 (
            .O(N__22644),
            .I(n14158_cascade_));
    InMux I__2142 (
            .O(N__22641),
            .I(N__22638));
    LocalMux I__2141 (
            .O(N__22638),
            .I(N__22635));
    Odrv4 I__2140 (
            .O(N__22635),
            .I(n2790));
    CascadeMux I__2139 (
            .O(N__22632),
            .I(n2742_cascade_));
    InMux I__2138 (
            .O(N__22629),
            .I(n12783));
    InMux I__2137 (
            .O(N__22626),
            .I(n12784));
    InMux I__2136 (
            .O(N__22623),
            .I(n12785));
    CascadeMux I__2135 (
            .O(N__22620),
            .I(N__22617));
    InMux I__2134 (
            .O(N__22617),
            .I(N__22613));
    InMux I__2133 (
            .O(N__22616),
            .I(N__22610));
    LocalMux I__2132 (
            .O(N__22613),
            .I(n2719));
    LocalMux I__2131 (
            .O(N__22610),
            .I(n2719));
    InMux I__2130 (
            .O(N__22605),
            .I(N__22602));
    LocalMux I__2129 (
            .O(N__22602),
            .I(n2786));
    InMux I__2128 (
            .O(N__22599),
            .I(n12786));
    InMux I__2127 (
            .O(N__22596),
            .I(N__22593));
    LocalMux I__2126 (
            .O(N__22593),
            .I(n2785));
    InMux I__2125 (
            .O(N__22590),
            .I(bfn_2_25_0_));
    CascadeMux I__2124 (
            .O(N__22587),
            .I(N__22584));
    InMux I__2123 (
            .O(N__22584),
            .I(N__22581));
    LocalMux I__2122 (
            .O(N__22581),
            .I(n2784));
    InMux I__2121 (
            .O(N__22578),
            .I(n12788));
    InMux I__2120 (
            .O(N__22575),
            .I(N__22572));
    LocalMux I__2119 (
            .O(N__22572),
            .I(n2783));
    InMux I__2118 (
            .O(N__22569),
            .I(n12789));
    InMux I__2117 (
            .O(N__22566),
            .I(N__22563));
    LocalMux I__2116 (
            .O(N__22563),
            .I(n2782));
    InMux I__2115 (
            .O(N__22560),
            .I(n12790));
    InMux I__2114 (
            .O(N__22557),
            .I(N__22554));
    LocalMux I__2113 (
            .O(N__22554),
            .I(N__22551));
    Odrv4 I__2112 (
            .O(N__22551),
            .I(n2798));
    InMux I__2111 (
            .O(N__22548),
            .I(n12774));
    InMux I__2110 (
            .O(N__22545),
            .I(N__22542));
    LocalMux I__2109 (
            .O(N__22542),
            .I(N__22539));
    Odrv4 I__2108 (
            .O(N__22539),
            .I(n2797));
    InMux I__2107 (
            .O(N__22536),
            .I(n12775));
    InMux I__2106 (
            .O(N__22533),
            .I(n12776));
    InMux I__2105 (
            .O(N__22530),
            .I(n12777));
    InMux I__2104 (
            .O(N__22527),
            .I(n12778));
    InMux I__2103 (
            .O(N__22524),
            .I(bfn_2_24_0_));
    InMux I__2102 (
            .O(N__22521),
            .I(n12780));
    InMux I__2101 (
            .O(N__22518),
            .I(n12781));
    InMux I__2100 (
            .O(N__22515),
            .I(n12782));
    InMux I__2099 (
            .O(N__22512),
            .I(N__22509));
    LocalMux I__2098 (
            .O(N__22509),
            .I(n2586));
    CascadeMux I__2097 (
            .O(N__22506),
            .I(N__22503));
    InMux I__2096 (
            .O(N__22503),
            .I(N__22500));
    LocalMux I__2095 (
            .O(N__22500),
            .I(N__22496));
    InMux I__2094 (
            .O(N__22499),
            .I(N__22493));
    Span4Mux_v I__2093 (
            .O(N__22496),
            .I(N__22487));
    LocalMux I__2092 (
            .O(N__22493),
            .I(N__22487));
    InMux I__2091 (
            .O(N__22492),
            .I(N__22484));
    Span4Mux_v I__2090 (
            .O(N__22487),
            .I(N__22481));
    LocalMux I__2089 (
            .O(N__22484),
            .I(N__22478));
    Odrv4 I__2088 (
            .O(N__22481),
            .I(n2519));
    Odrv4 I__2087 (
            .O(N__22478),
            .I(n2519));
    InMux I__2086 (
            .O(N__22473),
            .I(N__22470));
    LocalMux I__2085 (
            .O(N__22470),
            .I(N__22467));
    Span4Mux_v I__2084 (
            .O(N__22467),
            .I(N__22464));
    Odrv4 I__2083 (
            .O(N__22464),
            .I(n2484));
    InMux I__2082 (
            .O(N__22461),
            .I(N__22458));
    LocalMux I__2081 (
            .O(N__22458),
            .I(n2583));
    CascadeMux I__2080 (
            .O(N__22455),
            .I(n2516_cascade_));
    InMux I__2079 (
            .O(N__22452),
            .I(N__22449));
    LocalMux I__2078 (
            .O(N__22449),
            .I(n2588));
    CascadeMux I__2077 (
            .O(N__22446),
            .I(N__22443));
    InMux I__2076 (
            .O(N__22443),
            .I(N__22440));
    LocalMux I__2075 (
            .O(N__22440),
            .I(n2580));
    CascadeMux I__2074 (
            .O(N__22437),
            .I(n2612_cascade_));
    CascadeMux I__2073 (
            .O(N__22434),
            .I(N__22431));
    InMux I__2072 (
            .O(N__22431),
            .I(N__22428));
    LocalMux I__2071 (
            .O(N__22428),
            .I(N__22425));
    Sp12to4 I__2070 (
            .O(N__22425),
            .I(N__22422));
    Odrv12 I__2069 (
            .O(N__22422),
            .I(n2801));
    InMux I__2068 (
            .O(N__22419),
            .I(bfn_2_23_0_));
    InMux I__2067 (
            .O(N__22416),
            .I(n12772));
    InMux I__2066 (
            .O(N__22413),
            .I(N__22410));
    LocalMux I__2065 (
            .O(N__22410),
            .I(N__22407));
    Odrv4 I__2064 (
            .O(N__22407),
            .I(n2799));
    InMux I__2063 (
            .O(N__22404),
            .I(n12773));
    CascadeMux I__2062 (
            .O(N__22401),
            .I(n14650_cascade_));
    InMux I__2061 (
            .O(N__22398),
            .I(N__22395));
    LocalMux I__2060 (
            .O(N__22395),
            .I(n2595));
    CascadeMux I__2059 (
            .O(N__22392),
            .I(N__22389));
    InMux I__2058 (
            .O(N__22389),
            .I(N__22385));
    InMux I__2057 (
            .O(N__22388),
            .I(N__22382));
    LocalMux I__2056 (
            .O(N__22385),
            .I(N__22378));
    LocalMux I__2055 (
            .O(N__22382),
            .I(N__22375));
    InMux I__2054 (
            .O(N__22381),
            .I(N__22372));
    Odrv12 I__2053 (
            .O(N__22378),
            .I(n2528));
    Odrv4 I__2052 (
            .O(N__22375),
            .I(n2528));
    LocalMux I__2051 (
            .O(N__22372),
            .I(n2528));
    CascadeMux I__2050 (
            .O(N__22365),
            .I(n2627_cascade_));
    InMux I__2049 (
            .O(N__22362),
            .I(N__22359));
    LocalMux I__2048 (
            .O(N__22359),
            .I(n14646));
    InMux I__2047 (
            .O(N__22356),
            .I(N__22352));
    InMux I__2046 (
            .O(N__22355),
            .I(N__22349));
    LocalMux I__2045 (
            .O(N__22352),
            .I(N__22343));
    LocalMux I__2044 (
            .O(N__22349),
            .I(N__22343));
    InMux I__2043 (
            .O(N__22348),
            .I(N__22340));
    Odrv4 I__2042 (
            .O(N__22343),
            .I(n2520));
    LocalMux I__2041 (
            .O(N__22340),
            .I(n2520));
    CascadeMux I__2040 (
            .O(N__22335),
            .I(N__22332));
    InMux I__2039 (
            .O(N__22332),
            .I(N__22329));
    LocalMux I__2038 (
            .O(N__22329),
            .I(n2587));
    InMux I__2037 (
            .O(N__22326),
            .I(N__22323));
    LocalMux I__2036 (
            .O(N__22323),
            .I(n2589));
    InMux I__2035 (
            .O(N__22320),
            .I(N__22316));
    InMux I__2034 (
            .O(N__22319),
            .I(N__22313));
    LocalMux I__2033 (
            .O(N__22316),
            .I(N__22307));
    LocalMux I__2032 (
            .O(N__22313),
            .I(N__22307));
    InMux I__2031 (
            .O(N__22312),
            .I(N__22304));
    Odrv4 I__2030 (
            .O(N__22307),
            .I(n2522));
    LocalMux I__2029 (
            .O(N__22304),
            .I(n2522));
    InMux I__2028 (
            .O(N__22299),
            .I(N__22296));
    LocalMux I__2027 (
            .O(N__22296),
            .I(N__22293));
    Odrv4 I__2026 (
            .O(N__22293),
            .I(n2596));
    CascadeMux I__2025 (
            .O(N__22290),
            .I(n2628_cascade_));
    InMux I__2024 (
            .O(N__22287),
            .I(N__22284));
    LocalMux I__2023 (
            .O(N__22284),
            .I(n14644));
    InMux I__2022 (
            .O(N__22281),
            .I(N__22277));
    CascadeMux I__2021 (
            .O(N__22280),
            .I(N__22274));
    LocalMux I__2020 (
            .O(N__22277),
            .I(N__22271));
    InMux I__2019 (
            .O(N__22274),
            .I(N__22268));
    Odrv12 I__2018 (
            .O(N__22271),
            .I(n2527));
    LocalMux I__2017 (
            .O(N__22268),
            .I(n2527));
    CascadeMux I__2016 (
            .O(N__22263),
            .I(N__22260));
    InMux I__2015 (
            .O(N__22260),
            .I(N__22257));
    LocalMux I__2014 (
            .O(N__22257),
            .I(N__22254));
    Odrv4 I__2013 (
            .O(N__22254),
            .I(n2594));
    InMux I__2012 (
            .O(N__22251),
            .I(N__22248));
    LocalMux I__2011 (
            .O(N__22248),
            .I(n2579));
    InMux I__2010 (
            .O(N__22245),
            .I(N__22242));
    LocalMux I__2009 (
            .O(N__22242),
            .I(N__22239));
    Odrv4 I__2008 (
            .O(N__22239),
            .I(n2491));
    CascadeMux I__2007 (
            .O(N__22236),
            .I(N__22233));
    InMux I__2006 (
            .O(N__22233),
            .I(N__22230));
    LocalMux I__2005 (
            .O(N__22230),
            .I(n2481));
    CascadeMux I__2004 (
            .O(N__22227),
            .I(N__22224));
    InMux I__2003 (
            .O(N__22224),
            .I(N__22221));
    LocalMux I__2002 (
            .O(N__22221),
            .I(n14310));
    CascadeMux I__2001 (
            .O(N__22218),
            .I(N__22215));
    InMux I__2000 (
            .O(N__22215),
            .I(N__22212));
    LocalMux I__1999 (
            .O(N__22212),
            .I(N__22209));
    Odrv4 I__1998 (
            .O(N__22209),
            .I(n2494));
    InMux I__1997 (
            .O(N__22206),
            .I(N__22203));
    LocalMux I__1996 (
            .O(N__22203),
            .I(N__22200));
    Odrv4 I__1995 (
            .O(N__22200),
            .I(n2483));
    InMux I__1994 (
            .O(N__22197),
            .I(N__22192));
    InMux I__1993 (
            .O(N__22196),
            .I(N__22189));
    InMux I__1992 (
            .O(N__22195),
            .I(N__22186));
    LocalMux I__1991 (
            .O(N__22192),
            .I(n2416));
    LocalMux I__1990 (
            .O(N__22189),
            .I(n2416));
    LocalMux I__1989 (
            .O(N__22186),
            .I(n2416));
    InMux I__1988 (
            .O(N__22179),
            .I(N__22176));
    LocalMux I__1987 (
            .O(N__22176),
            .I(n2480));
    CascadeMux I__1986 (
            .O(N__22173),
            .I(N__22170));
    InMux I__1985 (
            .O(N__22170),
            .I(N__22167));
    LocalMux I__1984 (
            .O(N__22167),
            .I(n2482));
    CascadeMux I__1983 (
            .O(N__22164),
            .I(n2418_cascade_));
    InMux I__1982 (
            .O(N__22161),
            .I(N__22158));
    LocalMux I__1981 (
            .O(N__22158),
            .I(N__22155));
    Odrv4 I__1980 (
            .O(N__22155),
            .I(n2495));
    CascadeMux I__1979 (
            .O(N__22152),
            .I(n2428_cascade_));
    CascadeMux I__1978 (
            .O(N__22149),
            .I(n2527_cascade_));
    InMux I__1977 (
            .O(N__22146),
            .I(N__22143));
    LocalMux I__1976 (
            .O(N__22143),
            .I(n2488));
    CascadeMux I__1975 (
            .O(N__22140),
            .I(N__22137));
    InMux I__1974 (
            .O(N__22137),
            .I(N__22134));
    LocalMux I__1973 (
            .O(N__22134),
            .I(n2493));
    InMux I__1972 (
            .O(N__22131),
            .I(N__22128));
    LocalMux I__1971 (
            .O(N__22128),
            .I(n2490));
    CascadeMux I__1970 (
            .O(N__22125),
            .I(N__22121));
    InMux I__1969 (
            .O(N__22124),
            .I(N__22118));
    InMux I__1968 (
            .O(N__22121),
            .I(N__22115));
    LocalMux I__1967 (
            .O(N__22118),
            .I(n2418));
    LocalMux I__1966 (
            .O(N__22115),
            .I(n2418));
    CascadeMux I__1965 (
            .O(N__22110),
            .I(N__22107));
    InMux I__1964 (
            .O(N__22107),
            .I(N__22104));
    LocalMux I__1963 (
            .O(N__22104),
            .I(n2485));
    InMux I__1962 (
            .O(N__22101),
            .I(N__22098));
    LocalMux I__1961 (
            .O(N__22098),
            .I(n2498));
    InMux I__1960 (
            .O(N__22095),
            .I(N__22092));
    LocalMux I__1959 (
            .O(N__22092),
            .I(n2487));
    InMux I__1958 (
            .O(N__22089),
            .I(N__22086));
    LocalMux I__1957 (
            .O(N__22086),
            .I(n2497));
    InMux I__1956 (
            .O(N__22083),
            .I(N__22080));
    LocalMux I__1955 (
            .O(N__22080),
            .I(n2499));
    CascadeMux I__1954 (
            .O(N__22077),
            .I(N__22074));
    InMux I__1953 (
            .O(N__22074),
            .I(N__22071));
    LocalMux I__1952 (
            .O(N__22071),
            .I(n2496));
    InMux I__1951 (
            .O(N__22068),
            .I(\debounce.n13020 ));
    InMux I__1950 (
            .O(N__22065),
            .I(\debounce.n13021 ));
    InMux I__1949 (
            .O(N__22062),
            .I(\debounce.n13022 ));
    InMux I__1948 (
            .O(N__22059),
            .I(bfn_1_32_0_));
    InMux I__1947 (
            .O(N__22056),
            .I(\debounce.n13024 ));
    InMux I__1946 (
            .O(N__22053),
            .I(N__22050));
    LocalMux I__1945 (
            .O(N__22050),
            .I(n2501));
    InMux I__1944 (
            .O(N__22047),
            .I(N__22044));
    LocalMux I__1943 (
            .O(N__22044),
            .I(n2500));
    CascadeMux I__1942 (
            .O(N__22041),
            .I(n2433_cascade_));
    CascadeMux I__1941 (
            .O(N__22038),
            .I(n2532_cascade_));
    InMux I__1940 (
            .O(N__22035),
            .I(N__22032));
    LocalMux I__1939 (
            .O(N__22032),
            .I(N__22029));
    Odrv12 I__1938 (
            .O(N__22029),
            .I(n2900));
    CascadeMux I__1937 (
            .O(N__22026),
            .I(n2833_cascade_));
    CascadeMux I__1936 (
            .O(N__22023),
            .I(n2932_cascade_));
    InMux I__1935 (
            .O(N__22020),
            .I(N__22017));
    LocalMux I__1934 (
            .O(N__22017),
            .I(N__22014));
    Span4Mux_v I__1933 (
            .O(N__22014),
            .I(N__22011));
    Odrv4 I__1932 (
            .O(N__22011),
            .I(n2901));
    CascadeMux I__1931 (
            .O(N__22008),
            .I(n2933_cascade_));
    InMux I__1930 (
            .O(N__22005),
            .I(bfn_1_31_0_));
    InMux I__1929 (
            .O(N__22002),
            .I(\debounce.n13016 ));
    InMux I__1928 (
            .O(N__21999),
            .I(\debounce.n13017 ));
    InMux I__1927 (
            .O(N__21996),
            .I(\debounce.n13018 ));
    InMux I__1926 (
            .O(N__21993),
            .I(\debounce.n13019 ));
    InMux I__1925 (
            .O(N__21990),
            .I(n12818));
    InMux I__1924 (
            .O(N__21987),
            .I(n12819));
    InMux I__1923 (
            .O(N__21984),
            .I(bfn_1_29_0_));
    InMux I__1922 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__1921 (
            .O(N__21978),
            .I(N__21975));
    Odrv12 I__1920 (
            .O(N__21975),
            .I(n2876));
    InMux I__1919 (
            .O(N__21972),
            .I(n12821));
    InMux I__1918 (
            .O(N__21969),
            .I(n12822));
    InMux I__1917 (
            .O(N__21966),
            .I(N__21963));
    LocalMux I__1916 (
            .O(N__21963),
            .I(N__21960));
    Span4Mux_s1_h I__1915 (
            .O(N__21960),
            .I(N__21957));
    Odrv4 I__1914 (
            .O(N__21957),
            .I(n11956));
    InMux I__1913 (
            .O(N__21954),
            .I(N__21951));
    LocalMux I__1912 (
            .O(N__21951),
            .I(N__21948));
    Odrv12 I__1911 (
            .O(N__21948),
            .I(n2899));
    CascadeMux I__1910 (
            .O(N__21945),
            .I(N__21942));
    InMux I__1909 (
            .O(N__21942),
            .I(N__21939));
    LocalMux I__1908 (
            .O(N__21939),
            .I(N__21936));
    Span4Mux_s1_h I__1907 (
            .O(N__21936),
            .I(N__21932));
    InMux I__1906 (
            .O(N__21935),
            .I(N__21929));
    Odrv4 I__1905 (
            .O(N__21932),
            .I(n2833));
    LocalMux I__1904 (
            .O(N__21929),
            .I(n2833));
    InMux I__1903 (
            .O(N__21924),
            .I(n12809));
    InMux I__1902 (
            .O(N__21921),
            .I(n12810));
    InMux I__1901 (
            .O(N__21918),
            .I(n12811));
    InMux I__1900 (
            .O(N__21915),
            .I(bfn_1_28_0_));
    InMux I__1899 (
            .O(N__21912),
            .I(n12813));
    InMux I__1898 (
            .O(N__21909),
            .I(n12814));
    InMux I__1897 (
            .O(N__21906),
            .I(n12815));
    InMux I__1896 (
            .O(N__21903),
            .I(n12816));
    InMux I__1895 (
            .O(N__21900),
            .I(n12817));
    InMux I__1894 (
            .O(N__21897),
            .I(n12800));
    InMux I__1893 (
            .O(N__21894),
            .I(n12801));
    InMux I__1892 (
            .O(N__21891),
            .I(n12802));
    InMux I__1891 (
            .O(N__21888),
            .I(n12803));
    InMux I__1890 (
            .O(N__21885),
            .I(bfn_1_27_0_));
    InMux I__1889 (
            .O(N__21882),
            .I(n12805));
    InMux I__1888 (
            .O(N__21879),
            .I(n12806));
    InMux I__1887 (
            .O(N__21876),
            .I(n12807));
    InMux I__1886 (
            .O(N__21873),
            .I(n12808));
    CascadeMux I__1885 (
            .O(N__21870),
            .I(n13845_cascade_));
    InMux I__1884 (
            .O(N__21867),
            .I(N__21864));
    LocalMux I__1883 (
            .O(N__21864),
            .I(n14702));
    InMux I__1882 (
            .O(N__21861),
            .I(bfn_1_26_0_));
    InMux I__1881 (
            .O(N__21858),
            .I(n12797));
    InMux I__1880 (
            .O(N__21855),
            .I(n12798));
    InMux I__1879 (
            .O(N__21852),
            .I(n12799));
    CascadeMux I__1878 (
            .O(N__21849),
            .I(N__21846));
    InMux I__1877 (
            .O(N__21846),
            .I(N__21843));
    LocalMux I__1876 (
            .O(N__21843),
            .I(N__21840));
    Odrv12 I__1875 (
            .O(N__21840),
            .I(n2486));
    CascadeMux I__1874 (
            .O(N__21837),
            .I(n2816_cascade_));
    CascadeMux I__1873 (
            .O(N__21834),
            .I(n2829_cascade_));
    InMux I__1872 (
            .O(N__21831),
            .I(bfn_1_22_0_));
    InMux I__1871 (
            .O(N__21828),
            .I(n12741));
    InMux I__1870 (
            .O(N__21825),
            .I(n12742));
    InMux I__1869 (
            .O(N__21822),
            .I(n12743));
    InMux I__1868 (
            .O(N__21819),
            .I(n12744));
    InMux I__1867 (
            .O(N__21816),
            .I(n12745));
    InMux I__1866 (
            .O(N__21813),
            .I(n12746));
    InMux I__1865 (
            .O(N__21810),
            .I(n12747));
    CascadeMux I__1864 (
            .O(N__21807),
            .I(n2719_cascade_));
    InMux I__1863 (
            .O(N__21804),
            .I(n12731));
    InMux I__1862 (
            .O(N__21801),
            .I(bfn_1_21_0_));
    InMux I__1861 (
            .O(N__21798),
            .I(n12733));
    InMux I__1860 (
            .O(N__21795),
            .I(n12734));
    InMux I__1859 (
            .O(N__21792),
            .I(n12735));
    InMux I__1858 (
            .O(N__21789),
            .I(n12736));
    InMux I__1857 (
            .O(N__21786),
            .I(n12737));
    InMux I__1856 (
            .O(N__21783),
            .I(n12738));
    InMux I__1855 (
            .O(N__21780),
            .I(n12739));
    InMux I__1854 (
            .O(N__21777),
            .I(n12723));
    InMux I__1853 (
            .O(N__21774),
            .I(n12724));
    InMux I__1852 (
            .O(N__21771),
            .I(bfn_1_20_0_));
    InMux I__1851 (
            .O(N__21768),
            .I(n12725));
    InMux I__1850 (
            .O(N__21765),
            .I(n12726));
    InMux I__1849 (
            .O(N__21762),
            .I(n12727));
    InMux I__1848 (
            .O(N__21759),
            .I(n12728));
    InMux I__1847 (
            .O(N__21756),
            .I(n12729));
    InMux I__1846 (
            .O(N__21753),
            .I(n12730));
    InMux I__1845 (
            .O(N__21750),
            .I(n12714));
    InMux I__1844 (
            .O(N__21747),
            .I(n12715));
    InMux I__1843 (
            .O(N__21744),
            .I(n12716));
    InMux I__1842 (
            .O(N__21741),
            .I(n12717));
    InMux I__1841 (
            .O(N__21738),
            .I(bfn_1_19_0_));
    InMux I__1840 (
            .O(N__21735),
            .I(n12719));
    InMux I__1839 (
            .O(N__21732),
            .I(n12720));
    InMux I__1838 (
            .O(N__21729),
            .I(n12721));
    InMux I__1837 (
            .O(N__21726),
            .I(n12722));
    InMux I__1836 (
            .O(N__21723),
            .I(n12705));
    InMux I__1835 (
            .O(N__21720),
            .I(n12706));
    InMux I__1834 (
            .O(N__21717),
            .I(n12707));
    InMux I__1833 (
            .O(N__21714),
            .I(n12708));
    InMux I__1832 (
            .O(N__21711),
            .I(n12709));
    InMux I__1831 (
            .O(N__21708),
            .I(bfn_1_18_0_));
    InMux I__1830 (
            .O(N__21705),
            .I(n12711));
    InMux I__1829 (
            .O(N__21702),
            .I(n12712));
    InMux I__1828 (
            .O(N__21699),
            .I(n12713));
    InMux I__1827 (
            .O(N__21696),
            .I(bfn_1_17_0_));
    InMux I__1826 (
            .O(N__21693),
            .I(n12703));
    InMux I__1825 (
            .O(N__21690),
            .I(n12704));
    IoInMux I__1824 (
            .O(N__21687),
            .I(N__21684));
    LocalMux I__1823 (
            .O(N__21684),
            .I(N__21681));
    IoSpan4Mux I__1822 (
            .O(N__21681),
            .I(N__21678));
    IoSpan4Mux I__1821 (
            .O(N__21678),
            .I(N__21675));
    IoSpan4Mux I__1820 (
            .O(N__21675),
            .I(N__21672));
    Odrv4 I__1819 (
            .O(N__21672),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_7_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_29_0_));
    defparam IN_MUX_bfv_7_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_30_0_ (
            .carryinitin(n12914),
            .carryinitout(bfn_7_30_0_));
    defparam IN_MUX_bfv_7_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_31_0_ (
            .carryinitin(n12922),
            .carryinitout(bfn_7_31_0_));
    defparam IN_MUX_bfv_7_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_32_0_ (
            .carryinitin(n12930),
            .carryinitout(bfn_7_32_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(n12442),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(n12450),
            .carryinitout(bfn_15_27_0_));
    defparam IN_MUX_bfv_15_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_28_0_ (
            .carryinitin(n12458),
            .carryinitout(bfn_15_28_0_));
    defparam IN_MUX_bfv_9_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_30_0_));
    defparam IN_MUX_bfv_9_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_31_0_ (
            .carryinitin(n12419),
            .carryinitout(bfn_9_31_0_));
    defparam IN_MUX_bfv_9_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_32_0_ (
            .carryinitin(n12427),
            .carryinitout(bfn_9_32_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_17_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_27_0_ (
            .carryinitin(n13006),
            .carryinitout(bfn_17_27_0_));
    defparam IN_MUX_bfv_17_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_28_0_ (
            .carryinitin(n13014),
            .carryinitout(bfn_17_28_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(\quad_counter0.n13032 ),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\quad_counter0.n13040 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(\quad_counter0.n13048 ),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_12_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_26_0_));
    defparam IN_MUX_bfv_12_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_27_0_ (
            .carryinitin(n12466),
            .carryinitout(bfn_12_27_0_));
    defparam IN_MUX_bfv_12_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_28_0_ (
            .carryinitin(n12474),
            .carryinitout(bfn_12_28_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(n12975),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(n12983),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(n12991),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(n12545),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(n12534),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(n12524),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(n12515),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(n12507),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_5_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_26_0_ (
            .carryinitin(n12885),
            .carryinitout(bfn_5_26_0_));
    defparam IN_MUX_bfv_5_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_27_0_ (
            .carryinitin(n12893),
            .carryinitout(bfn_5_27_0_));
    defparam IN_MUX_bfv_5_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_28_0_ (
            .carryinitin(n12901),
            .carryinitout(bfn_5_28_0_));
    defparam IN_MUX_bfv_3_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_29_0_));
    defparam IN_MUX_bfv_3_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_30_0_ (
            .carryinitin(n12857),
            .carryinitout(bfn_3_30_0_));
    defparam IN_MUX_bfv_3_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_31_0_ (
            .carryinitin(n12865),
            .carryinitout(bfn_3_31_0_));
    defparam IN_MUX_bfv_3_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_32_0_ (
            .carryinitin(n12873),
            .carryinitout(bfn_3_32_0_));
    defparam IN_MUX_bfv_2_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_29_0_));
    defparam IN_MUX_bfv_2_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_30_0_ (
            .carryinitin(n12830),
            .carryinitout(bfn_2_30_0_));
    defparam IN_MUX_bfv_2_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_31_0_ (
            .carryinitin(n12838),
            .carryinitout(bfn_2_31_0_));
    defparam IN_MUX_bfv_2_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_32_0_ (
            .carryinitin(n12846),
            .carryinitout(bfn_2_32_0_));
    defparam IN_MUX_bfv_1_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_26_0_));
    defparam IN_MUX_bfv_1_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_27_0_ (
            .carryinitin(n12804),
            .carryinitout(bfn_1_27_0_));
    defparam IN_MUX_bfv_1_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_28_0_ (
            .carryinitin(n12812),
            .carryinitout(bfn_1_28_0_));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(n12820),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(n12779),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(n12787),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(n12795),
            .carryinitout(bfn_2_26_0_));
    defparam IN_MUX_bfv_4_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_21_0_));
    defparam IN_MUX_bfv_4_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_22_0_ (
            .carryinitin(n12755),
            .carryinitout(bfn_4_22_0_));
    defparam IN_MUX_bfv_4_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_23_0_ (
            .carryinitin(n12763),
            .carryinitout(bfn_4_23_0_));
    defparam IN_MUX_bfv_4_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_24_0_ (
            .carryinitin(n12771),
            .carryinitout(bfn_4_24_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(n12732),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(n12740),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(n12710),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(n12718),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(n12689),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(n12697),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_5_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_20_0_));
    defparam IN_MUX_bfv_5_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_21_0_ (
            .carryinitin(n12669),
            .carryinitout(bfn_5_21_0_));
    defparam IN_MUX_bfv_5_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_22_0_ (
            .carryinitin(n12677),
            .carryinitout(bfn_5_22_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(n12650),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_5_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_19_0_ (
            .carryinitin(n12658),
            .carryinitout(bfn_5_19_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_7_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_18_0_ (
            .carryinitin(n12632),
            .carryinitout(bfn_7_18_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(n12640),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(n12615),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(n12623),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(n12599),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(n12607),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(n12584),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(n12570),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(n12557),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_15_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_31_0_));
    defparam IN_MUX_bfv_1_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_31_0_));
    defparam IN_MUX_bfv_1_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_32_0_ (
            .carryinitin(\debounce.n13023 ),
            .carryinitout(bfn_1_32_0_));
    defparam IN_MUX_bfv_11_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_29_0_));
    defparam IN_MUX_bfv_11_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_30_0_ (
            .carryinitin(n13094),
            .carryinitout(bfn_11_30_0_));
    defparam IN_MUX_bfv_11_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_31_0_ (
            .carryinitin(n13102),
            .carryinitout(bfn_11_31_0_));
    defparam IN_MUX_bfv_11_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_32_0_ (
            .carryinitin(n13110),
            .carryinitout(bfn_11_32_0_));
    defparam IN_MUX_bfv_7_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_23_0_));
    defparam IN_MUX_bfv_7_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_24_0_ (
            .carryinitin(n12945),
            .carryinitout(bfn_7_24_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(n12953),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_12_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_27_0_ (
            .carryinitin(\PWM.n13063 ),
            .carryinitout(bfn_13_27_0_));
    defparam IN_MUX_bfv_13_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_28_0_ (
            .carryinitin(\PWM.n13071 ),
            .carryinitout(bfn_13_28_0_));
    defparam IN_MUX_bfv_13_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_29_0_ (
            .carryinitin(\PWM.n13079 ),
            .carryinitout(bfn_13_29_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21687),
            .GLOBALBUFFEROUTPUT(CLK_N));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_1_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_1_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_1_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_2_lut_LC_1_17_0 (
            .in0(_gnd_net_),
            .in1(N__37816),
            .in2(_gnd_net_),
            .in3(N__21696),
            .lcout(n2501),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(n12703),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_1_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_1_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_1_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_3_lut_LC_1_17_1 (
            .in0(_gnd_net_),
            .in1(N__53441),
            .in2(N__23211),
            .in3(N__21693),
            .lcout(n2500),
            .ltout(),
            .carryin(n12703),
            .carryout(n12704),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_1_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_1_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_1_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_4_lut_LC_1_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23232),
            .in3(N__21690),
            .lcout(n2499),
            .ltout(),
            .carryin(n12704),
            .carryout(n12705),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_1_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_1_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_1_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_5_lut_LC_1_17_3 (
            .in0(_gnd_net_),
            .in1(N__23191),
            .in2(N__53813),
            .in3(N__21723),
            .lcout(n2498),
            .ltout(),
            .carryin(n12705),
            .carryout(n12706),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_1_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_1_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_1_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_6_lut_LC_1_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23174),
            .in3(N__21720),
            .lcout(n2497),
            .ltout(),
            .carryin(n12706),
            .carryout(n12707),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_1_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_1_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_1_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_7_lut_LC_1_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23148),
            .in3(N__21717),
            .lcout(n2496),
            .ltout(),
            .carryin(n12707),
            .carryout(n12708),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_1_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_1_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_1_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_8_lut_LC_1_17_6 (
            .in0(_gnd_net_),
            .in1(N__23076),
            .in2(N__53812),
            .in3(N__21714),
            .lcout(n2495),
            .ltout(),
            .carryin(n12708),
            .carryout(n12709),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_1_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_1_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_1_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_9_lut_LC_1_17_7 (
            .in0(_gnd_net_),
            .in1(N__53445),
            .in2(N__23124),
            .in3(N__21711),
            .lcout(n2494),
            .ltout(),
            .carryin(n12709),
            .carryout(n12710),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_1_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_1_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_1_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_10_lut_LC_1_18_0 (
            .in0(_gnd_net_),
            .in1(N__53433),
            .in2(N__23376),
            .in3(N__21708),
            .lcout(n2493),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(n12711),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_1_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_1_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_1_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_11_lut_LC_1_18_1 (
            .in0(_gnd_net_),
            .in1(N__53437),
            .in2(N__25689),
            .in3(N__21705),
            .lcout(n2492),
            .ltout(),
            .carryin(n12711),
            .carryout(n12712),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_1_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_1_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_1_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_12_lut_LC_1_18_2 (
            .in0(_gnd_net_),
            .in1(N__53434),
            .in2(N__23102),
            .in3(N__21702),
            .lcout(n2491),
            .ltout(),
            .carryin(n12712),
            .carryout(n12713),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_1_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_1_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_1_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_13_lut_LC_1_18_3 (
            .in0(_gnd_net_),
            .in1(N__53438),
            .in2(N__23631),
            .in3(N__21699),
            .lcout(n2490),
            .ltout(),
            .carryin(n12713),
            .carryout(n12714),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_1_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_1_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_1_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_14_lut_LC_1_18_4 (
            .in0(_gnd_net_),
            .in1(N__53435),
            .in2(N__23711),
            .in3(N__21750),
            .lcout(n2489),
            .ltout(),
            .carryin(n12714),
            .carryout(n12715),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_1_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_1_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_1_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_15_lut_LC_1_18_5 (
            .in0(_gnd_net_),
            .in1(N__53439),
            .in2(N__23352),
            .in3(N__21747),
            .lcout(n2488),
            .ltout(),
            .carryin(n12715),
            .carryout(n12716),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_1_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_1_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_1_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_16_lut_LC_1_18_6 (
            .in0(_gnd_net_),
            .in1(N__53436),
            .in2(N__23409),
            .in3(N__21744),
            .lcout(n2487),
            .ltout(),
            .carryin(n12716),
            .carryout(n12717),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_1_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_1_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_1_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_17_lut_LC_1_18_7 (
            .in0(_gnd_net_),
            .in1(N__53440),
            .in2(N__23598),
            .in3(N__21741),
            .lcout(n2486),
            .ltout(),
            .carryin(n12717),
            .carryout(n12718),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_1_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_1_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_1_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_18_lut_LC_1_19_0 (
            .in0(_gnd_net_),
            .in1(N__53418),
            .in2(N__22125),
            .in3(N__21738),
            .lcout(n2485),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(n12719),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_1_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_1_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_1_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_19_lut_LC_1_19_1 (
            .in0(_gnd_net_),
            .in1(N__53425),
            .in2(N__23537),
            .in3(N__21735),
            .lcout(n2484),
            .ltout(),
            .carryin(n12719),
            .carryout(n12720),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_1_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_1_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_1_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_20_lut_LC_1_19_2 (
            .in0(_gnd_net_),
            .in1(N__22196),
            .in2(N__53810),
            .in3(N__21732),
            .lcout(n2483),
            .ltout(),
            .carryin(n12720),
            .carryout(n12721),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_1_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_1_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_1_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_21_lut_LC_1_19_3 (
            .in0(_gnd_net_),
            .in1(N__23565),
            .in2(N__53808),
            .in3(N__21729),
            .lcout(n2482),
            .ltout(),
            .carryin(n12721),
            .carryout(n12722),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_1_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_1_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_1_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_22_lut_LC_1_19_4 (
            .in0(_gnd_net_),
            .in1(N__23508),
            .in2(N__53811),
            .in3(N__21726),
            .lcout(n2481),
            .ltout(),
            .carryin(n12722),
            .carryout(n12723),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_1_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_1_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_1_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_23_lut_LC_1_19_5 (
            .in0(_gnd_net_),
            .in1(N__23325),
            .in2(N__53809),
            .in3(N__21777),
            .lcout(n2480),
            .ltout(),
            .carryin(n12723),
            .carryout(n12724),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_1_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_1_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_1_19_6.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1637_24_lut_LC_1_19_6 (
            .in0(N__53432),
            .in1(N__33024),
            .in2(N__25521),
            .in3(N__21774),
            .lcout(n2511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_1_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_1_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_1_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_2_lut_LC_1_20_0 (
            .in0(_gnd_net_),
            .in1(N__28671),
            .in2(_gnd_net_),
            .in3(N__21771),
            .lcout(n2601),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(n12725),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_1_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_1_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_1_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_3_lut_LC_1_20_1 (
            .in0(_gnd_net_),
            .in1(N__53412),
            .in2(N__28637),
            .in3(N__21768),
            .lcout(n2600),
            .ltout(),
            .carryin(n12725),
            .carryout(n12726),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_1_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_1_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_1_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_4_lut_LC_1_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28586),
            .in3(N__21765),
            .lcout(n2599),
            .ltout(),
            .carryin(n12726),
            .carryout(n12727),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_1_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_1_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_1_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_5_lut_LC_1_20_3 (
            .in0(_gnd_net_),
            .in1(N__53413),
            .in2(N__24113),
            .in3(N__21762),
            .lcout(n2598),
            .ltout(),
            .carryin(n12727),
            .carryout(n12728),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_1_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_1_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_1_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_6_lut_LC_1_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23850),
            .in3(N__21759),
            .lcout(n2597),
            .ltout(),
            .carryin(n12728),
            .carryout(n12729),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_1_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_1_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_1_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_7_lut_LC_1_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23459),
            .in3(N__21756),
            .lcout(n2596),
            .ltout(),
            .carryin(n12729),
            .carryout(n12730),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_1_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_1_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_1_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_8_lut_LC_1_20_6 (
            .in0(_gnd_net_),
            .in1(N__22388),
            .in2(N__53807),
            .in3(N__21753),
            .lcout(n2595),
            .ltout(),
            .carryin(n12730),
            .carryout(n12731),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_1_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_1_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_1_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_9_lut_LC_1_20_7 (
            .in0(_gnd_net_),
            .in1(N__53417),
            .in2(N__22280),
            .in3(N__21804),
            .lcout(n2594),
            .ltout(),
            .carryin(n12731),
            .carryout(n12732),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_1_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_1_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_1_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_10_lut_LC_1_21_0 (
            .in0(_gnd_net_),
            .in1(N__54529),
            .in2(N__23658),
            .in3(N__21801),
            .lcout(n2593),
            .ltout(),
            .carryin(bfn_1_21_0_),
            .carryout(n12733),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_1_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_1_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_1_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_11_lut_LC_1_21_1 (
            .in0(_gnd_net_),
            .in1(N__54534),
            .in2(N__24188),
            .in3(N__21798),
            .lcout(n2592),
            .ltout(),
            .carryin(n12733),
            .carryout(n12734),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_1_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_1_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_1_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_12_lut_LC_1_21_2 (
            .in0(_gnd_net_),
            .in1(N__54530),
            .in2(N__25665),
            .in3(N__21795),
            .lcout(n2591),
            .ltout(),
            .carryin(n12734),
            .carryout(n12735),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_1_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_1_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_1_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_13_lut_LC_1_21_3 (
            .in0(_gnd_net_),
            .in1(N__54535),
            .in2(N__23892),
            .in3(N__21792),
            .lcout(n2590),
            .ltout(),
            .carryin(n12735),
            .carryout(n12736),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_1_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_1_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_1_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_14_lut_LC_1_21_4 (
            .in0(_gnd_net_),
            .in1(N__22319),
            .in2(N__54545),
            .in3(N__21789),
            .lcout(n2589),
            .ltout(),
            .carryin(n12736),
            .carryout(n12737),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_1_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_1_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_1_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_15_lut_LC_1_21_5 (
            .in0(_gnd_net_),
            .in1(N__54539),
            .in2(N__23676),
            .in3(N__21786),
            .lcout(n2588),
            .ltout(),
            .carryin(n12737),
            .carryout(n12738),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_1_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_1_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_1_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_16_lut_LC_1_21_6 (
            .in0(_gnd_net_),
            .in1(N__22355),
            .in2(N__54546),
            .in3(N__21783),
            .lcout(n2587),
            .ltout(),
            .carryin(n12738),
            .carryout(n12739),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_1_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_1_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_1_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_17_lut_LC_1_21_7 (
            .in0(_gnd_net_),
            .in1(N__22499),
            .in2(N__54544),
            .in3(N__21780),
            .lcout(n2586),
            .ltout(),
            .carryin(n12739),
            .carryout(n12740),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_1_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_1_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_1_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_18_lut_LC_1_22_0 (
            .in0(_gnd_net_),
            .in1(N__24016),
            .in2(N__54185),
            .in3(N__21831),
            .lcout(n2585),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(n12741),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_1_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_1_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_1_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_19_lut_LC_1_22_1 (
            .in0(_gnd_net_),
            .in1(N__53925),
            .in2(N__23766),
            .in3(N__21828),
            .lcout(n2584),
            .ltout(),
            .carryin(n12741),
            .carryout(n12742),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_1_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_1_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_1_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_20_lut_LC_1_22_2 (
            .in0(_gnd_net_),
            .in1(N__52886),
            .in2(N__23979),
            .in3(N__21825),
            .lcout(n2583),
            .ltout(),
            .carryin(n12742),
            .carryout(n12743),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_1_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_1_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_1_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_21_lut_LC_1_22_3 (
            .in0(_gnd_net_),
            .in1(N__53926),
            .in2(N__24143),
            .in3(N__21822),
            .lcout(n2582),
            .ltout(),
            .carryin(n12743),
            .carryout(n12744),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_1_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_1_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_1_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_22_lut_LC_1_22_4 (
            .in0(_gnd_net_),
            .in1(N__24287),
            .in2(N__54186),
            .in3(N__21819),
            .lcout(n2581),
            .ltout(),
            .carryin(n12744),
            .carryout(n12745),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_1_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_1_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_1_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_23_lut_LC_1_22_5 (
            .in0(_gnd_net_),
            .in1(N__23936),
            .in2(N__53195),
            .in3(N__21816),
            .lcout(n2580),
            .ltout(),
            .carryin(n12745),
            .carryout(n12746),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_1_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_1_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_1_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_24_lut_LC_1_22_6 (
            .in0(_gnd_net_),
            .in1(N__23962),
            .in2(N__54187),
            .in3(N__21813),
            .lcout(n2579),
            .ltout(),
            .carryin(n12746),
            .carryout(n12747),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_1_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_1_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_1_22_7.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1704_25_lut_LC_1_22_7 (
            .in0(N__52890),
            .in1(N__23912),
            .in2(N__33188),
            .in3(N__21810),
            .lcout(n2610),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_1_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_1_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_1_23_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1783_3_lut_LC_1_23_0 (
            .in0(_gnd_net_),
            .in1(N__26219),
            .in2(N__26199),
            .in3(N__33349),
            .lcout(n2719),
            .ltout(n2719_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_145_LC_1_23_1.C_ON=1'b0;
    defparam i1_3_lut_adj_145_LC_1_23_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_145_LC_1_23_1.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_145_LC_1_23_1 (
            .in0(_gnd_net_),
            .in1(N__24061),
            .in2(N__21807),
            .in3(N__24649),
            .lcout(n14138),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13096_1_lut_LC_1_23_2.C_ON=1'b0;
    defparam i13096_1_lut_LC_1_23_2.SEQ_MODE=4'b0000;
    defparam i13096_1_lut_LC_1_23_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 i13096_1_lut_LC_1_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33170),
            .lcout(n15821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_1_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_1_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_1_23_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1646_3_lut_LC_1_23_3 (
            .in0(_gnd_net_),
            .in1(N__23597),
            .in2(N__21849),
            .in3(N__33000),
            .lcout(n2518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i0_LC_1_23_5 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i0_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i0_LC_1_23_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \debounce.reg_out_i0_i0_LC_1_23_5  (
            .in0(N__47662),
            .in1(N__34854),
            .in2(_gnd_net_),
            .in3(N__39543),
            .lcout(h3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55773),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_1_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_1_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_1_24_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1908_3_lut_LC_1_24_1 (
            .in0(N__24897),
            .in1(N__21981),
            .in2(_gnd_net_),
            .in3(N__33713),
            .lcout(n2908),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_1_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_1_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_1_24_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1848_3_lut_LC_1_24_2 (
            .in0(_gnd_net_),
            .in1(N__24498),
            .in2(N__22587),
            .in3(N__33517),
            .lcout(n2816),
            .ltout(n2816_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_40_LC_1_24_3.C_ON=1'b0;
    defparam i1_4_lut_adj_40_LC_1_24_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_40_LC_1_24_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_40_LC_1_24_3 (
            .in0(N__26998),
            .in1(N__24985),
            .in2(N__21837),
            .in3(N__21867),
            .lcout(n14708),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_1_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_1_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_1_24_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1850_3_lut_LC_1_24_4 (
            .in0(_gnd_net_),
            .in1(N__22605),
            .in2(N__22620),
            .in3(N__33516),
            .lcout(n2818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_1_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_1_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_1_25_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1861_3_lut_LC_1_25_0 (
            .in0(_gnd_net_),
            .in1(N__26474),
            .in2(N__33522),
            .in3(N__22545),
            .lcout(n2829),
            .ltout(n2829_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_38_LC_1_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_38_LC_1_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_38_LC_1_25_1.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_38_LC_1_25_1 (
            .in0(N__24730),
            .in1(N__22864),
            .in2(N__21834),
            .in3(N__21966),
            .lcout(),
            .ltout(n13845_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_39_LC_1_25_2.C_ON=1'b0;
    defparam i1_4_lut_adj_39_LC_1_25_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_39_LC_1_25_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_39_LC_1_25_2 (
            .in0(N__27037),
            .in1(N__22912),
            .in2(N__21870),
            .in3(N__26577),
            .lcout(n14702),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_1_25_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_1_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_1_25_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1862_3_lut_LC_1_25_3 (
            .in0(_gnd_net_),
            .in1(N__22557),
            .in2(N__26514),
            .in3(N__33492),
            .lcout(n2830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_1_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_1_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_1_25_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1846_3_lut_LC_1_25_4 (
            .in0(N__24405),
            .in1(_gnd_net_),
            .in2(N__33523),
            .in3(N__22566),
            .lcout(n2814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_1_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_1_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_1_25_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1847_3_lut_LC_1_25_5 (
            .in0(N__22575),
            .in1(N__24435),
            .in2(_gnd_net_),
            .in3(N__33502),
            .lcout(n2815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_1_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_1_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_1_25_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1849_3_lut_LC_1_25_6 (
            .in0(N__24477),
            .in1(_gnd_net_),
            .in2(N__33521),
            .in3(N__22596),
            .lcout(n2817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_1_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_1_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_1_25_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1863_3_lut_LC_1_25_7 (
            .in0(_gnd_net_),
            .in1(N__22413),
            .in2(N__26901),
            .in3(N__33491),
            .lcout(n2831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_1_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_1_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_1_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_2_lut_LC_1_26_0 (
            .in0(_gnd_net_),
            .in1(N__38956),
            .in2(_gnd_net_),
            .in3(N__21861),
            .lcout(n2901),
            .ltout(),
            .carryin(bfn_1_26_0_),
            .carryout(n12797),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_1_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_1_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_1_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_3_lut_LC_1_26_1 (
            .in0(_gnd_net_),
            .in1(N__53028),
            .in2(N__21945),
            .in3(N__21858),
            .lcout(n2900),
            .ltout(),
            .carryin(n12797),
            .carryout(n12798),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_1_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_1_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_1_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_4_lut_LC_1_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22727),
            .in3(N__21855),
            .lcout(n2899),
            .ltout(),
            .carryin(n12798),
            .carryout(n12799),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_1_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_1_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_1_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_5_lut_LC_1_26_3 (
            .in0(_gnd_net_),
            .in1(N__53029),
            .in2(N__24737),
            .in3(N__21852),
            .lcout(n2898),
            .ltout(),
            .carryin(n12799),
            .carryout(n12800),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_1_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_1_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_1_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_6_lut_LC_1_26_4 (
            .in0(_gnd_net_),
            .in1(N__22865),
            .in2(_gnd_net_),
            .in3(N__21897),
            .lcout(n2897),
            .ltout(),
            .carryin(n12800),
            .carryout(n12801),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_1_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_1_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_1_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_7_lut_LC_1_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24680),
            .in3(N__21894),
            .lcout(n2896),
            .ltout(),
            .carryin(n12801),
            .carryout(n12802),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_1_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_1_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_1_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_8_lut_LC_1_26_6 (
            .in0(_gnd_net_),
            .in1(N__53031),
            .in2(N__27099),
            .in3(N__21891),
            .lcout(n2895),
            .ltout(),
            .carryin(n12802),
            .carryout(n12803),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_1_26_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_1_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_1_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_9_lut_LC_1_26_7 (
            .in0(_gnd_net_),
            .in1(N__53030),
            .in2(N__26787),
            .in3(N__21888),
            .lcout(n2894),
            .ltout(),
            .carryin(n12803),
            .carryout(n12804),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_1_27_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_1_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_1_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_10_lut_LC_1_27_0 (
            .in0(_gnd_net_),
            .in1(N__54415),
            .in2(N__25031),
            .in3(N__21885),
            .lcout(n2893),
            .ltout(),
            .carryin(bfn_1_27_0_),
            .carryout(n12805),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_1_27_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_1_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_1_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_11_lut_LC_1_27_1 (
            .in0(_gnd_net_),
            .in1(N__54422),
            .in2(N__27885),
            .in3(N__21882),
            .lcout(n2892),
            .ltout(),
            .carryin(n12805),
            .carryout(n12806),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_1_27_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_1_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_1_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_12_lut_LC_1_27_2 (
            .in0(_gnd_net_),
            .in1(N__54416),
            .in2(N__30710),
            .in3(N__21879),
            .lcout(n2891),
            .ltout(),
            .carryin(n12806),
            .carryout(n12807),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_1_27_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_1_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_1_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_13_lut_LC_1_27_3 (
            .in0(_gnd_net_),
            .in1(N__54423),
            .in2(N__24822),
            .in3(N__21876),
            .lcout(n2890),
            .ltout(),
            .carryin(n12807),
            .carryout(n12808),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_1_27_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_1_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_1_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_14_lut_LC_1_27_4 (
            .in0(_gnd_net_),
            .in1(N__54417),
            .in2(N__24540),
            .in3(N__21873),
            .lcout(n2889),
            .ltout(),
            .carryin(n12808),
            .carryout(n12809),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_1_27_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_1_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_1_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_15_lut_LC_1_27_5 (
            .in0(_gnd_net_),
            .in1(N__54424),
            .in2(N__24519),
            .in3(N__21924),
            .lcout(n2888),
            .ltout(),
            .carryin(n12809),
            .carryout(n12810),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_1_27_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_1_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_1_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_16_lut_LC_1_27_6 (
            .in0(_gnd_net_),
            .in1(N__54418),
            .in2(N__26616),
            .in3(N__21921),
            .lcout(n2887),
            .ltout(),
            .carryin(n12810),
            .carryout(n12811),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_1_27_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_1_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_1_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_17_lut_LC_1_27_7 (
            .in0(_gnd_net_),
            .in1(N__26826),
            .in2(N__54507),
            .in3(N__21918),
            .lcout(n2886),
            .ltout(),
            .carryin(n12811),
            .carryout(n12812),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_1_28_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_1_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_1_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_18_lut_LC_1_28_0 (
            .in0(_gnd_net_),
            .in1(N__27044),
            .in2(N__54508),
            .in3(N__21915),
            .lcout(n2885),
            .ltout(),
            .carryin(bfn_1_28_0_),
            .carryout(n12813),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_1_28_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_1_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_1_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_19_lut_LC_1_28_1 (
            .in0(_gnd_net_),
            .in1(N__22919),
            .in2(N__54512),
            .in3(N__21912),
            .lcout(n2884),
            .ltout(),
            .carryin(n12813),
            .carryout(n12814),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_1_28_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_1_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_1_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_20_lut_LC_1_28_2 (
            .in0(_gnd_net_),
            .in1(N__26282),
            .in2(N__54509),
            .in3(N__21909),
            .lcout(n2883),
            .ltout(),
            .carryin(n12814),
            .carryout(n12815),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_1_28_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_1_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_1_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_21_lut_LC_1_28_3 (
            .in0(_gnd_net_),
            .in1(N__24992),
            .in2(N__54513),
            .in3(N__21906),
            .lcout(n2882),
            .ltout(),
            .carryin(n12815),
            .carryout(n12816),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_1_28_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_1_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_1_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_22_lut_LC_1_28_4 (
            .in0(_gnd_net_),
            .in1(N__27005),
            .in2(N__54510),
            .in3(N__21903),
            .lcout(n2881),
            .ltout(),
            .carryin(n12816),
            .carryout(n12817),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_1_28_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_1_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_1_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_23_lut_LC_1_28_5 (
            .in0(_gnd_net_),
            .in1(N__24971),
            .in2(N__54514),
            .in3(N__21900),
            .lcout(n2880),
            .ltout(),
            .carryin(n12817),
            .carryout(n12818),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_1_28_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_1_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_1_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_24_lut_LC_1_28_6 (
            .in0(_gnd_net_),
            .in1(N__24704),
            .in2(N__54511),
            .in3(N__21990),
            .lcout(n2879),
            .ltout(),
            .carryin(n12818),
            .carryout(n12819),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_1_28_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_1_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_1_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_25_lut_LC_1_28_7 (
            .in0(_gnd_net_),
            .in1(N__22847),
            .in2(N__54515),
            .in3(N__21987),
            .lcout(n2878),
            .ltout(),
            .carryin(n12819),
            .carryout(n12820),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_1_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_1_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_1_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_26_lut_LC_1_29_0 (
            .in0(_gnd_net_),
            .in1(N__24872),
            .in2(N__54516),
            .in3(N__21984),
            .lcout(n2877),
            .ltout(),
            .carryin(bfn_1_29_0_),
            .carryout(n12821),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_1_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_1_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_1_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_27_lut_LC_1_29_1 (
            .in0(_gnd_net_),
            .in1(N__24896),
            .in2(N__54517),
            .in3(N__21972),
            .lcout(n2876),
            .ltout(),
            .carryin(n12821),
            .carryout(n12822),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_1_29_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_1_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_1_29_2.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1905_28_lut_LC_1_29_2 (
            .in0(N__24849),
            .in1(N__54455),
            .in2(N__33731),
            .in3(N__21969),
            .lcout(n2907),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9988_3_lut_LC_1_29_3.C_ON=1'b0;
    defparam i9988_3_lut_LC_1_29_3.SEQ_MODE=4'b0000;
    defparam i9988_3_lut_LC_1_29_3.LUT_INIT=16'b1100110010001000;
    LogicCell40 i9988_3_lut_LC_1_29_3 (
            .in0(N__38957),
            .in1(N__22723),
            .in2(_gnd_net_),
            .in3(N__21935),
            .lcout(n11956),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i1_LC_1_29_7 .C_ON=1'b0;
    defparam \debounce.reg_B_i1_LC_1_29_7 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i1_LC_1_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounce.reg_B_i1_LC_1_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34823),
            .lcout(reg_B_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55777),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_1_30_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_1_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_1_30_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1931_3_lut_LC_1_30_0 (
            .in0(_gnd_net_),
            .in1(N__21954),
            .in2(N__22731),
            .in3(N__33707),
            .lcout(n2931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_1_30_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_1_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_1_30_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1865_3_lut_LC_1_30_1 (
            .in0(_gnd_net_),
            .in1(N__44866),
            .in2(N__22434),
            .in3(N__33524),
            .lcout(n2833),
            .ltout(n2833_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_1_30_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_1_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_1_30_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1932_3_lut_LC_1_30_2 (
            .in0(_gnd_net_),
            .in1(N__22035),
            .in2(N__22026),
            .in3(N__33708),
            .lcout(n2932),
            .ltout(n2932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10070_4_lut_LC_1_30_3.C_ON=1'b0;
    defparam i10070_4_lut_LC_1_30_3.SEQ_MODE=4'b0000;
    defparam i10070_4_lut_LC_1_30_3.LUT_INIT=16'b1111110011101100;
    LogicCell40 i10070_4_lut_LC_1_30_3 (
            .in0(N__32432),
            .in1(N__27445),
            .in2(N__22023),
            .in3(N__22823),
            .lcout(n12038),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_1_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_1_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_1_30_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1933_3_lut_LC_1_30_6 (
            .in0(N__22020),
            .in1(_gnd_net_),
            .in2(N__38961),
            .in3(N__33706),
            .lcout(n2933),
            .ltout(n2933_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_1_30_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_1_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_1_30_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2000_3_lut_LC_1_30_7 (
            .in0(_gnd_net_),
            .in1(N__22812),
            .in2(N__22008),
            .in3(N__33886),
            .lcout(n3032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.cnt_reg_662__i0_LC_1_31_0 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i0_LC_1_31_0 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i0_LC_1_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i0_LC_1_31_0  (
            .in0(_gnd_net_),
            .in1(N__23034),
            .in2(_gnd_net_),
            .in3(N__22005),
            .lcout(\debounce.cnt_reg_0 ),
            .ltout(),
            .carryin(bfn_1_31_0_),
            .carryout(\debounce.n13016 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i1_LC_1_31_1 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i1_LC_1_31_1 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i1_LC_1_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i1_LC_1_31_1  (
            .in0(_gnd_net_),
            .in1(N__23009),
            .in2(_gnd_net_),
            .in3(N__22002),
            .lcout(\debounce.cnt_reg_1 ),
            .ltout(),
            .carryin(\debounce.n13016 ),
            .carryout(\debounce.n13017 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i2_LC_1_31_2 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i2_LC_1_31_2 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i2_LC_1_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i2_LC_1_31_2  (
            .in0(_gnd_net_),
            .in1(N__22995),
            .in2(_gnd_net_),
            .in3(N__21999),
            .lcout(\debounce.cnt_reg_2 ),
            .ltout(),
            .carryin(\debounce.n13017 ),
            .carryout(\debounce.n13018 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i3_LC_1_31_3 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i3_LC_1_31_3 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i3_LC_1_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i3_LC_1_31_3  (
            .in0(_gnd_net_),
            .in1(N__25154),
            .in2(_gnd_net_),
            .in3(N__21996),
            .lcout(\debounce.cnt_reg_3 ),
            .ltout(),
            .carryin(\debounce.n13018 ),
            .carryout(\debounce.n13019 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i4_LC_1_31_4 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i4_LC_1_31_4 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i4_LC_1_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i4_LC_1_31_4  (
            .in0(_gnd_net_),
            .in1(N__23267),
            .in2(_gnd_net_),
            .in3(N__21993),
            .lcout(\debounce.cnt_reg_4 ),
            .ltout(),
            .carryin(\debounce.n13019 ),
            .carryout(\debounce.n13020 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i5_LC_1_31_5 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i5_LC_1_31_5 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i5_LC_1_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i5_LC_1_31_5  (
            .in0(_gnd_net_),
            .in1(N__23253),
            .in2(_gnd_net_),
            .in3(N__22068),
            .lcout(\debounce.cnt_reg_5 ),
            .ltout(),
            .carryin(\debounce.n13020 ),
            .carryout(\debounce.n13021 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i6_LC_1_31_6 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i6_LC_1_31_6 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i6_LC_1_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i6_LC_1_31_6  (
            .in0(_gnd_net_),
            .in1(N__25181),
            .in2(_gnd_net_),
            .in3(N__22065),
            .lcout(\debounce.cnt_reg_6 ),
            .ltout(),
            .carryin(\debounce.n13021 ),
            .carryout(\debounce.n13022 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i7_LC_1_31_7 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i7_LC_1_31_7 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i7_LC_1_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i7_LC_1_31_7  (
            .in0(_gnd_net_),
            .in1(N__23022),
            .in2(_gnd_net_),
            .in3(N__22062),
            .lcout(\debounce.cnt_reg_7 ),
            .ltout(),
            .carryin(\debounce.n13022 ),
            .carryout(\debounce.n13023 ),
            .clk(N__55781),
            .ce(),
            .sr(N__27978));
    defparam \debounce.cnt_reg_662__i8_LC_1_32_0 .C_ON=1'b1;
    defparam \debounce.cnt_reg_662__i8_LC_1_32_0 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i8_LC_1_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i8_LC_1_32_0  (
            .in0(_gnd_net_),
            .in1(N__23286),
            .in2(_gnd_net_),
            .in3(N__22059),
            .lcout(\debounce.cnt_reg_8 ),
            .ltout(),
            .carryin(bfn_1_32_0_),
            .carryout(\debounce.n13024 ),
            .clk(N__55785),
            .ce(),
            .sr(N__27974));
    defparam \debounce.cnt_reg_662__i9_LC_1_32_1 .C_ON=1'b0;
    defparam \debounce.cnt_reg_662__i9_LC_1_32_1 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_662__i9_LC_1_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_662__i9_LC_1_32_1  (
            .in0(_gnd_net_),
            .in1(N__23298),
            .in2(_gnd_net_),
            .in3(N__22056),
            .lcout(\debounce.cnt_reg_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55785),
            .ce(),
            .sr(N__27974));
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_2_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_2_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_2_17_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1661_3_lut_LC_2_17_0 (
            .in0(N__37818),
            .in1(N__22053),
            .in2(_gnd_net_),
            .in3(N__32904),
            .lcout(n2533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_2_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_2_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_2_17_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1593_3_lut_LC_2_17_1 (
            .in0(N__30579),
            .in1(N__25134),
            .in2(_gnd_net_),
            .in3(N__32818),
            .lcout(n2433),
            .ltout(n2433_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_2_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_2_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_2_17_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1660_3_lut_LC_2_17_2 (
            .in0(_gnd_net_),
            .in1(N__22047),
            .in2(N__22041),
            .in3(N__32905),
            .lcout(n2532),
            .ltout(n2532_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9974_3_lut_LC_2_17_3.C_ON=1'b0;
    defparam i9974_3_lut_LC_2_17_3.SEQ_MODE=4'b0000;
    defparam i9974_3_lut_LC_2_17_3.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9974_3_lut_LC_2_17_3 (
            .in0(_gnd_net_),
            .in1(N__28670),
            .in2(N__22038),
            .in3(N__28618),
            .lcout(n11942),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_2_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_2_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_2_17_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1658_3_lut_LC_2_17_4 (
            .in0(_gnd_net_),
            .in1(N__22101),
            .in2(N__23196),
            .in3(N__32907),
            .lcout(n2530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_2_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_2_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_2_17_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1647_3_lut_LC_2_17_5 (
            .in0(N__23405),
            .in1(_gnd_net_),
            .in2(N__32952),
            .in3(N__22095),
            .lcout(n2519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_2_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_2_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_2_17_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1657_3_lut_LC_2_17_6 (
            .in0(_gnd_net_),
            .in1(N__22089),
            .in2(N__23175),
            .in3(N__32906),
            .lcout(n2529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_2_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_2_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_2_17_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1659_3_lut_LC_2_17_7 (
            .in0(_gnd_net_),
            .in1(N__22083),
            .in2(N__32953),
            .in3(N__23231),
            .lcout(n2531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_2_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_2_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_2_18_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1591_3_lut_LC_2_18_1 (
            .in0(_gnd_net_),
            .in1(N__30098),
            .in2(N__32820),
            .in3(N__25347),
            .lcout(n2431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_2_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_2_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_2_18_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1584_3_lut_LC_2_18_2 (
            .in0(_gnd_net_),
            .in1(N__28143),
            .in2(N__25215),
            .in3(N__32782),
            .lcout(n2424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_2_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_2_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_2_18_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1590_3_lut_LC_2_18_3 (
            .in0(_gnd_net_),
            .in1(N__28713),
            .in2(N__32821),
            .in3(N__25332),
            .lcout(n2430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_2_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_2_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_2_18_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1656_3_lut_LC_2_18_4 (
            .in0(_gnd_net_),
            .in1(N__23144),
            .in2(N__22077),
            .in3(N__32946),
            .lcout(n2528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_2_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_2_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_2_18_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1582_3_lut_LC_2_18_5 (
            .in0(_gnd_net_),
            .in1(N__29703),
            .in2(N__32819),
            .in3(N__25425),
            .lcout(n2422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_2_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_2_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_2_18_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1578_3_lut_LC_2_18_6 (
            .in0(_gnd_net_),
            .in1(N__25386),
            .in2(N__25599),
            .in3(N__32792),
            .lcout(n2418),
            .ltout(n2418_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_121_LC_2_18_7.C_ON=1'b0;
    defparam i1_4_lut_adj_121_LC_2_18_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_121_LC_2_18_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_121_LC_2_18_7 (
            .in0(N__23560),
            .in1(N__22195),
            .in2(N__22164),
            .in3(N__23604),
            .lcout(n14638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_2_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_2_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_2_19_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1588_3_lut_LC_2_19_0 (
            .in0(_gnd_net_),
            .in1(N__25278),
            .in2(N__25304),
            .in3(N__32768),
            .lcout(n2428),
            .ltout(n2428_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_2_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_2_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_2_19_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1655_3_lut_LC_2_19_1 (
            .in0(N__22161),
            .in1(_gnd_net_),
            .in2(N__22152),
            .in3(N__32941),
            .lcout(n2527),
            .ltout(n2527_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_127_LC_2_19_2.C_ON=1'b0;
    defparam i1_4_lut_adj_127_LC_2_19_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_127_LC_2_19_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_127_LC_2_19_2 (
            .in0(N__24174),
            .in1(N__22312),
            .in2(N__22149),
            .in3(N__22381),
            .lcout(n14310),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_2_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_2_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_2_19_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1576_3_lut_LC_2_19_3 (
            .in0(N__30247),
            .in1(_gnd_net_),
            .in2(N__32812),
            .in3(N__25365),
            .lcout(n2416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_2_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_2_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_2_19_4.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1648_3_lut_LC_2_19_4 (
            .in0(N__22146),
            .in1(_gnd_net_),
            .in2(N__32977),
            .in3(N__23351),
            .lcout(n2520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1653_3_lut_LC_2_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1653_3_lut_LC_2_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1653_3_lut_LC_2_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1653_3_lut_LC_2_19_5 (
            .in0(_gnd_net_),
            .in1(N__23372),
            .in2(N__22140),
            .in3(N__32940),
            .lcout(n2525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_2_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_2_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_2_19_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1650_3_lut_LC_2_19_6 (
            .in0(_gnd_net_),
            .in1(N__23627),
            .in2(N__32976),
            .in3(N__22131),
            .lcout(n2522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_2_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_2_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_2_19_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1645_3_lut_LC_2_19_7 (
            .in0(_gnd_net_),
            .in1(N__22124),
            .in2(N__22110),
            .in3(N__32945),
            .lcout(n2517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_2_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_2_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_2_20_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1651_3_lut_LC_2_20_0 (
            .in0(_gnd_net_),
            .in1(N__23103),
            .in2(N__32984),
            .in3(N__22245),
            .lcout(n2523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_2_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_2_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_2_20_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1641_3_lut_LC_2_20_1 (
            .in0(N__23506),
            .in1(_gnd_net_),
            .in2(N__22236),
            .in3(N__32965),
            .lcout(n2513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_128_LC_2_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_128_LC_2_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_128_LC_2_20_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_128_LC_2_20_2 (
            .in0(N__22348),
            .in1(N__22492),
            .in2(N__22227),
            .in3(N__23637),
            .lcout(n14318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_2_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_2_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_2_20_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1654_3_lut_LC_2_20_3 (
            .in0(_gnd_net_),
            .in1(N__23123),
            .in2(N__22218),
            .in3(N__32954),
            .lcout(n2526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_2_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_2_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_2_20_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1643_3_lut_LC_2_20_4 (
            .in0(_gnd_net_),
            .in1(N__22206),
            .in2(N__32986),
            .in3(N__22197),
            .lcout(n2515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1720_3_lut_LC_2_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1720_3_lut_LC_2_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1720_3_lut_LC_2_20_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1720_3_lut_LC_2_20_5 (
            .in0(_gnd_net_),
            .in1(N__24178),
            .in2(N__24209),
            .in3(N__33095),
            .lcout(n2624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_2_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_2_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_2_20_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1640_3_lut_LC_2_20_6 (
            .in0(_gnd_net_),
            .in1(N__22179),
            .in2(N__32985),
            .in3(N__23324),
            .lcout(n2512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_2_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_2_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_2_20_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1642_3_lut_LC_2_20_7 (
            .in0(_gnd_net_),
            .in1(N__23564),
            .in2(N__22173),
            .in3(N__32958),
            .lcout(n2514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_138_LC_2_21_0.C_ON=1'b0;
    defparam i1_4_lut_adj_138_LC_2_21_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_138_LC_2_21_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_138_LC_2_21_0 (
            .in0(N__25762),
            .in1(N__25729),
            .in2(N__26242),
            .in3(N__22287),
            .lcout(),
            .ltout(n14650_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_139_LC_2_21_1.C_ON=1'b0;
    defparam i1_4_lut_adj_139_LC_2_21_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_139_LC_2_21_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_139_LC_2_21_1 (
            .in0(N__26215),
            .in1(N__26173),
            .in2(N__22401),
            .in3(N__22362),
            .lcout(n14656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1723_3_lut_LC_2_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1723_3_lut_LC_2_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1723_3_lut_LC_2_21_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1723_3_lut_LC_2_21_2 (
            .in0(_gnd_net_),
            .in1(N__22398),
            .in2(N__22392),
            .in3(N__33135),
            .lcout(n2627),
            .ltout(n2627_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_137_LC_2_21_3.C_ON=1'b0;
    defparam i1_3_lut_adj_137_LC_2_21_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_137_LC_2_21_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_137_LC_2_21_3 (
            .in0(_gnd_net_),
            .in1(N__25858),
            .in2(N__22365),
            .in3(N__25828),
            .lcout(n14646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_2_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_2_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_2_21_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1715_3_lut_LC_2_21_4 (
            .in0(_gnd_net_),
            .in1(N__22356),
            .in2(N__22335),
            .in3(N__33136),
            .lcout(n2619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_2_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_2_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_2_21_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1717_3_lut_LC_2_21_5 (
            .in0(N__22326),
            .in1(_gnd_net_),
            .in2(N__33159),
            .in3(N__22320),
            .lcout(n2621),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_2_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_2_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_2_21_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1724_3_lut_LC_2_21_6 (
            .in0(_gnd_net_),
            .in1(N__22299),
            .in2(N__23466),
            .in3(N__33131),
            .lcout(n2628),
            .ltout(n2628_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_135_LC_2_21_7.C_ON=1'b0;
    defparam i1_2_lut_adj_135_LC_2_21_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_135_LC_2_21_7.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_135_LC_2_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22290),
            .in3(N__25796),
            .lcout(n14644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_2_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_2_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_2_22_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1722_3_lut_LC_2_22_0 (
            .in0(_gnd_net_),
            .in1(N__22281),
            .in2(N__22263),
            .in3(N__33121),
            .lcout(n2626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_2_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_2_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_2_22_1.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1707_3_lut_LC_2_22_1 (
            .in0(N__22251),
            .in1(_gnd_net_),
            .in2(N__33158),
            .in3(N__23963),
            .lcout(n2611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_2_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_2_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_2_22_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1714_3_lut_LC_2_22_2 (
            .in0(_gnd_net_),
            .in1(N__22512),
            .in2(N__22506),
            .in3(N__33125),
            .lcout(n2618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_2_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_2_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_2_22_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1644_3_lut_LC_2_22_3 (
            .in0(_gnd_net_),
            .in1(N__22473),
            .in2(N__23538),
            .in3(N__32997),
            .lcout(n2516),
            .ltout(n2516_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_2_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_2_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_2_22_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1711_3_lut_LC_2_22_4 (
            .in0(N__22461),
            .in1(_gnd_net_),
            .in2(N__22455),
            .in3(N__33126),
            .lcout(n2615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_2_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_2_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_2_22_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1716_3_lut_LC_2_22_5 (
            .in0(_gnd_net_),
            .in1(N__23672),
            .in2(N__33157),
            .in3(N__22452),
            .lcout(n2620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_2_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_2_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_2_22_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1708_3_lut_LC_2_22_6 (
            .in0(_gnd_net_),
            .in1(N__23937),
            .in2(N__22446),
            .in3(N__33127),
            .lcout(n2612),
            .ltout(n2612_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_2_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_2_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_2_22_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1775_3_lut_LC_2_22_7 (
            .in0(_gnd_net_),
            .in1(N__26391),
            .in2(N__22437),
            .in3(N__33344),
            .lcout(n2711),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_2_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_2_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_2_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_2_lut_LC_2_23_0 (
            .in0(_gnd_net_),
            .in1(N__44870),
            .in2(_gnd_net_),
            .in3(N__22419),
            .lcout(n2801),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(n12772),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_2_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_2_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_2_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_3_lut_LC_2_23_1 (
            .in0(_gnd_net_),
            .in1(N__53708),
            .in2(N__26928),
            .in3(N__22416),
            .lcout(n2800),
            .ltout(),
            .carryin(n12772),
            .carryout(n12773),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_2_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_2_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_2_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_4_lut_LC_2_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26893),
            .in3(N__22404),
            .lcout(n2799),
            .ltout(),
            .carryin(n12773),
            .carryout(n12774),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_2_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_2_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_2_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_5_lut_LC_2_23_3 (
            .in0(_gnd_net_),
            .in1(N__53709),
            .in2(N__26513),
            .in3(N__22548),
            .lcout(n2798),
            .ltout(),
            .carryin(n12774),
            .carryout(n12775),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_2_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_2_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_2_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_6_lut_LC_2_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26478),
            .in3(N__22536),
            .lcout(n2797),
            .ltout(),
            .carryin(n12775),
            .carryout(n12776),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_2_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_2_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_2_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_7_lut_LC_2_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26862),
            .in3(N__22533),
            .lcout(n2796),
            .ltout(),
            .carryin(n12776),
            .carryout(n12777),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_2_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_2_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_2_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_8_lut_LC_2_23_6 (
            .in0(_gnd_net_),
            .in1(N__24329),
            .in2(N__54009),
            .in3(N__22530),
            .lcout(n2795),
            .ltout(),
            .carryin(n12777),
            .carryout(n12778),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_2_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_2_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_2_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_9_lut_LC_2_23_7 (
            .in0(_gnd_net_),
            .in1(N__53713),
            .in2(N__24062),
            .in3(N__22527),
            .lcout(n2794),
            .ltout(),
            .carryin(n12778),
            .carryout(n12779),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_2_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_2_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_2_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_10_lut_LC_2_24_0 (
            .in0(_gnd_net_),
            .in1(N__53783),
            .in2(N__26718),
            .in3(N__22524),
            .lcout(n2793),
            .ltout(),
            .carryin(bfn_2_24_0_),
            .carryout(n12780),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_2_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_2_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_2_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_11_lut_LC_2_24_1 (
            .in0(_gnd_net_),
            .in1(N__53792),
            .in2(N__24650),
            .in3(N__22521),
            .lcout(n2792),
            .ltout(),
            .carryin(n12780),
            .carryout(n12781),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_2_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_2_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_2_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_12_lut_LC_2_24_2 (
            .in0(_gnd_net_),
            .in1(N__53784),
            .in2(N__26696),
            .in3(N__22518),
            .lcout(n2791),
            .ltout(),
            .carryin(n12781),
            .carryout(n12782),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_2_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_2_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_2_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_13_lut_LC_2_24_3 (
            .in0(_gnd_net_),
            .in1(N__53793),
            .in2(N__26669),
            .in3(N__22515),
            .lcout(n2790),
            .ltout(),
            .carryin(n12782),
            .carryout(n12783),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_2_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_2_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_2_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_14_lut_LC_2_24_4 (
            .in0(_gnd_net_),
            .in1(N__53785),
            .in2(N__24374),
            .in3(N__22629),
            .lcout(n2789),
            .ltout(),
            .carryin(n12783),
            .carryout(n12784),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_2_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_2_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_2_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_15_lut_LC_2_24_5 (
            .in0(_gnd_net_),
            .in1(N__24611),
            .in2(N__54079),
            .in3(N__22626),
            .lcout(n2788),
            .ltout(),
            .carryin(n12784),
            .carryout(n12785),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_2_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_2_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_2_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_16_lut_LC_2_24_6 (
            .in0(_gnd_net_),
            .in1(N__26735),
            .in2(N__54081),
            .in3(N__22623),
            .lcout(n2787),
            .ltout(),
            .carryin(n12785),
            .carryout(n12786),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_2_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_2_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_2_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_17_lut_LC_2_24_7 (
            .in0(_gnd_net_),
            .in1(N__22616),
            .in2(N__54080),
            .in3(N__22599),
            .lcout(n2786),
            .ltout(),
            .carryin(n12786),
            .carryout(n12787),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_2_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_2_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_2_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_18_lut_LC_2_25_0 (
            .in0(_gnd_net_),
            .in1(N__53616),
            .in2(N__24476),
            .in3(N__22590),
            .lcout(n2785),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(n12788),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_2_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_2_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_2_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_19_lut_LC_2_25_1 (
            .in0(_gnd_net_),
            .in1(N__24494),
            .in2(N__53981),
            .in3(N__22578),
            .lcout(n2784),
            .ltout(),
            .carryin(n12788),
            .carryout(n12789),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_2_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_2_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_2_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_20_lut_LC_2_25_2 (
            .in0(_gnd_net_),
            .in1(N__53620),
            .in2(N__24434),
            .in3(N__22569),
            .lcout(n2783),
            .ltout(),
            .carryin(n12789),
            .carryout(n12790),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_2_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_2_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_2_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_21_lut_LC_2_25_3 (
            .in0(_gnd_net_),
            .in1(N__24401),
            .in2(N__53982),
            .in3(N__22560),
            .lcout(n2782),
            .ltout(),
            .carryin(n12790),
            .carryout(n12791),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_2_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_2_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_2_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_22_lut_LC_2_25_4 (
            .in0(_gnd_net_),
            .in1(N__22757),
            .in2(N__53985),
            .in3(N__22662),
            .lcout(n2781),
            .ltout(),
            .carryin(n12791),
            .carryout(n12792),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_2_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_2_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_2_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_23_lut_LC_2_25_5 (
            .in0(_gnd_net_),
            .in1(N__24232),
            .in2(N__53983),
            .in3(N__22659),
            .lcout(n2780),
            .ltout(),
            .carryin(n12792),
            .carryout(n12793),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_2_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_2_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_2_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_24_lut_LC_2_25_6 (
            .in0(_gnd_net_),
            .in1(N__24310),
            .in2(N__53986),
            .in3(N__22656),
            .lcout(n2779),
            .ltout(),
            .carryin(n12793),
            .carryout(n12794),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_2_25_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_2_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_2_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_25_lut_LC_2_25_7 (
            .in0(_gnd_net_),
            .in1(N__22794),
            .in2(N__53984),
            .in3(N__22653),
            .lcout(n2778),
            .ltout(),
            .carryin(n12794),
            .carryout(n12795),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_2_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_2_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_2_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_26_lut_LC_2_26_0 (
            .in0(_gnd_net_),
            .in1(N__24911),
            .in2(N__53411),
            .in3(N__22650),
            .lcout(n2777),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(n12796),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_2_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_2_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_2_26_1.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1838_27_lut_LC_2_26_1 (
            .in0(N__54297),
            .in1(N__26298),
            .in2(N__33551),
            .in3(N__22647),
            .lcout(n2808),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_2_26_2.C_ON=1'b0;
    defparam i1_4_lut_LC_2_26_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_2_26_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_LC_2_26_2 (
            .in0(N__22756),
            .in1(N__24233),
            .in2(N__24312),
            .in3(N__24381),
            .lcout(),
            .ltout(n14158_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12589_4_lut_LC_2_26_3.C_ON=1'b0;
    defparam i12589_4_lut_LC_2_26_3.SEQ_MODE=4'b0000;
    defparam i12589_4_lut_LC_2_26_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12589_4_lut_LC_2_26_3 (
            .in0(N__24910),
            .in1(N__22792),
            .in2(N__22644),
            .in3(N__26297),
            .lcout(n2742),
            .ltout(n2742_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12449_3_lut_LC_2_26_4.C_ON=1'b0;
    defparam i12449_3_lut_LC_2_26_4.SEQ_MODE=4'b0000;
    defparam i12449_3_lut_LC_2_26_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 i12449_3_lut_LC_2_26_4 (
            .in0(_gnd_net_),
            .in1(N__22641),
            .in2(N__22632),
            .in3(N__26670),
            .lcout(n2822),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_2_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_2_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_2_26_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1853_3_lut_LC_2_26_5 (
            .in0(_gnd_net_),
            .in1(N__22803),
            .in2(N__24375),
            .in3(N__33456),
            .lcout(n2821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_2_26_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_2_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_2_26_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1842_3_lut_LC_2_26_6 (
            .in0(N__22793),
            .in1(_gnd_net_),
            .in2(N__33506),
            .in3(N__22776),
            .lcout(n2810),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_2_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_2_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_2_26_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1778_3_lut_LC_2_26_7 (
            .in0(N__26013),
            .in1(_gnd_net_),
            .in2(N__33351),
            .in3(N__26043),
            .lcout(n2714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_2_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_2_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_2_27_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1845_3_lut_LC_2_27_0 (
            .in0(N__22767),
            .in1(N__22758),
            .in2(_gnd_net_),
            .in3(N__33452),
            .lcout(n2813),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_2_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_2_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_2_27_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1864_3_lut_LC_2_27_1 (
            .in0(_gnd_net_),
            .in1(N__26927),
            .in2(N__33503),
            .in3(N__22740),
            .lcout(n2832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_2_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_2_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_2_27_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1858_3_lut_LC_2_27_2 (
            .in0(_gnd_net_),
            .in1(N__22701),
            .in2(N__24069),
            .in3(N__33445),
            .lcout(n2826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_2_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_2_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_2_27_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1919_3_lut_LC_2_27_3 (
            .in0(_gnd_net_),
            .in1(N__26609),
            .in2(N__22692),
            .in3(N__33647),
            .lcout(n2919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_2_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_2_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_2_27_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1843_3_lut_LC_2_27_5 (
            .in0(_gnd_net_),
            .in1(N__22683),
            .in2(N__33505),
            .in3(N__24311),
            .lcout(n2811),
            .ltout(n2811_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_41_LC_2_27_6.C_ON=1'b0;
    defparam i1_4_lut_adj_41_LC_2_27_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_41_LC_2_27_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_41_LC_2_27_6 (
            .in0(N__24703),
            .in1(N__24970),
            .in2(N__22674),
            .in3(N__22671),
            .lcout(n14714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_2_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_2_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_2_27_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1844_3_lut_LC_2_27_7 (
            .in0(_gnd_net_),
            .in1(N__24234),
            .in2(N__33504),
            .in3(N__22929),
            .lcout(n2812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_2_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_2_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_2_28_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1916_3_lut_LC_2_28_1 (
            .in0(_gnd_net_),
            .in1(N__22920),
            .in2(N__22896),
            .in3(N__33667),
            .lcout(n2916),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_2_28_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_2_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_2_28_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1909_3_lut_LC_2_28_2 (
            .in0(_gnd_net_),
            .in1(N__22887),
            .in2(N__33701),
            .in3(N__24873),
            .lcout(n2909),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_2_28_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_2_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_2_28_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1929_3_lut_LC_2_28_3 (
            .in0(_gnd_net_),
            .in1(N__22881),
            .in2(N__22872),
            .in3(N__33668),
            .lcout(n2929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_2_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_2_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_2_28_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2054_3_lut_LC_2_28_4 (
            .in0(N__27575),
            .in1(_gnd_net_),
            .in2(N__25110),
            .in3(N__37219),
            .lcout(n3118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12621_1_lut_LC_2_28_5.C_ON=1'b0;
    defparam i12621_1_lut_LC_2_28_5.SEQ_MODE=4'b0000;
    defparam i12621_1_lut_LC_2_28_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12621_1_lut_LC_2_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33669),
            .lcout(n15346),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_2_28_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_2_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_2_28_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1910_3_lut_LC_2_28_6 (
            .in0(_gnd_net_),
            .in1(N__22848),
            .in2(N__33700),
            .in3(N__22836),
            .lcout(n2910),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_2_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_2_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_2_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_2_lut_LC_2_29_0 (
            .in0(_gnd_net_),
            .in1(N__32433),
            .in2(_gnd_net_),
            .in3(N__22830),
            .lcout(n3001),
            .ltout(),
            .carryin(bfn_2_29_0_),
            .carryout(n12823),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_2_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_2_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_2_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_3_lut_LC_2_29_1 (
            .in0(_gnd_net_),
            .in1(N__53763),
            .in2(N__22827),
            .in3(N__22806),
            .lcout(n3000),
            .ltout(),
            .carryin(n12823),
            .carryout(n12824),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_2_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_2_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_2_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_4_lut_LC_2_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29417),
            .in3(N__22956),
            .lcout(n2999),
            .ltout(),
            .carryin(n12824),
            .carryout(n12825),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_2_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_2_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_2_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_5_lut_LC_2_29_3 (
            .in0(_gnd_net_),
            .in1(N__53764),
            .in2(N__27452),
            .in3(N__22953),
            .lcout(n2998),
            .ltout(),
            .carryin(n12825),
            .carryout(n12826),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_2_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_2_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_2_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_6_lut_LC_2_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27167),
            .in3(N__22950),
            .lcout(n2997),
            .ltout(),
            .carryin(n12826),
            .carryout(n12827),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_2_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_2_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_2_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_7_lut_LC_2_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27285),
            .in3(N__22947),
            .lcout(n2996),
            .ltout(),
            .carryin(n12827),
            .carryout(n12828),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_2_29_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_2_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_2_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_8_lut_LC_2_29_6 (
            .in0(_gnd_net_),
            .in1(N__54062),
            .in2(N__27198),
            .in3(N__22944),
            .lcout(n2995),
            .ltout(),
            .carryin(n12828),
            .carryout(n12829),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_2_29_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_2_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_2_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_9_lut_LC_2_29_7 (
            .in0(_gnd_net_),
            .in1(N__53765),
            .in2(N__27378),
            .in3(N__22941),
            .lcout(n2994),
            .ltout(),
            .carryin(n12829),
            .carryout(n12830),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_2_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_2_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_2_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_10_lut_LC_2_30_0 (
            .in0(_gnd_net_),
            .in1(N__54010),
            .in2(N__28917),
            .in3(N__22938),
            .lcout(n2993),
            .ltout(),
            .carryin(bfn_2_30_0_),
            .carryout(n12831),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_2_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_2_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_2_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_11_lut_LC_2_30_1 (
            .in0(_gnd_net_),
            .in1(N__54354),
            .in2(N__28986),
            .in3(N__22935),
            .lcout(n2992),
            .ltout(),
            .carryin(n12831),
            .carryout(n12832),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_2_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_2_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_2_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_12_lut_LC_2_30_2 (
            .in0(_gnd_net_),
            .in1(N__54011),
            .in2(N__27837),
            .in3(N__22932),
            .lcout(n2991),
            .ltout(),
            .carryin(n12832),
            .carryout(n12833),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_2_30_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_2_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_2_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_13_lut_LC_2_30_3 (
            .in0(_gnd_net_),
            .in1(N__30671),
            .in2(N__54262),
            .in3(N__22983),
            .lcout(n2990),
            .ltout(),
            .carryin(n12833),
            .carryout(n12834),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_2_30_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_2_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_2_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_14_lut_LC_2_30_4 (
            .in0(_gnd_net_),
            .in1(N__27551),
            .in2(N__54458),
            .in3(N__22980),
            .lcout(n2989),
            .ltout(),
            .carryin(n12834),
            .carryout(n12835),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_2_30_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_2_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_2_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_15_lut_LC_2_30_5 (
            .in0(_gnd_net_),
            .in1(N__27249),
            .in2(N__54263),
            .in3(N__22977),
            .lcout(n2988),
            .ltout(),
            .carryin(n12835),
            .carryout(n12836),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_2_30_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_2_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_2_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_16_lut_LC_2_30_6 (
            .in0(_gnd_net_),
            .in1(N__54018),
            .in2(N__24792),
            .in3(N__22974),
            .lcout(n2987),
            .ltout(),
            .carryin(n12836),
            .carryout(n12837),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_2_30_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_2_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_2_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_17_lut_LC_2_30_7 (
            .in0(_gnd_net_),
            .in1(N__54358),
            .in2(N__27686),
            .in3(N__22971),
            .lcout(n2986),
            .ltout(),
            .carryin(n12837),
            .carryout(n12838),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_2_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_2_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_2_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_18_lut_LC_2_31_0 (
            .in0(_gnd_net_),
            .in1(N__27933),
            .in2(N__54272),
            .in3(N__22968),
            .lcout(n2985),
            .ltout(),
            .carryin(bfn_2_31_0_),
            .carryout(n12839),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_2_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_2_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_2_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_19_lut_LC_2_31_1 (
            .in0(_gnd_net_),
            .in1(N__27482),
            .in2(N__54278),
            .in3(N__22965),
            .lcout(n2984),
            .ltout(),
            .carryin(n12839),
            .carryout(n12840),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_2_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_2_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_2_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_20_lut_LC_2_31_2 (
            .in0(_gnd_net_),
            .in1(N__29356),
            .in2(N__54273),
            .in3(N__22962),
            .lcout(n2983),
            .ltout(),
            .carryin(n12840),
            .carryout(n12841),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_2_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_2_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_2_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_21_lut_LC_2_31_3 (
            .in0(_gnd_net_),
            .in1(N__27762),
            .in2(N__54279),
            .in3(N__22959),
            .lcout(n2982),
            .ltout(),
            .carryin(n12841),
            .carryout(n12842),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_2_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_2_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_2_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_22_lut_LC_2_31_4 (
            .in0(_gnd_net_),
            .in1(N__27617),
            .in2(N__54274),
            .in3(N__23058),
            .lcout(n2981),
            .ltout(),
            .carryin(n12842),
            .carryout(n12843),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_2_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_2_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_2_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_23_lut_LC_2_31_5 (
            .in0(_gnd_net_),
            .in1(N__54052),
            .in2(N__27804),
            .in3(N__23055),
            .lcout(n2980),
            .ltout(),
            .carryin(n12843),
            .carryout(n12844),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_2_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_2_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_2_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_24_lut_LC_2_31_6 (
            .in0(_gnd_net_),
            .in1(N__27716),
            .in2(N__54275),
            .in3(N__23052),
            .lcout(n2979),
            .ltout(),
            .carryin(n12844),
            .carryout(n12845),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_2_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_2_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_2_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_25_lut_LC_2_31_7 (
            .in0(_gnd_net_),
            .in1(N__27911),
            .in2(N__54280),
            .in3(N__23049),
            .lcout(n2978),
            .ltout(),
            .carryin(n12845),
            .carryout(n12846),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_2_32_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_2_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_2_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_26_lut_LC_2_32_0 (
            .in0(_gnd_net_),
            .in1(N__28031),
            .in2(N__54283),
            .in3(N__23046),
            .lcout(n2977),
            .ltout(),
            .carryin(bfn_2_32_0_),
            .carryout(n12847),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_2_32_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_2_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_2_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_27_lut_LC_2_32_1 (
            .in0(_gnd_net_),
            .in1(N__27335),
            .in2(N__54285),
            .in3(N__23043),
            .lcout(n2976),
            .ltout(),
            .carryin(n12847),
            .carryout(n12848),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_2_32_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_2_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_2_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_28_lut_LC_2_32_2 (
            .in0(_gnd_net_),
            .in1(N__28086),
            .in2(N__54284),
            .in3(N__23040),
            .lcout(n2975),
            .ltout(),
            .carryin(n12848),
            .carryout(n12849),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_2_32_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_2_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_2_32_3.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1972_29_lut_LC_2_32_3 (
            .in0(N__54091),
            .in1(N__27311),
            .in2(N__32306),
            .in3(N__23037),
            .lcout(n3006),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i6_4_lut_LC_2_32_4 .C_ON=1'b0;
    defparam \debounce.i6_4_lut_LC_2_32_4 .SEQ_MODE=4'b0000;
    defparam \debounce.i6_4_lut_LC_2_32_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \debounce.i6_4_lut_LC_2_32_4  (
            .in0(N__23033),
            .in1(N__23021),
            .in2(N__23010),
            .in3(N__22994),
            .lcout(\debounce.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12653_1_lut_LC_2_32_5.C_ON=1'b0;
    defparam i12653_1_lut_LC_2_32_5.SEQ_MODE=4'b0000;
    defparam i12653_1_lut_LC_2_32_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12653_1_lut_LC_2_32_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33895),
            .lcout(n15378),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i7_4_lut_LC_2_32_6 .C_ON=1'b0;
    defparam \debounce.i7_4_lut_LC_2_32_6 .SEQ_MODE=4'b0000;
    defparam \debounce.i7_4_lut_LC_2_32_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \debounce.i7_4_lut_LC_2_32_6  (
            .in0(N__23297),
            .in1(N__23285),
            .in2(N__23274),
            .in3(N__23252),
            .lcout(\debounce.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_2_32_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_2_32_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_2_32_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1976_3_lut_LC_2_32_7 (
            .in0(_gnd_net_),
            .in1(N__27336),
            .in2(N__23241),
            .in3(N__33896),
            .lcout(n3008),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_3_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_3_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_3_17_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1592_3_lut_LC_3_17_0 (
            .in0(_gnd_net_),
            .in1(N__25122),
            .in2(N__28458),
            .in3(N__32813),
            .lcout(n2432),
            .ltout(n2432_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9978_3_lut_LC_3_17_1.C_ON=1'b0;
    defparam i9978_3_lut_LC_3_17_1.SEQ_MODE=4'b0000;
    defparam i9978_3_lut_LC_3_17_1.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9978_3_lut_LC_3_17_1 (
            .in0(_gnd_net_),
            .in1(N__37817),
            .in2(N__23214),
            .in3(N__23207),
            .lcout(),
            .ltout(n11946_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_114_LC_3_17_2.C_ON=1'b0;
    defparam i1_4_lut_adj_114_LC_3_17_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_114_LC_3_17_2.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_114_LC_3_17_2 (
            .in0(N__23192),
            .in1(N__23170),
            .in2(N__23151),
            .in3(N__23143),
            .lcout(n13816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_3_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_3_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_3_17_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1589_3_lut_LC_3_17_4 (
            .in0(N__29873),
            .in1(_gnd_net_),
            .in2(N__25317),
            .in3(N__32817),
            .lcout(n2429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_3_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_3_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_3_17_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1587_3_lut_LC_3_17_5 (
            .in0(N__25262),
            .in1(_gnd_net_),
            .in2(N__32828),
            .in3(N__25245),
            .lcout(n2427),
            .ltout(n2427_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_111_LC_3_17_6.C_ON=1'b0;
    defparam i1_4_lut_adj_111_LC_3_17_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_111_LC_3_17_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_111_LC_3_17_6 (
            .in0(N__23095),
            .in1(N__23368),
            .in2(N__23079),
            .in3(N__23075),
            .lcout(n14612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_129_LC_3_17_7.C_ON=1'b0;
    defparam i1_4_lut_adj_129_LC_3_17_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_129_LC_3_17_7.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_129_LC_3_17_7 (
            .in0(N__23446),
            .in1(N__23833),
            .in2(N__24106),
            .in3(N__23433),
            .lcout(n13790),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_123_LC_3_18_0.C_ON=1'b0;
    defparam i1_4_lut_adj_123_LC_3_18_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_123_LC_3_18_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_123_LC_3_18_0 (
            .in0(N__23314),
            .in1(N__23524),
            .in2(N__23427),
            .in3(N__23382),
            .lcout(),
            .ltout(n14622_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13070_4_lut_LC_3_18_1.C_ON=1'b0;
    defparam i13070_4_lut_LC_3_18_1.SEQ_MODE=4'b0000;
    defparam i13070_4_lut_LC_3_18_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13070_4_lut_LC_3_18_1 (
            .in0(N__23507),
            .in1(N__25514),
            .in2(N__23418),
            .in3(N__23415),
            .lcout(n2445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_3_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_3_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_3_18_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1580_3_lut_LC_3_18_2 (
            .in0(_gnd_net_),
            .in1(N__25404),
            .in2(N__28755),
            .in3(N__32798),
            .lcout(n2420),
            .ltout(n2420_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_113_LC_3_18_3.C_ON=1'b0;
    defparam i1_3_lut_adj_113_LC_3_18_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_113_LC_3_18_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_113_LC_3_18_3 (
            .in0(_gnd_net_),
            .in1(N__23341),
            .in2(N__23391),
            .in3(N__23388),
            .lcout(n14616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1586_3_lut_LC_3_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1586_3_lut_LC_3_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1586_3_lut_LC_3_18_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1586_3_lut_LC_3_18_4 (
            .in0(_gnd_net_),
            .in1(N__25236),
            .in2(N__25485),
            .in3(N__32793),
            .lcout(n2426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_3_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_3_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_3_18_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1581_3_lut_LC_3_18_5 (
            .in0(_gnd_net_),
            .in1(N__30056),
            .in2(N__32822),
            .in3(N__25413),
            .lcout(n2421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1583_3_lut_LC_3_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1583_3_lut_LC_3_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1583_3_lut_LC_3_18_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1583_3_lut_LC_3_18_6 (
            .in0(_gnd_net_),
            .in1(N__25434),
            .in2(N__29817),
            .in3(N__32794),
            .lcout(n2423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_3_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_3_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_3_18_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1573_3_lut_LC_3_18_7 (
            .in0(N__25533),
            .in1(_gnd_net_),
            .in2(N__32823),
            .in3(N__25503),
            .lcout(n2413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_3_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_3_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_3_19_0.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i1585_3_lut_LC_3_19_0 (
            .in0(N__32805),
            .in1(_gnd_net_),
            .in2(N__25227),
            .in3(N__25460),
            .lcout(n2425),
            .ltout(n2425_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_112_LC_3_19_1.C_ON=1'b0;
    defparam i1_4_lut_adj_112_LC_3_19_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_112_LC_3_19_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_112_LC_3_19_1 (
            .in0(N__23581),
            .in1(N__23623),
            .in2(N__23607),
            .in3(N__23704),
            .lcout(n14632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_3_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_3_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_3_19_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1579_3_lut_LC_3_19_2 (
            .in0(_gnd_net_),
            .in1(N__25619),
            .in2(N__32824),
            .in3(N__25395),
            .lcout(n2419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_3_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_3_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_3_19_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1575_3_lut_LC_3_19_3 (
            .in0(_gnd_net_),
            .in1(N__32806),
            .in2(N__32511),
            .in3(N__25353),
            .lcout(n2415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_110_LC_3_19_4.C_ON=1'b0;
    defparam i1_4_lut_adj_110_LC_3_19_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_110_LC_3_19_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_110_LC_3_19_4 (
            .in0(N__32500),
            .in1(N__25636),
            .in2(N__30251),
            .in3(N__23730),
            .lcout(),
            .ltout(n14456_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13043_4_lut_LC_3_19_5.C_ON=1'b0;
    defparam i13043_4_lut_LC_3_19_5.SEQ_MODE=4'b0000;
    defparam i13043_4_lut_LC_3_19_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13043_4_lut_LC_3_19_5 (
            .in0(N__28162),
            .in1(N__25501),
            .in2(N__23544),
            .in3(N__28389),
            .lcout(n2346),
            .ltout(n2346_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_3_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_3_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_3_19_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1577_3_lut_LC_3_19_6 (
            .in0(_gnd_net_),
            .in1(N__25637),
            .in2(N__23541),
            .in3(N__25374),
            .lcout(n2417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_3_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_3_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_3_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1574_3_lut_LC_3_19_7 (
            .in0(_gnd_net_),
            .in1(N__25542),
            .in2(N__28167),
            .in3(N__32807),
            .lcout(n2414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_130_LC_3_20_0.C_ON=1'b0;
    defparam i1_4_lut_adj_130_LC_3_20_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_130_LC_3_20_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_130_LC_3_20_0 (
            .in0(N__24024),
            .in1(N__23755),
            .in2(N__23484),
            .in3(N__23472),
            .lcout(n14324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_3_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_3_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_3_20_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1521_3_lut_LC_3_20_1 (
            .in0(_gnd_net_),
            .in1(N__28338),
            .in2(N__28236),
            .in3(N__32664),
            .lcout(n2329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_3_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_3_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_3_20_2.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i1520_3_lut_LC_3_20_2 (
            .in0(N__28221),
            .in1(N__30003),
            .in2(N__32682),
            .in3(_gnd_net_),
            .lcout(n2328),
            .ltout(n2328_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_107_LC_3_20_3.C_ON=1'b0;
    defparam i1_4_lut_adj_107_LC_3_20_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_107_LC_3_20_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_107_LC_3_20_3 (
            .in0(N__28744),
            .in1(N__29701),
            .in2(N__23739),
            .in3(N__29815),
            .lcout(),
            .ltout(n14442_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_108_LC_3_20_4.C_ON=1'b0;
    defparam i1_4_lut_adj_108_LC_3_20_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_108_LC_3_20_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_108_LC_3_20_4 (
            .in0(N__25585),
            .in1(N__25615),
            .in2(N__23736),
            .in3(N__25440),
            .lcout(),
            .ltout(n14448_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_109_LC_3_20_5.C_ON=1'b0;
    defparam i1_4_lut_adj_109_LC_3_20_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_109_LC_3_20_5.LUT_INIT=16'b1111100011110000;
    LogicCell40 i1_4_lut_adj_109_LC_3_20_5 (
            .in0(N__25297),
            .in1(N__29872),
            .in2(N__23733),
            .in3(N__28683),
            .lcout(n14450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1721_3_lut_LC_3_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1721_3_lut_LC_3_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1721_3_lut_LC_3_21_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1721_3_lut_LC_3_21_0 (
            .in0(_gnd_net_),
            .in1(N__23654),
            .in2(N__23724),
            .in3(N__33119),
            .lcout(n2625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_3_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_3_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_3_21_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1649_3_lut_LC_3_21_1 (
            .in0(_gnd_net_),
            .in1(N__23712),
            .in2(N__32998),
            .in3(N__23688),
            .lcout(n2521),
            .ltout(n2521_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_125_LC_3_21_2.C_ON=1'b0;
    defparam i1_4_lut_adj_125_LC_3_21_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_125_LC_3_21_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_125_LC_3_21_2 (
            .in0(N__23887),
            .in1(N__23653),
            .in2(N__23640),
            .in3(N__25654),
            .lcout(n14312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_131_LC_3_21_3.C_ON=1'b0;
    defparam i1_4_lut_adj_131_LC_3_21_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_131_LC_3_21_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_131_LC_3_21_3 (
            .in0(N__24280),
            .in1(N__24130),
            .in2(N__23988),
            .in3(N__23975),
            .lcout(),
            .ltout(n14330_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13099_4_lut_LC_3_21_4.C_ON=1'b0;
    defparam i13099_4_lut_LC_3_21_4.SEQ_MODE=4'b0000;
    defparam i13099_4_lut_LC_3_21_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13099_4_lut_LC_3_21_4 (
            .in0(N__23964),
            .in1(N__23929),
            .in2(N__23916),
            .in3(N__23913),
            .lcout(n2544),
            .ltout(n2544_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1718_rep_16_3_lut_LC_3_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1718_rep_16_3_lut_LC_3_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1718_rep_16_3_lut_LC_3_21_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1718_rep_16_3_lut_LC_3_21_5 (
            .in0(_gnd_net_),
            .in1(N__23888),
            .in2(N__23874),
            .in3(N__23871),
            .lcout(n2622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1719_3_lut_LC_3_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1719_3_lut_LC_3_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1719_3_lut_LC_3_21_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1719_3_lut_LC_3_21_6 (
            .in0(_gnd_net_),
            .in1(N__25655),
            .in2(N__23862),
            .in3(N__33120),
            .lcout(n2623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_3_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_3_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_3_22_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1725_3_lut_LC_3_22_0 (
            .in0(_gnd_net_),
            .in1(N__23849),
            .in2(N__23817),
            .in3(N__33114),
            .lcout(n2629),
            .ltout(n2629_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_140_LC_3_22_1.C_ON=1'b0;
    defparam i1_4_lut_adj_140_LC_3_22_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_140_LC_3_22_1.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_140_LC_3_22_1 (
            .in0(N__26530),
            .in1(N__28482),
            .in2(N__23799),
            .in3(N__23796),
            .lcout(n14658),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_3_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_3_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_3_22_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1729_3_lut_LC_3_22_2 (
            .in0(N__23790),
            .in1(N__28669),
            .in2(_gnd_net_),
            .in3(N__33110),
            .lcout(n2633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_3_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_3_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_3_22_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1782_3_lut_LC_3_22_3 (
            .in0(_gnd_net_),
            .in1(N__26177),
            .in2(N__26157),
            .in3(N__33343),
            .lcout(n2718),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_3_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_3_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_3_22_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1712_3_lut_LC_3_22_5 (
            .in0(_gnd_net_),
            .in1(N__23775),
            .in2(N__33156),
            .in3(N__23765),
            .lcout(n2616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_3_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_3_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_3_22_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1710_3_lut_LC_3_22_6 (
            .in0(_gnd_net_),
            .in1(N__24153),
            .in2(N__24144),
            .in3(N__33118),
            .lcout(n2614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_3_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_3_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_3_22_7.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1726_3_lut_LC_3_22_7 (
            .in0(N__24114),
            .in1(N__24081),
            .in2(N__33155),
            .in3(_gnd_net_),
            .lcout(n2630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_3_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_3_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_3_23_0.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1791_3_lut_LC_3_23_0 (
            .in0(N__25940),
            .in1(_gnd_net_),
            .in2(N__33328),
            .in3(N__25920),
            .lcout(n2727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_3_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_3_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_3_23_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1796_3_lut_LC_3_23_1 (
            .in0(_gnd_net_),
            .in1(N__25566),
            .in2(N__28535),
            .in3(N__33273),
            .lcout(n2732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_3_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_3_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_3_23_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1780_3_lut_LC_3_23_2 (
            .in0(N__26085),
            .in1(_gnd_net_),
            .in2(N__33329),
            .in3(N__26099),
            .lcout(n2716),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_3_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_3_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_3_23_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1713_3_lut_LC_3_23_3 (
            .in0(_gnd_net_),
            .in1(N__24036),
            .in2(N__33165),
            .in3(N__24023),
            .lcout(n2617),
            .ltout(n2617_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_141_LC_3_23_4.C_ON=1'b0;
    defparam i1_4_lut_adj_141_LC_3_23_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_141_LC_3_23_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_141_LC_3_23_4 (
            .in0(N__26075),
            .in1(N__23997),
            .in2(N__23991),
            .in3(N__26125),
            .lcout(n14664),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1788_3_lut_LC_3_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1788_3_lut_LC_3_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1788_3_lut_LC_3_23_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1788_3_lut_LC_3_23_5 (
            .in0(N__25833),
            .in1(N__25812),
            .in2(_gnd_net_),
            .in3(N__33278),
            .lcout(n2724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_3_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_3_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_3_23_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1789_3_lut_LC_3_23_7 (
            .in0(_gnd_net_),
            .in1(N__25842),
            .in2(N__25866),
            .in3(N__33274),
            .lcout(n2725),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_3_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_3_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_3_24_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1781_3_lut_LC_3_24_0 (
            .in0(_gnd_net_),
            .in1(N__26109),
            .in2(N__26145),
            .in3(N__33301),
            .lcout(n2717),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_3_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_3_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_3_24_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1792_3_lut_LC_3_24_1 (
            .in0(N__25971),
            .in1(_gnd_net_),
            .in2(N__33339),
            .in3(N__25953),
            .lcout(n2728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_3_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_3_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_3_24_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1709_3_lut_LC_3_24_2 (
            .in0(_gnd_net_),
            .in1(N__24291),
            .in2(N__24264),
            .in3(N__33148),
            .lcout(n2613),
            .ltout(n2613_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_142_LC_3_24_3.C_ON=1'b0;
    defparam i1_4_lut_adj_142_LC_3_24_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_142_LC_3_24_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_142_LC_3_24_3 (
            .in0(N__26032),
            .in1(N__25997),
            .in2(N__24249),
            .in3(N__24246),
            .lcout(),
            .ltout(n14670_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13130_4_lut_LC_3_24_4.C_ON=1'b0;
    defparam i13130_4_lut_LC_3_24_4.SEQ_MODE=4'b0000;
    defparam i13130_4_lut_LC_3_24_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13130_4_lut_LC_3_24_4 (
            .in0(N__26408),
            .in1(N__26368),
            .in2(N__24240),
            .in3(N__26321),
            .lcout(n2643),
            .ltout(n2643_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_3_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_3_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_3_24_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1777_3_lut_LC_3_24_5 (
            .in0(N__25980),
            .in1(_gnd_net_),
            .in2(N__24237),
            .in3(N__25998),
            .lcout(n2713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1720_rep_14_3_lut_LC_3_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1720_rep_14_3_lut_LC_3_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1720_rep_14_3_lut_LC_3_24_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1720_rep_14_3_lut_LC_3_24_6 (
            .in0(_gnd_net_),
            .in1(N__24213),
            .in2(N__25785),
            .in3(N__33296),
            .lcout(),
            .ltout(n14889_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1787_3_lut_4_lut_LC_3_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1787_3_lut_4_lut_LC_3_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1787_3_lut_4_lut_LC_3_24_7.LUT_INIT=16'b1111100001110000;
    LogicCell40 encoder0_position_31__I_0_i1787_3_lut_4_lut_LC_3_24_7 (
            .in0(N__33297),
            .in1(N__33166),
            .in2(N__24192),
            .in3(N__24189),
            .lcout(n2723),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_3_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_3_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_3_25_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1779_3_lut_LC_3_25_0 (
            .in0(N__26055),
            .in1(_gnd_net_),
            .in2(N__33341),
            .in3(N__26076),
            .lcout(n2715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1790_3_lut_LC_3_25_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1790_3_lut_LC_3_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1790_3_lut_LC_3_25_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1790_3_lut_LC_3_25_1 (
            .in0(_gnd_net_),
            .in1(N__25908),
            .in2(N__25884),
            .in3(N__33302),
            .lcout(n2726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1785_3_lut_LC_3_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1785_3_lut_LC_3_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1785_3_lut_LC_3_25_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1785_3_lut_LC_3_25_2 (
            .in0(N__25713),
            .in1(_gnd_net_),
            .in2(N__33340),
            .in3(N__25734),
            .lcout(n2721),
            .ltout(n2721_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_146_LC_3_25_3.C_ON=1'b0;
    defparam i1_4_lut_adj_146_LC_3_25_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_146_LC_3_25_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_146_LC_3_25_3 (
            .in0(N__24367),
            .in1(N__24328),
            .in2(N__24501),
            .in3(N__26646),
            .lcout(),
            .ltout(n14140_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_147_LC_3_25_4.C_ON=1'b0;
    defparam i1_4_lut_adj_147_LC_3_25_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_147_LC_3_25_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_147_LC_3_25_4 (
            .in0(N__24493),
            .in1(N__24469),
            .in2(N__24450),
            .in3(N__24447),
            .lcout(),
            .ltout(n14146_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_149_LC_3_25_5.C_ON=1'b0;
    defparam i1_4_lut_adj_149_LC_3_25_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_149_LC_3_25_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_149_LC_3_25_5 (
            .in0(N__24427),
            .in1(N__24400),
            .in2(N__24384),
            .in3(N__26445),
            .lcout(n14152),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1786_3_lut_LC_3_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1786_3_lut_LC_3_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1786_3_lut_LC_3_25_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1786_3_lut_LC_3_25_7 (
            .in0(_gnd_net_),
            .in1(N__25746),
            .in2(N__25770),
            .in3(N__33303),
            .lcout(n2722),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_3_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_3_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_3_26_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1851_3_lut_LC_3_26_0 (
            .in0(_gnd_net_),
            .in1(N__26736),
            .in2(N__33515),
            .in3(N__24351),
            .lcout(n2819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_3_26_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_3_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_3_26_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1859_3_lut_LC_3_26_2 (
            .in0(_gnd_net_),
            .in1(N__24342),
            .in2(N__33512),
            .in3(N__24333),
            .lcout(n2827),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_3_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_3_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_3_26_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1776_3_lut_LC_3_26_3 (
            .in0(N__26439),
            .in1(N__26424),
            .in2(_gnd_net_),
            .in3(N__33334),
            .lcout(n2712),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_3_26_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_3_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_3_26_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1856_3_lut_LC_3_26_4 (
            .in0(N__24651),
            .in1(_gnd_net_),
            .in2(N__33513),
            .in3(N__24624),
            .lcout(n2824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_3_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_3_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_3_26_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1774_3_lut_LC_3_26_5 (
            .in0(_gnd_net_),
            .in1(N__26375),
            .in2(N__26346),
            .in3(N__33335),
            .lcout(n2710),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12515_3_lut_LC_3_26_6.C_ON=1'b0;
    defparam i12515_3_lut_LC_3_26_6.SEQ_MODE=4'b0000;
    defparam i12515_3_lut_LC_3_26_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12515_3_lut_LC_3_26_6 (
            .in0(N__24612),
            .in1(_gnd_net_),
            .in2(N__33514),
            .in3(N__24600),
            .lcout(n2820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1857_3_lut_LC_3_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1857_3_lut_LC_3_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1857_3_lut_LC_3_26_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1857_3_lut_LC_3_26_7 (
            .in0(_gnd_net_),
            .in1(N__26717),
            .in2(N__24591),
            .in3(N__33470),
            .lcout(n2825),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_3_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_3_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_3_27_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1921_3_lut_LC_3_27_0 (
            .in0(N__24536),
            .in1(_gnd_net_),
            .in2(N__24579),
            .in3(N__33646),
            .lcout(n2921),
            .ltout(n2921_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_43_LC_3_27_1.C_ON=1'b0;
    defparam i1_4_lut_adj_43_LC_3_27_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_43_LC_3_27_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_43_LC_3_27_1 (
            .in0(N__27544),
            .in1(N__27673),
            .in2(N__24567),
            .in3(N__24784),
            .lcout(n14346),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_3_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_3_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_3_27_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1920_3_lut_LC_3_27_2 (
            .in0(_gnd_net_),
            .in1(N__24515),
            .in2(N__24564),
            .in3(N__33645),
            .lcout(n2920),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1855_3_lut_LC_3_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1855_3_lut_LC_3_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1855_3_lut_LC_3_27_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1855_3_lut_LC_3_27_3 (
            .in0(N__26697),
            .in1(_gnd_net_),
            .in2(N__24552),
            .in3(N__33463),
            .lcout(n2823),
            .ltout(n2823_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_28_LC_3_27_4.C_ON=1'b0;
    defparam i1_4_lut_adj_28_LC_3_27_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_28_LC_3_27_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_28_LC_3_27_4 (
            .in0(N__24535),
            .in1(N__25024),
            .in2(N__24522),
            .in3(N__24514),
            .lcout(n14690),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_3_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_3_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_3_27_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1841_3_lut_LC_3_27_5 (
            .in0(N__24921),
            .in1(_gnd_net_),
            .in2(N__24915),
            .in3(N__33464),
            .lcout(n2809),
            .ltout(n2809_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12625_4_lut_LC_3_27_6.C_ON=1'b0;
    defparam i12625_4_lut_LC_3_27_6.SEQ_MODE=4'b0000;
    defparam i12625_4_lut_LC_3_27_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12625_4_lut_LC_3_27_6 (
            .in0(N__24871),
            .in1(N__24842),
            .in2(N__24831),
            .in3(N__24828),
            .lcout(n2841),
            .ltout(n2841_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_3_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_3_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_3_27_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1922_3_lut_LC_3_27_7 (
            .in0(N__24818),
            .in1(_gnd_net_),
            .in2(N__24804),
            .in3(N__24801),
            .lcout(n2922),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_3_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_3_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_3_28_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1987_3_lut_LC_3_28_0 (
            .in0(_gnd_net_),
            .in1(N__24788),
            .in2(N__24768),
            .in3(N__33845),
            .lcout(n3019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_3_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_3_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_3_28_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1930_3_lut_LC_3_28_1 (
            .in0(_gnd_net_),
            .in1(N__24756),
            .in2(N__24744),
            .in3(N__33655),
            .lcout(n2930),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_3_28_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_3_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_3_28_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1911_3_lut_LC_3_28_2 (
            .in0(_gnd_net_),
            .in1(N__24714),
            .in2(N__33698),
            .in3(N__24705),
            .lcout(n2911),
            .ltout(n2911_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_48_LC_3_28_3.C_ON=1'b0;
    defparam i1_4_lut_adj_48_LC_3_28_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_48_LC_3_28_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_48_LC_3_28_3 (
            .in0(N__28024),
            .in1(N__27709),
            .in2(N__24687),
            .in3(N__26961),
            .lcout(n14372),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_3_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_3_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_3_28_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1928_3_lut_LC_3_28_4 (
            .in0(_gnd_net_),
            .in1(N__24684),
            .in2(N__33697),
            .in3(N__24663),
            .lcout(n2928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_3_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_3_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_3_28_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1925_3_lut_LC_3_28_5 (
            .in0(_gnd_net_),
            .in1(N__25044),
            .in2(N__25032),
            .in3(N__33651),
            .lcout(n2925),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_3_28_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_3_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_3_28_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i1914_3_lut_LC_3_28_6 (
            .in0(N__33656),
            .in1(_gnd_net_),
            .in2(N__25008),
            .in3(N__24996),
            .lcout(n2914),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_3_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_3_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_3_28_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1912_3_lut_LC_3_28_7 (
            .in0(_gnd_net_),
            .in1(N__24972),
            .in2(N__24954),
            .in3(N__33657),
            .lcout(n2912),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_3_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_3_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_3_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_2_lut_LC_3_29_0 (
            .in0(_gnd_net_),
            .in1(N__42225),
            .in2(_gnd_net_),
            .in3(N__24939),
            .lcout(n3101),
            .ltout(),
            .carryin(bfn_3_29_0_),
            .carryout(n12850),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_3_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_3_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_3_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_3_lut_LC_3_29_1 (
            .in0(_gnd_net_),
            .in1(N__53714),
            .in2(N__29118),
            .in3(N__24936),
            .lcout(n3100),
            .ltout(),
            .carryin(n12850),
            .carryout(n12851),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_3_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_3_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_3_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_4_lut_LC_3_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29097),
            .in3(N__24933),
            .lcout(n3099),
            .ltout(),
            .carryin(n12851),
            .carryout(n12852),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_3_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_3_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_3_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_5_lut_LC_3_29_3 (
            .in0(_gnd_net_),
            .in1(N__53715),
            .in2(N__29400),
            .in3(N__24930),
            .lcout(n3098),
            .ltout(),
            .carryin(n12852),
            .carryout(n12853),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_3_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_3_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_3_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_6_lut_LC_3_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29052),
            .in3(N__24927),
            .lcout(n3097),
            .ltout(),
            .carryin(n12853),
            .carryout(n12854),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_3_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_3_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_3_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_7_lut_LC_3_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29037),
            .in3(N__24924),
            .lcout(n3096),
            .ltout(),
            .carryin(n12854),
            .carryout(n12855),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_3_29_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_3_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_3_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_8_lut_LC_3_29_6 (
            .in0(_gnd_net_),
            .in1(N__53717),
            .in2(N__29235),
            .in3(N__25071),
            .lcout(n3095),
            .ltout(),
            .carryin(n12855),
            .carryout(n12856),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_3_29_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_3_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_3_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_9_lut_LC_3_29_7 (
            .in0(_gnd_net_),
            .in1(N__53716),
            .in2(N__28877),
            .in3(N__25068),
            .lcout(n3094),
            .ltout(),
            .carryin(n12856),
            .carryout(n12857),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_3_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_3_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_3_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_10_lut_LC_3_30_0 (
            .in0(_gnd_net_),
            .in1(N__31385),
            .in2(N__54456),
            .in3(N__25065),
            .lcout(n3093),
            .ltout(),
            .carryin(bfn_3_30_0_),
            .carryout(n12858),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_3_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_3_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_3_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_11_lut_LC_3_30_1 (
            .in0(_gnd_net_),
            .in1(N__54345),
            .in2(N__29475),
            .in3(N__25062),
            .lcout(n3092),
            .ltout(),
            .carryin(n12858),
            .carryout(n12859),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_3_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_3_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_3_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_12_lut_LC_3_30_2 (
            .in0(_gnd_net_),
            .in1(N__54352),
            .in2(N__37269),
            .in3(N__25059),
            .lcout(n3091),
            .ltout(),
            .carryin(n12859),
            .carryout(n12860),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_3_30_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_3_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_3_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_13_lut_LC_3_30_3 (
            .in0(_gnd_net_),
            .in1(N__54346),
            .in2(N__31169),
            .in3(N__25056),
            .lcout(n3090),
            .ltout(),
            .carryin(n12860),
            .carryout(n12861),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_3_30_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_3_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_3_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_14_lut_LC_3_30_4 (
            .in0(_gnd_net_),
            .in1(N__29264),
            .in2(N__54457),
            .in3(N__25053),
            .lcout(n3089),
            .ltout(),
            .carryin(n12861),
            .carryout(n12862),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_3_30_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_3_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_3_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_15_lut_LC_3_30_5 (
            .in0(_gnd_net_),
            .in1(N__54350),
            .in2(N__31496),
            .in3(N__25050),
            .lcout(n3088),
            .ltout(),
            .carryin(n12862),
            .carryout(n12863),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_3_30_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_3_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_3_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_16_lut_LC_3_30_6 (
            .in0(_gnd_net_),
            .in1(N__54353),
            .in2(N__27405),
            .in3(N__25047),
            .lcout(n3087),
            .ltout(),
            .carryin(n12863),
            .carryout(n12864),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_3_30_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_3_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_3_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_17_lut_LC_3_30_7 (
            .in0(_gnd_net_),
            .in1(N__54351),
            .in2(N__27579),
            .in3(N__25098),
            .lcout(n3086),
            .ltout(),
            .carryin(n12864),
            .carryout(n12865),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_3_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_3_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_3_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_18_lut_LC_3_31_0 (
            .in0(_gnd_net_),
            .in1(N__29540),
            .in2(N__54264),
            .in3(N__25095),
            .lcout(n3085),
            .ltout(),
            .carryin(bfn_3_31_0_),
            .carryout(n12866),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_3_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_3_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_3_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_19_lut_LC_3_31_1 (
            .in0(_gnd_net_),
            .in1(N__29504),
            .in2(N__54268),
            .in3(N__25092),
            .lcout(n3084),
            .ltout(),
            .carryin(n12866),
            .carryout(n12867),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_3_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_3_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_3_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_20_lut_LC_3_31_2 (
            .in0(_gnd_net_),
            .in1(N__27641),
            .in2(N__54265),
            .in3(N__25089),
            .lcout(n3083),
            .ltout(),
            .carryin(n12867),
            .carryout(n12868),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_3_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_3_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_3_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_21_lut_LC_3_31_3 (
            .in0(_gnd_net_),
            .in1(N__29313),
            .in2(N__54269),
            .in3(N__25086),
            .lcout(n3082),
            .ltout(),
            .carryin(n12868),
            .carryout(n12869),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_3_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_3_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_3_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_22_lut_LC_3_31_4 (
            .in0(_gnd_net_),
            .in1(N__29171),
            .in2(N__54266),
            .in3(N__25083),
            .lcout(n3081),
            .ltout(),
            .carryin(n12869),
            .carryout(n12870),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_3_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_3_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_3_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_23_lut_LC_3_31_5 (
            .in0(_gnd_net_),
            .in1(N__34331),
            .in2(N__54270),
            .in3(N__25080),
            .lcout(n3080),
            .ltout(),
            .carryin(n12870),
            .carryout(n12871),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_3_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_3_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_3_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_24_lut_LC_3_31_6 (
            .in0(_gnd_net_),
            .in1(N__29570),
            .in2(N__54267),
            .in3(N__25077),
            .lcout(n3079),
            .ltout(),
            .carryin(n12871),
            .carryout(n12872),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_3_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_3_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_3_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_25_lut_LC_3_31_7 (
            .in0(_gnd_net_),
            .in1(N__29207),
            .in2(N__54271),
            .in3(N__25074),
            .lcout(n3078),
            .ltout(),
            .carryin(n12872),
            .carryout(n12873),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_3_32_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_3_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_3_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_26_lut_LC_3_32_0 (
            .in0(_gnd_net_),
            .in1(N__29753),
            .in2(N__54281),
            .in3(N__25200),
            .lcout(n3077),
            .ltout(),
            .carryin(bfn_3_32_0_),
            .carryout(n12874),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_3_32_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_3_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_3_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_27_lut_LC_3_32_1 (
            .in0(_gnd_net_),
            .in1(N__29666),
            .in2(N__54276),
            .in3(N__25197),
            .lcout(n3076),
            .ltout(),
            .carryin(n12874),
            .carryout(n12875),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_3_32_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_3_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_3_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_28_lut_LC_3_32_2 (
            .in0(_gnd_net_),
            .in1(N__29623),
            .in2(N__54282),
            .in3(N__25194),
            .lcout(n3075),
            .ltout(),
            .carryin(n12875),
            .carryout(n12876),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_3_32_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_3_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_3_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_29_lut_LC_3_32_3 (
            .in0(_gnd_net_),
            .in1(N__29649),
            .in2(N__54277),
            .in3(N__25191),
            .lcout(n3074),
            .ltout(),
            .carryin(n12876),
            .carryout(n12877),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_3_32_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_3_32_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_3_32_4.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_2039_30_lut_LC_3_32_4 (
            .in0(N__54078),
            .in1(N__29597),
            .in2(N__32336),
            .in3(N__25188),
            .lcout(n3105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i9_4_lut_LC_3_32_5 .C_ON=1'b0;
    defparam \debounce.i9_4_lut_LC_3_32_5 .SEQ_MODE=4'b0000;
    defparam \debounce.i9_4_lut_LC_3_32_5 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \debounce.i9_4_lut_LC_3_32_5  (
            .in0(N__25185),
            .in1(N__25167),
            .in2(N__25161),
            .in3(N__25140),
            .lcout(n14125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i2_LC_3_32_6 .C_ON=1'b0;
    defparam \debounce.reg_B_i2_LC_3_32_6 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i2_LC_3_32_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \debounce.reg_B_i2_LC_3_32_6  (
            .in0(N__27996),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(reg_B_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55788),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_4_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_4_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_4_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_2_lut_LC_4_17_0 (
            .in0(_gnd_net_),
            .in1(N__30578),
            .in2(_gnd_net_),
            .in3(N__25125),
            .lcout(n2401),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(n12682),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_4_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_4_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_4_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_3_lut_LC_4_17_1 (
            .in0(_gnd_net_),
            .in1(N__28454),
            .in2(N__54505),
            .in3(N__25113),
            .lcout(n2400),
            .ltout(),
            .carryin(n12682),
            .carryout(n12683),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_4_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_4_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_4_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_4_lut_LC_4_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30099),
            .in3(N__25335),
            .lcout(n2399),
            .ltout(),
            .carryin(n12683),
            .carryout(n12684),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_4_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_4_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_4_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_5_lut_LC_4_17_3 (
            .in0(_gnd_net_),
            .in1(N__28712),
            .in2(N__54506),
            .in3(N__25320),
            .lcout(n2398),
            .ltout(),
            .carryin(n12684),
            .carryout(n12685),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_4_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_4_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_4_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_6_lut_LC_4_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29874),
            .in3(N__25308),
            .lcout(n2397),
            .ltout(),
            .carryin(n12685),
            .carryout(n12686),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_4_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_4_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_4_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_7_lut_LC_4_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25305),
            .in3(N__25266),
            .lcout(n2396),
            .ltout(),
            .carryin(n12686),
            .carryout(n12687),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_4_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_4_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_4_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_8_lut_LC_4_17_6 (
            .in0(_gnd_net_),
            .in1(N__54413),
            .in2(N__25263),
            .in3(N__25239),
            .lcout(n2395),
            .ltout(),
            .carryin(n12687),
            .carryout(n12688),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_4_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_4_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_4_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_9_lut_LC_4_17_7 (
            .in0(_gnd_net_),
            .in1(N__54414),
            .in2(N__25484),
            .in3(N__25230),
            .lcout(n2394),
            .ltout(),
            .carryin(n12688),
            .carryout(n12689),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_4_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_4_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_4_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_10_lut_LC_4_18_0 (
            .in0(_gnd_net_),
            .in1(N__54519),
            .in2(N__25461),
            .in3(N__25218),
            .lcout(n2393),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(n12690),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_4_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_4_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_4_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_11_lut_LC_4_18_1 (
            .in0(_gnd_net_),
            .in1(N__54526),
            .in2(N__28139),
            .in3(N__25203),
            .lcout(n2392),
            .ltout(),
            .carryin(n12690),
            .carryout(n12691),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_4_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_4_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_4_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_12_lut_LC_4_18_2 (
            .in0(_gnd_net_),
            .in1(N__54520),
            .in2(N__29816),
            .in3(N__25428),
            .lcout(n2391),
            .ltout(),
            .carryin(n12691),
            .carryout(n12692),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_4_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_4_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_4_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_13_lut_LC_4_18_3 (
            .in0(_gnd_net_),
            .in1(N__54527),
            .in2(N__29702),
            .in3(N__25416),
            .lcout(n2390),
            .ltout(),
            .carryin(n12692),
            .carryout(n12693),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_4_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_4_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_4_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_14_lut_LC_4_18_4 (
            .in0(_gnd_net_),
            .in1(N__54521),
            .in2(N__30057),
            .in3(N__25407),
            .lcout(n2389),
            .ltout(),
            .carryin(n12693),
            .carryout(n12694),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_4_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_4_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_4_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_15_lut_LC_4_18_5 (
            .in0(_gnd_net_),
            .in1(N__54528),
            .in2(N__28754),
            .in3(N__25398),
            .lcout(n2388),
            .ltout(),
            .carryin(n12694),
            .carryout(n12695),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_4_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_4_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_4_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_16_lut_LC_4_18_6 (
            .in0(_gnd_net_),
            .in1(N__54522),
            .in2(N__25623),
            .in3(N__25389),
            .lcout(n2387),
            .ltout(),
            .carryin(n12695),
            .carryout(n12696),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_4_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_4_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_4_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_17_lut_LC_4_18_7 (
            .in0(_gnd_net_),
            .in1(N__25592),
            .in2(N__54543),
            .in3(N__25377),
            .lcout(n2386),
            .ltout(),
            .carryin(n12696),
            .carryout(n12697),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_4_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_4_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_4_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_18_lut_LC_4_19_0 (
            .in0(_gnd_net_),
            .in1(N__54096),
            .in2(N__25641),
            .in3(N__25368),
            .lcout(n2385),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(n12698),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_4_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_4_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_4_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_19_lut_LC_4_19_1 (
            .in0(_gnd_net_),
            .in1(N__53916),
            .in2(N__30252),
            .in3(N__25356),
            .lcout(n2384),
            .ltout(),
            .carryin(n12698),
            .carryout(n12699),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_4_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_4_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_4_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_20_lut_LC_4_19_2 (
            .in0(_gnd_net_),
            .in1(N__54097),
            .in2(N__32507),
            .in3(N__25545),
            .lcout(n2383),
            .ltout(),
            .carryin(n12699),
            .carryout(n12700),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_4_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_4_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_4_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_21_lut_LC_4_19_3 (
            .in0(_gnd_net_),
            .in1(N__53917),
            .in2(N__28166),
            .in3(N__25536),
            .lcout(n2382),
            .ltout(),
            .carryin(n12700),
            .carryout(n12701),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_4_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_4_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_4_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_22_lut_LC_4_19_4 (
            .in0(_gnd_net_),
            .in1(N__25502),
            .in2(N__54184),
            .in3(N__25527),
            .lcout(n2381),
            .ltout(),
            .carryin(n12701),
            .carryout(n12702),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_4_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_4_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_4_19_5.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1570_23_lut_LC_4_19_5 (
            .in0(N__54098),
            .in1(N__28388),
            .in2(N__32846),
            .in3(N__25524),
            .lcout(n2412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_4_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_4_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_4_19_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1506_3_lut_LC_4_19_6 (
            .in0(_gnd_net_),
            .in1(N__28407),
            .in2(N__32685),
            .in3(N__29925),
            .lcout(n2314_adj_622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_4_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_4_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_4_19_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1518_3_lut_LC_4_19_7 (
            .in0(_gnd_net_),
            .in1(N__30451),
            .in2(N__28197),
            .in3(N__32676),
            .lcout(n2326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13040_1_lut_LC_4_20_0.C_ON=1'b0;
    defparam i13040_1_lut_LC_4_20_0.SEQ_MODE=4'b0000;
    defparam i13040_1_lut_LC_4_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i13040_1_lut_LC_4_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32808),
            .lcout(n15765),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1519_3_lut_LC_4_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1519_3_lut_LC_4_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1519_3_lut_LC_4_20_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1519_3_lut_LC_4_20_2 (
            .in0(_gnd_net_),
            .in1(N__30507),
            .in2(N__28209),
            .in3(N__32656),
            .lcout(n2327),
            .ltout(n2327_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_106_LC_4_20_3.C_ON=1'b0;
    defparam i1_4_lut_adj_106_LC_4_20_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_106_LC_4_20_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_106_LC_4_20_3 (
            .in0(N__30046),
            .in1(N__28132),
            .in2(N__25464),
            .in3(N__25456),
            .lcout(n14440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1652_3_lut_LC_4_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1652_3_lut_LC_4_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1652_3_lut_LC_4_20_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1652_3_lut_LC_4_20_4 (
            .in0(_gnd_net_),
            .in1(N__25701),
            .in2(N__25685),
            .in3(N__32966),
            .lcout(n2524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_4_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_4_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_4_20_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1510_3_lut_LC_4_20_5 (
            .in0(_gnd_net_),
            .in1(N__28266),
            .in2(N__32681),
            .in3(N__30153),
            .lcout(n2318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_4_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_4_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_4_20_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1512_3_lut_LC_4_20_6 (
            .in0(N__28284),
            .in1(_gnd_net_),
            .in2(N__30357),
            .in3(N__32660),
            .lcout(n2320),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_4_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_4_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_4_20_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1511_3_lut_LC_4_20_7 (
            .in0(N__28275),
            .in1(_gnd_net_),
            .in2(N__32680),
            .in3(N__30327),
            .lcout(n2319),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_4_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_4_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_4_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_2_lut_LC_4_21_0 (
            .in0(_gnd_net_),
            .in1(N__40117),
            .in2(_gnd_net_),
            .in3(N__25569),
            .lcout(n2701),
            .ltout(),
            .carryin(bfn_4_21_0_),
            .carryout(n12748),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_4_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_4_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_4_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_3_lut_LC_4_21_1 (
            .in0(_gnd_net_),
            .in1(N__54460),
            .in2(N__28534),
            .in3(N__25557),
            .lcout(n2700),
            .ltout(),
            .carryin(n12748),
            .carryout(n12749),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_4_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_4_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_4_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_4_lut_LC_4_21_2 (
            .in0(_gnd_net_),
            .in1(N__28503),
            .in2(_gnd_net_),
            .in3(N__25554),
            .lcout(n2699),
            .ltout(),
            .carryin(n12749),
            .carryout(n12750),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_4_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_4_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_4_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_5_lut_LC_4_21_3 (
            .in0(_gnd_net_),
            .in1(N__28551),
            .in2(N__54518),
            .in3(N__25551),
            .lcout(n2698),
            .ltout(),
            .carryin(n12750),
            .carryout(n12751),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_4_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_4_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_4_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_6_lut_LC_4_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26537),
            .in3(N__25548),
            .lcout(n2697),
            .ltout(),
            .carryin(n12751),
            .carryout(n12752),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_4_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_4_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_4_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_7_lut_LC_4_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25970),
            .in3(N__25944),
            .lcout(n2696),
            .ltout(),
            .carryin(n12752),
            .carryout(n12753),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_4_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_4_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_4_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_8_lut_LC_4_21_6 (
            .in0(_gnd_net_),
            .in1(N__54465),
            .in2(N__25941),
            .in3(N__25911),
            .lcout(n2695),
            .ltout(),
            .carryin(n12753),
            .carryout(n12754),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_4_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_4_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_4_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_9_lut_LC_4_21_7 (
            .in0(_gnd_net_),
            .in1(N__54461),
            .in2(N__25904),
            .in3(N__25869),
            .lcout(n2694),
            .ltout(),
            .carryin(n12754),
            .carryout(n12755),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_4_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_4_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_4_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_10_lut_LC_4_22_0 (
            .in0(_gnd_net_),
            .in1(N__25865),
            .in2(N__53187),
            .in3(N__25836),
            .lcout(n2693),
            .ltout(),
            .carryin(bfn_4_22_0_),
            .carryout(n12756),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_4_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_4_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_4_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_11_lut_LC_4_22_1 (
            .in0(_gnd_net_),
            .in1(N__25829),
            .in2(N__53191),
            .in3(N__25806),
            .lcout(n2692),
            .ltout(),
            .carryin(n12756),
            .carryout(n12757),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_4_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_4_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_4_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_12_lut_LC_4_22_2 (
            .in0(_gnd_net_),
            .in1(N__25803),
            .in2(N__53188),
            .in3(N__25773),
            .lcout(n2691),
            .ltout(),
            .carryin(n12757),
            .carryout(n12758),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_4_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_4_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_4_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_13_lut_LC_4_22_3 (
            .in0(_gnd_net_),
            .in1(N__25763),
            .in2(N__53192),
            .in3(N__25737),
            .lcout(n2690),
            .ltout(),
            .carryin(n12758),
            .carryout(n12759),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_4_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_4_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_4_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_14_lut_LC_4_22_4 (
            .in0(_gnd_net_),
            .in1(N__25730),
            .in2(N__53189),
            .in3(N__25704),
            .lcout(n2689),
            .ltout(),
            .carryin(n12759),
            .carryout(n12760),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_4_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_4_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_4_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_15_lut_LC_4_22_5 (
            .in0(_gnd_net_),
            .in1(N__26249),
            .in2(N__53193),
            .in3(N__26223),
            .lcout(n2688),
            .ltout(),
            .carryin(n12760),
            .carryout(n12761),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_4_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_4_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_4_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_16_lut_LC_4_22_6 (
            .in0(_gnd_net_),
            .in1(N__26220),
            .in2(N__53190),
            .in3(N__26184),
            .lcout(n2687),
            .ltout(),
            .carryin(n12761),
            .carryout(n12762),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_4_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_4_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_4_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_17_lut_LC_4_22_7 (
            .in0(_gnd_net_),
            .in1(N__26181),
            .in2(N__53194),
            .in3(N__26148),
            .lcout(n2686),
            .ltout(),
            .carryin(n12762),
            .carryout(n12763),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_4_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_4_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_4_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_18_lut_LC_4_23_0 (
            .in0(_gnd_net_),
            .in1(N__26138),
            .in2(N__54092),
            .in3(N__26103),
            .lcout(n2685),
            .ltout(),
            .carryin(bfn_4_23_0_),
            .carryout(n12764),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_4_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_4_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_4_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_19_lut_LC_4_23_1 (
            .in0(_gnd_net_),
            .in1(N__53818),
            .in2(N__26100),
            .in3(N__26079),
            .lcout(n2684),
            .ltout(),
            .carryin(n12764),
            .carryout(n12765),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_4_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_4_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_4_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_20_lut_LC_4_23_2 (
            .in0(_gnd_net_),
            .in1(N__26074),
            .in2(N__54093),
            .in3(N__26046),
            .lcout(n2683),
            .ltout(),
            .carryin(n12765),
            .carryout(n12766),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_4_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_4_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_4_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_21_lut_LC_4_23_3 (
            .in0(_gnd_net_),
            .in1(N__26039),
            .in2(N__54176),
            .in3(N__26001),
            .lcout(n2682),
            .ltout(),
            .carryin(n12766),
            .carryout(n12767),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_4_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_4_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_4_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_22_lut_LC_4_23_4 (
            .in0(_gnd_net_),
            .in1(N__25996),
            .in2(N__54094),
            .in3(N__25974),
            .lcout(n2681),
            .ltout(),
            .carryin(n12767),
            .carryout(n12768),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_4_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_4_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_4_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_23_lut_LC_4_23_5 (
            .in0(_gnd_net_),
            .in1(N__26435),
            .in2(N__54177),
            .in3(N__26415),
            .lcout(n2680),
            .ltout(),
            .carryin(n12768),
            .carryout(n12769),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_4_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_4_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_4_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_24_lut_LC_4_23_6 (
            .in0(_gnd_net_),
            .in1(N__26412),
            .in2(N__54095),
            .in3(N__26379),
            .lcout(n2679),
            .ltout(),
            .carryin(n12769),
            .carryout(n12770),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_4_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_4_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_4_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_25_lut_LC_4_23_7 (
            .in0(_gnd_net_),
            .in1(N__26376),
            .in2(N__54178),
            .in3(N__26331),
            .lcout(n2678),
            .ltout(),
            .carryin(n12770),
            .carryout(n12771),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_4_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_4_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_4_24_0.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1771_26_lut_LC_4_24_0 (
            .in0(N__53814),
            .in1(N__33362),
            .in2(N__26328),
            .in3(N__26301),
            .lcout(n2709),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13066_1_lut_LC_4_24_1.C_ON=1'b0;
    defparam i13066_1_lut_LC_4_24_1.SEQ_MODE=4'b0000;
    defparam i13066_1_lut_LC_4_24_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i13066_1_lut_LC_4_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32987),
            .lcout(n15791),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_4_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_4_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_4_24_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i13_3_lut_LC_4_24_2 (
            .in0(N__38697),
            .in1(N__46200),
            .in2(_gnd_net_),
            .in3(N__36609),
            .lcout(n307),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13127_1_lut_LC_4_24_3.C_ON=1'b0;
    defparam i13127_1_lut_LC_4_24_3.SEQ_MODE=4'b0000;
    defparam i13127_1_lut_LC_4_24_3.LUT_INIT=16'b0000111100001111;
    LogicCell40 i13127_1_lut_LC_4_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33345),
            .in3(_gnd_net_),
            .lcout(n15852),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_4_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_4_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_4_24_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1915_3_lut_LC_4_24_5 (
            .in0(_gnd_net_),
            .in1(N__26283),
            .in2(N__26265),
            .in3(N__33709),
            .lcout(n2915),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_4_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_4_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_4_24_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1784_3_lut_LC_4_24_6 (
            .in0(_gnd_net_),
            .in1(N__26250),
            .in2(N__26748),
            .in3(N__33321),
            .lcout(n2720),
            .ltout(n2720_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_143_LC_4_24_7.C_ON=1'b0;
    defparam i1_4_lut_adj_143_LC_4_24_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_143_LC_4_24_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_143_LC_4_24_7 (
            .in0(N__26713),
            .in1(N__26689),
            .in2(N__26673),
            .in3(N__26662),
            .lcout(n14136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_4_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_4_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_4_25_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1795_3_lut_LC_4_25_0 (
            .in0(_gnd_net_),
            .in1(N__28502),
            .in2(N__26640),
            .in3(N__33310),
            .lcout(n2731),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_4_25_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_4_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_4_25_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1794_3_lut_LC_4_25_1 (
            .in0(_gnd_net_),
            .in1(N__28550),
            .in2(N__33342),
            .in3(N__26625),
            .lcout(n2730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_27_LC_4_25_2.C_ON=1'b0;
    defparam i1_4_lut_adj_27_LC_4_25_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_27_LC_4_25_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_27_LC_4_25_2 (
            .in0(N__27868),
            .in1(N__26779),
            .in2(N__30697),
            .in3(N__27091),
            .lcout(),
            .ltout(n14688_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_29_LC_4_25_3.C_ON=1'b0;
    defparam i1_4_lut_adj_29_LC_4_25_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_29_LC_4_25_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_29_LC_4_25_3 (
            .in0(N__26605),
            .in1(N__26818),
            .in2(N__26589),
            .in3(N__26586),
            .lcout(n14696),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_new_i0_LC_4_25_4 .C_ON=1'b0;
    defparam \quad_counter0.b_new_i0_LC_4_25_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_new_i0_LC_4_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.b_new_i0_LC_4_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26568),
            .lcout(\quad_counter0.b_new_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55775),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_4_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_4_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_4_25_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1793_3_lut_LC_4_25_6 (
            .in0(_gnd_net_),
            .in1(N__26550),
            .in2(N__26541),
            .in3(N__33314),
            .lcout(n2729),
            .ltout(n2729_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_148_LC_4_25_7.C_ON=1'b0;
    defparam i1_4_lut_adj_148_LC_4_25_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_148_LC_4_25_7.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_148_LC_4_25_7 (
            .in0(N__26497),
            .in1(N__26467),
            .in2(N__26448),
            .in3(N__26868),
            .lcout(n13796),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_4_26_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_4_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_4_26_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2062_3_lut_LC_4_26_2 (
            .in0(_gnd_net_),
            .in1(N__28878),
            .in2(N__26955),
            .in3(N__37210),
            .lcout(n3126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_4_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_4_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_4_26_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1797_3_lut_LC_4_26_3 (
            .in0(N__26940),
            .in1(N__40125),
            .in2(_gnd_net_),
            .in3(N__33330),
            .lcout(n2733),
            .ltout(n2733_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9968_3_lut_LC_4_26_4.C_ON=1'b0;
    defparam i9968_3_lut_LC_4_26_4.SEQ_MODE=4'b0000;
    defparam i9968_3_lut_LC_4_26_4.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9968_3_lut_LC_4_26_4 (
            .in0(_gnd_net_),
            .in1(N__44871),
            .in2(N__26904),
            .in3(N__26894),
            .lcout(n11936),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12585_1_lut_LC_4_26_5.C_ON=1'b0;
    defparam i12585_1_lut_LC_4_26_5.SEQ_MODE=4'b0000;
    defparam i12585_1_lut_LC_4_26_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12585_1_lut_LC_4_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33511),
            .lcout(n15310),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_4_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_4_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_4_26_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1860_3_lut_LC_4_26_7 (
            .in0(N__26855),
            .in1(_gnd_net_),
            .in2(N__26841),
            .in3(N__33510),
            .lcout(n2828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_4_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_4_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_4_27_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1918_3_lut_LC_4_27_0 (
            .in0(_gnd_net_),
            .in1(N__26822),
            .in2(N__26802),
            .in3(N__33662),
            .lcout(n2918),
            .ltout(n2918_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_4_27_1.C_ON=1'b0;
    defparam i1_3_lut_LC_4_27_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_4_27_1.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_LC_4_27_1 (
            .in0(_gnd_net_),
            .in1(N__28975),
            .in2(N__26790),
            .in3(N__27367),
            .lcout(n14350),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_4_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_4_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_4_27_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1926_3_lut_LC_4_27_2 (
            .in0(_gnd_net_),
            .in1(N__26783),
            .in2(N__26763),
            .in3(N__33663),
            .lcout(n2926),
            .ltout(n2926_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_42_LC_4_27_3.C_ON=1'b0;
    defparam i1_2_lut_adj_42_LC_4_27_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_42_LC_4_27_3.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_42_LC_4_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27120),
            .in3(N__27193),
            .lcout(),
            .ltout(n14336_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_44_LC_4_27_4.C_ON=1'b0;
    defparam i1_4_lut_adj_44_LC_4_27_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_44_LC_4_27_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_44_LC_4_27_4 (
            .in0(N__30664),
            .in1(N__27117),
            .in2(N__27111),
            .in3(N__27833),
            .lcout(),
            .ltout(n14352_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_45_LC_4_27_5.C_ON=1'b0;
    defparam i1_4_lut_adj_45_LC_4_27_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_45_LC_4_27_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_45_LC_4_27_5 (
            .in0(N__27469),
            .in1(N__29360),
            .in2(N__27108),
            .in3(N__27105),
            .lcout(n14358),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_4_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_4_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_4_27_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1927_3_lut_LC_4_27_6 (
            .in0(_gnd_net_),
            .in1(N__27095),
            .in2(N__27075),
            .in3(N__33661),
            .lcout(n2927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_4_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_4_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_4_27_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1917_3_lut_LC_4_27_7 (
            .in0(N__27060),
            .in1(_gnd_net_),
            .in2(N__33699),
            .in3(N__27048),
            .lcout(n2917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_4_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_4_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_4_28_0.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1913_3_lut_LC_4_28_0 (
            .in0(N__27021),
            .in1(_gnd_net_),
            .in2(N__27012),
            .in3(N__33676),
            .lcout(n2913),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_46_LC_4_28_1.C_ON=1'b0;
    defparam i1_4_lut_adj_46_LC_4_28_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_46_LC_4_28_1.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_46_LC_4_28_1 (
            .in0(N__27160),
            .in1(N__27283),
            .in2(N__26985),
            .in3(N__26970),
            .lcout(),
            .ltout(n14360_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_47_LC_4_28_2.C_ON=1'b0;
    defparam i1_4_lut_adj_47_LC_4_28_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_47_LC_4_28_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_47_LC_4_28_2 (
            .in0(N__27610),
            .in1(N__27790),
            .in2(N__26964),
            .in3(N__27751),
            .lcout(n14366),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i0_LC_4_28_3 .C_ON=1'b0;
    defparam \debounce.reg_B_i0_LC_4_28_3 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i0_LC_4_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounce.reg_B_i0_LC_4_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34874),
            .lcout(reg_B_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55782),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_4_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_4_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_4_28_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1994_3_lut_LC_4_28_4 (
            .in0(_gnd_net_),
            .in1(N__27371),
            .in2(N__27351),
            .in3(N__33795),
            .lcout(n3026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12657_4_lut_LC_4_28_5.C_ON=1'b0;
    defparam i12657_4_lut_LC_4_28_5.SEQ_MODE=4'b0000;
    defparam i12657_4_lut_LC_4_28_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12657_4_lut_LC_4_28_5 (
            .in0(N__27334),
            .in1(N__28075),
            .in2(N__27315),
            .in3(N__27291),
            .lcout(n2940),
            .ltout(n2940_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_4_28_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_4_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_4_28_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1996_3_lut_LC_4_28_6 (
            .in0(N__27284),
            .in1(_gnd_net_),
            .in2(N__27264),
            .in3(N__27261),
            .lcout(n3028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_4_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_4_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_4_29_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1988_3_lut_LC_4_29_0 (
            .in0(_gnd_net_),
            .in1(N__27248),
            .in2(N__33850),
            .in3(N__27228),
            .lcout(n3020),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_4_29_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_4_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_4_29_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2051_3_lut_LC_4_29_1 (
            .in0(_gnd_net_),
            .in1(N__27642),
            .in2(N__37223),
            .in3(N__27216),
            .lcout(n3115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_4_29_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_4_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_4_29_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1995_3_lut_LC_4_29_2 (
            .in0(N__27207),
            .in1(_gnd_net_),
            .in2(N__33849),
            .in3(N__27197),
            .lcout(n3027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_4_29_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_4_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_4_29_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1997_3_lut_LC_4_29_3 (
            .in0(_gnd_net_),
            .in1(N__27177),
            .in2(N__27168),
            .in3(N__33803),
            .lcout(n3029),
            .ltout(n3029_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_4_29_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_4_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_4_29_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2064_3_lut_LC_4_29_4 (
            .in0(_gnd_net_),
            .in1(N__27144),
            .in2(N__27138),
            .in3(N__37211),
            .lcout(n3128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_4_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_4_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_4_29_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1991_3_lut_LC_4_29_5 (
            .in0(_gnd_net_),
            .in1(N__27829),
            .in2(N__27135),
            .in3(N__33804),
            .lcout(n3023),
            .ltout(n3023_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_68_LC_4_29_6.C_ON=1'b0;
    defparam i1_4_lut_adj_68_LC_4_29_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_68_LC_4_29_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_68_LC_4_29_6 (
            .in0(N__27400),
            .in1(N__27571),
            .in2(N__27555),
            .in3(N__28851),
            .lcout(n14738),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_4_29_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_4_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_4_29_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1989_3_lut_LC_4_29_7 (
            .in0(_gnd_net_),
            .in1(N__27552),
            .in2(N__27528),
            .in3(N__33796),
            .lcout(n3021),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_4_30_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_4_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_4_30_0.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i2046_3_lut_LC_4_30_0 (
            .in0(N__37153),
            .in1(_gnd_net_),
            .in2(N__27513),
            .in3(N__29208),
            .lcout(n3110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_4_30_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_4_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_4_30_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2043_3_lut_LC_4_30_1 (
            .in0(_gnd_net_),
            .in1(N__27504),
            .in2(N__29637),
            .in3(N__37154),
            .lcout(n3107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_4_30_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_4_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_4_30_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1984_3_lut_LC_4_30_2 (
            .in0(_gnd_net_),
            .in1(N__27495),
            .in2(N__27483),
            .in3(N__33858),
            .lcout(n3016),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_4_30_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_4_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_4_30_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1998_3_lut_LC_4_30_4 (
            .in0(_gnd_net_),
            .in1(N__27453),
            .in2(N__27429),
            .in3(N__33854),
            .lcout(n3030),
            .ltout(n3030_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_4_30_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_4_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_4_30_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2065_3_lut_LC_4_30_5 (
            .in0(_gnd_net_),
            .in1(N__27414),
            .in2(N__27408),
            .in3(N__37149),
            .lcout(n3129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_4_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_4_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_4_30_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2055_3_lut_LC_4_30_6 (
            .in0(_gnd_net_),
            .in1(N__27404),
            .in2(N__37203),
            .in3(N__27384),
            .lcout(n3119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_4_30_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_4_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_4_30_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1985_3_lut_LC_4_30_7 (
            .in0(N__27945),
            .in1(_gnd_net_),
            .in2(N__33887),
            .in3(N__27932),
            .lcout(n3017),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_4_31_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_4_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_4_31_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1978_3_lut_LC_4_31_0 (
            .in0(N__27912),
            .in1(N__27894),
            .in2(_gnd_net_),
            .in3(N__33873),
            .lcout(n3010),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_4_31_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_4_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_4_31_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1924_3_lut_LC_4_31_1 (
            .in0(N__27884),
            .in1(_gnd_net_),
            .in2(N__27852),
            .in3(N__33705),
            .lcout(n2924),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_4_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_4_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_4_31_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1980_3_lut_LC_4_31_2 (
            .in0(_gnd_net_),
            .in1(N__27800),
            .in2(N__27774),
            .in3(N__33871),
            .lcout(n3012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_4_31_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_4_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_4_31_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1982_3_lut_LC_4_31_4 (
            .in0(_gnd_net_),
            .in1(N__27761),
            .in2(N__27732),
            .in3(N__33867),
            .lcout(n3014),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_4_31_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_4_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_4_31_5.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1979_3_lut_LC_4_31_5 (
            .in0(N__27720),
            .in1(N__27696),
            .in2(N__33891),
            .in3(_gnd_net_),
            .lcout(n3011),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_4_31_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_4_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_4_31_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1986_3_lut_LC_4_31_6 (
            .in0(_gnd_net_),
            .in1(N__27687),
            .in2(N__27657),
            .in3(N__33872),
            .lcout(n3018),
            .ltout(n3018_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_164_LC_4_31_7.C_ON=1'b0;
    defparam i1_3_lut_adj_164_LC_4_31_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_164_LC_4_31_7.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_164_LC_4_31_7 (
            .in0(_gnd_net_),
            .in1(N__27640),
            .in2(N__27624),
            .in3(N__29170),
            .lcout(n14816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_4_32_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_4_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_4_32_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1981_3_lut_LC_4_32_0 (
            .in0(_gnd_net_),
            .in1(N__27621),
            .in2(N__27594),
            .in3(N__33892),
            .lcout(n3013),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12687_1_lut_LC_4_32_1.C_ON=1'b0;
    defparam i12687_1_lut_LC_4_32_1.SEQ_MODE=4'b0000;
    defparam i12687_1_lut_LC_4_32_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12687_1_lut_LC_4_32_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37171),
            .lcout(n15412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_4_32_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_4_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_4_32_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1975_3_lut_LC_4_32_2 (
            .in0(_gnd_net_),
            .in1(N__28085),
            .in2(N__28056),
            .in3(N__33894),
            .lcout(n3007),
            .ltout(n3007_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_4_32_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_4_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_4_32_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2042_3_lut_LC_4_32_3 (
            .in0(_gnd_net_),
            .in1(N__28044),
            .in2(N__28038),
            .in3(N__37172),
            .lcout(n3106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_4_32_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_4_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_4_32_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1977_3_lut_LC_4_32_6 (
            .in0(_gnd_net_),
            .in1(N__28035),
            .in2(N__28008),
            .in3(N__33893),
            .lcout(n3009),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i3_4_lut_LC_4_32_7 .C_ON=1'b0;
    defparam \debounce.i3_4_lut_LC_4_32_7 .SEQ_MODE=4'b0000;
    defparam \debounce.i3_4_lut_LC_4_32_7 .LUT_INIT=16'b1111011011111111;
    LogicCell40 \debounce.i3_4_lut_LC_4_32_7  (
            .in0(N__39554),
            .in1(N__27995),
            .in2(N__34809),
            .in3(N__39516),
            .lcout(\debounce.cnt_next_9__N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_5_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_5_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_5_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_2_lut_LC_5_17_0 (
            .in0(_gnd_net_),
            .in1(N__32184),
            .in2(_gnd_net_),
            .in3(N__27954),
            .lcout(n2201),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(n12643),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_5_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_5_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_5_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_3_lut_LC_5_17_1 (
            .in0(_gnd_net_),
            .in1(N__54403),
            .in2(N__32214),
            .in3(N__27951),
            .lcout(n2200),
            .ltout(),
            .carryin(n12643),
            .carryout(n12644),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_5_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_5_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_5_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_4_lut_LC_5_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32460),
            .in3(N__27948),
            .lcout(n2199),
            .ltout(),
            .carryin(n12644),
            .carryout(n12645),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_5_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_5_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_5_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_5_lut_LC_5_17_3 (
            .in0(_gnd_net_),
            .in1(N__54404),
            .in2(N__31970),
            .in3(N__28116),
            .lcout(n2198),
            .ltout(),
            .carryin(n12645),
            .carryout(n12646),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_5_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_5_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_5_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_6_lut_LC_5_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31998),
            .in3(N__28113),
            .lcout(n2197),
            .ltout(),
            .carryin(n12646),
            .carryout(n12647),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_5_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_5_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_5_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_7_lut_LC_5_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31936),
            .in3(N__28110),
            .lcout(n2196),
            .ltout(),
            .carryin(n12647),
            .carryout(n12648),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_5_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_5_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_5_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_8_lut_LC_5_17_6 (
            .in0(_gnd_net_),
            .in1(N__54406),
            .in2(N__31823),
            .in3(N__28107),
            .lcout(n2195),
            .ltout(),
            .carryin(n12648),
            .carryout(n12649),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_5_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_5_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_5_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_9_lut_LC_5_17_7 (
            .in0(_gnd_net_),
            .in1(N__54405),
            .in2(N__32289),
            .in3(N__28104),
            .lcout(n2194),
            .ltout(),
            .carryin(n12649),
            .carryout(n12650),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_5_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_5_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_5_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_10_lut_LC_5_18_0 (
            .in0(_gnd_net_),
            .in1(N__53562),
            .in2(N__31644),
            .in3(N__28101),
            .lcout(n2193),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(n12651),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_5_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_5_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_5_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_11_lut_LC_5_18_1 (
            .in0(_gnd_net_),
            .in1(N__53571),
            .in2(N__31848),
            .in3(N__28098),
            .lcout(n2192),
            .ltout(),
            .carryin(n12651),
            .carryout(n12652),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_5_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_5_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_5_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_12_lut_LC_5_18_2 (
            .in0(_gnd_net_),
            .in1(N__53563),
            .in2(N__31599),
            .in3(N__28095),
            .lcout(n2191),
            .ltout(),
            .carryin(n12652),
            .carryout(n12653),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_5_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_5_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_5_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_13_lut_LC_5_18_3 (
            .in0(_gnd_net_),
            .in1(N__53572),
            .in2(N__31670),
            .in3(N__28092),
            .lcout(n2190),
            .ltout(),
            .carryin(n12653),
            .carryout(n12654),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_5_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_5_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_5_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_14_lut_LC_5_18_4 (
            .in0(_gnd_net_),
            .in1(N__53564),
            .in2(N__31869),
            .in3(N__28089),
            .lcout(n2189),
            .ltout(),
            .carryin(n12654),
            .carryout(n12655),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_5_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_5_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_5_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_15_lut_LC_5_18_5 (
            .in0(_gnd_net_),
            .in1(N__31752),
            .in2(N__53933),
            .in3(N__28188),
            .lcout(n2188),
            .ltout(),
            .carryin(n12655),
            .carryout(n12656),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_5_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_5_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_5_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_16_lut_LC_5_18_6 (
            .in0(_gnd_net_),
            .in1(N__31793),
            .in2(N__53935),
            .in3(N__28185),
            .lcout(n2187),
            .ltout(),
            .carryin(n12656),
            .carryout(n12657),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_5_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_5_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_5_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_17_lut_LC_5_18_7 (
            .in0(_gnd_net_),
            .in1(N__31904),
            .in2(N__53934),
            .in3(N__28182),
            .lcout(n2186),
            .ltout(),
            .carryin(n12657),
            .carryout(n12658),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_5_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_5_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_5_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_18_lut_LC_5_19_0 (
            .in0(_gnd_net_),
            .in1(N__32061),
            .in2(N__54181),
            .in3(N__28179),
            .lcout(n2185),
            .ltout(),
            .carryin(bfn_5_19_0_),
            .carryout(n12659),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_5_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_5_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_5_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_19_lut_LC_5_19_1 (
            .in0(_gnd_net_),
            .in1(N__29957),
            .in2(N__54183),
            .in3(N__28176),
            .lcout(n2184),
            .ltout(),
            .carryin(n12659),
            .carryout(n12660),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_5_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_5_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_5_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_20_lut_LC_5_19_2 (
            .in0(_gnd_net_),
            .in1(N__30030),
            .in2(N__54182),
            .in3(N__28173),
            .lcout(n2183),
            .ltout(),
            .carryin(n12660),
            .carryout(n12661),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_5_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_5_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_5_19_3.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1436_21_lut_LC_5_19_3 (
            .in0(N__53915),
            .in1(N__34184),
            .in2(N__31698),
            .in3(N__28170),
            .lcout(n2214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_5_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_5_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_5_19_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1507_3_lut_LC_5_19_5 (
            .in0(N__29939),
            .in1(_gnd_net_),
            .in2(N__32655),
            .in3(N__28419),
            .lcout(n2315),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_5_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_5_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_5_19_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1517_3_lut_LC_5_19_6 (
            .in0(_gnd_net_),
            .in1(N__32250),
            .in2(N__28311),
            .in3(N__32614),
            .lcout(n2325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_5_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_5_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_5_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1451_3_lut_LC_5_19_7 (
            .in0(_gnd_net_),
            .in1(N__28257),
            .in2(N__31824),
            .in3(N__34127),
            .lcout(n2227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_5_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_5_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_5_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_2_lut_LC_5_20_0 (
            .in0(_gnd_net_),
            .in1(N__32036),
            .in2(_gnd_net_),
            .in3(N__28248),
            .lcout(n2301),
            .ltout(),
            .carryin(bfn_5_20_0_),
            .carryout(n12662),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_5_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_5_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_5_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_3_lut_LC_5_20_1 (
            .in0(_gnd_net_),
            .in1(N__53902),
            .in2(N__32145),
            .in3(N__28245),
            .lcout(n2300),
            .ltout(),
            .carryin(n12662),
            .carryout(n12663),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_5_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_5_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_5_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_4_lut_LC_5_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32097),
            .in3(N__28242),
            .lcout(n2299),
            .ltout(),
            .carryin(n12663),
            .carryout(n12664),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_5_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_5_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_5_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_5_lut_LC_5_20_3 (
            .in0(_gnd_net_),
            .in1(N__53903),
            .in2(N__32123),
            .in3(N__28239),
            .lcout(n2298),
            .ltout(),
            .carryin(n12664),
            .carryout(n12665),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_5_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_5_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_5_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_6_lut_LC_5_20_4 (
            .in0(_gnd_net_),
            .in1(N__28334),
            .in2(_gnd_net_),
            .in3(N__28224),
            .lcout(n2297),
            .ltout(),
            .carryin(n12665),
            .carryout(n12666),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_5_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_5_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_5_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_7_lut_LC_5_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30002),
            .in3(N__28212),
            .lcout(n2296),
            .ltout(),
            .carryin(n12666),
            .carryout(n12667),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_5_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_5_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_5_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_8_lut_LC_5_20_6 (
            .in0(_gnd_net_),
            .in1(N__53905),
            .in2(N__30506),
            .in3(N__28200),
            .lcout(n2295),
            .ltout(),
            .carryin(n12667),
            .carryout(n12668),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_5_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_5_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_5_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_9_lut_LC_5_20_7 (
            .in0(_gnd_net_),
            .in1(N__53904),
            .in2(N__30453),
            .in3(N__28314),
            .lcout(n2294),
            .ltout(),
            .carryin(n12668),
            .carryout(n12669),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_5_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_5_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_5_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_10_lut_LC_5_21_0 (
            .in0(_gnd_net_),
            .in1(N__53890),
            .in2(N__32249),
            .in3(N__28299),
            .lcout(n2293),
            .ltout(),
            .carryin(bfn_5_21_0_),
            .carryout(n12670),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_5_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_5_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_5_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_11_lut_LC_5_21_1 (
            .in0(_gnd_net_),
            .in1(N__53896),
            .in2(N__30426),
            .in3(N__28296),
            .lcout(n2292),
            .ltout(),
            .carryin(n12670),
            .carryout(n12671),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_5_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_5_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_5_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_12_lut_LC_5_21_2 (
            .in0(_gnd_net_),
            .in1(N__53891),
            .in2(N__30474),
            .in3(N__28293),
            .lcout(n2291),
            .ltout(),
            .carryin(n12671),
            .carryout(n12672),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_5_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_5_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_5_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_13_lut_LC_5_21_3 (
            .in0(_gnd_net_),
            .in1(N__53897),
            .in2(N__30405),
            .in3(N__28290),
            .lcout(n2290),
            .ltout(),
            .carryin(n12672),
            .carryout(n12673),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_5_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_5_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_5_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_14_lut_LC_5_21_4 (
            .in0(_gnd_net_),
            .in1(N__53892),
            .in2(N__30381),
            .in3(N__28287),
            .lcout(n2289),
            .ltout(),
            .carryin(n12673),
            .carryout(n12674),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_5_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_5_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_5_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_15_lut_LC_5_21_5 (
            .in0(_gnd_net_),
            .in1(N__53898),
            .in2(N__30353),
            .in3(N__28278),
            .lcout(n2288),
            .ltout(),
            .carryin(n12674),
            .carryout(n12675),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_5_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_5_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_5_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_16_lut_LC_5_21_6 (
            .in0(_gnd_net_),
            .in1(N__30320),
            .in2(N__54180),
            .in3(N__28269),
            .lcout(n2287),
            .ltout(),
            .carryin(n12675),
            .carryout(n12676),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_5_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_5_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_5_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_17_lut_LC_5_21_7 (
            .in0(_gnd_net_),
            .in1(N__30146),
            .in2(N__54179),
            .in3(N__28260),
            .lcout(n2286),
            .ltout(),
            .carryin(n12676),
            .carryout(n12677),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_5_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_5_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_5_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_18_lut_LC_5_22_0 (
            .in0(_gnd_net_),
            .in1(N__53491),
            .in2(N__30177),
            .in3(N__28425),
            .lcout(n2285),
            .ltout(),
            .carryin(bfn_5_22_0_),
            .carryout(n12678),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_5_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_5_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_5_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_19_lut_LC_5_22_1 (
            .in0(_gnd_net_),
            .in1(N__32522),
            .in2(N__53888),
            .in3(N__28422),
            .lcout(n2284),
            .ltout(),
            .carryin(n12678),
            .carryout(n12679),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_5_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_5_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_5_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_20_lut_LC_5_22_2 (
            .in0(_gnd_net_),
            .in1(N__29940),
            .in2(N__53921),
            .in3(N__28410),
            .lcout(n2283),
            .ltout(),
            .carryin(n12679),
            .carryout(n12680),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_5_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_5_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_5_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_21_lut_LC_5_22_3 (
            .in0(_gnd_net_),
            .in1(N__29924),
            .in2(N__53889),
            .in3(N__28395),
            .lcout(n2282),
            .ltout(),
            .carryin(n12680),
            .carryout(n12681),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_5_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_5_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_5_22_4.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1503_22_lut_LC_5_22_4 (
            .in0(N__53546),
            .in1(N__29901),
            .in2(N__32702),
            .in3(N__28392),
            .lcout(n2313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_5_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_5_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_5_22_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1523_3_lut_LC_5_22_5 (
            .in0(_gnd_net_),
            .in1(N__28368),
            .in2(N__32671),
            .in3(N__32096),
            .lcout(n2331),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_5_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_5_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_5_23_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1452_3_lut_LC_5_23_1 (
            .in0(_gnd_net_),
            .in1(N__28359),
            .in2(N__31944),
            .in3(N__34159),
            .lcout(n2228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_5_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_5_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_5_23_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1454_3_lut_LC_5_23_3 (
            .in0(_gnd_net_),
            .in1(N__28347),
            .in2(N__31977),
            .in3(N__34160),
            .lcout(n2230),
            .ltout(n2230_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_103_LC_5_23_4.C_ON=1'b0;
    defparam i1_2_lut_adj_103_LC_5_23_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_103_LC_5_23_4.LUT_INIT=16'b1010000010100000;
    LogicCell40 i1_2_lut_adj_103_LC_5_23_4 (
            .in0(N__30001),
            .in1(_gnd_net_),
            .in2(N__28317),
            .in3(_gnd_net_),
            .lcout(n14812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_5_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_5_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_5_23_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1513_3_lut_LC_5_23_5 (
            .in0(N__30380),
            .in1(_gnd_net_),
            .in2(N__32684),
            .in3(N__28764),
            .lcout(n2321),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9986_4_lut_LC_5_23_7.C_ON=1'b0;
    defparam i9986_4_lut_LC_5_23_7.SEQ_MODE=4'b0000;
    defparam i9986_4_lut_LC_5_23_7.LUT_INIT=16'b1111110011111000;
    LogicCell40 i9986_4_lut_LC_5_23_7 (
            .in0(N__30565),
            .in1(N__30077),
            .in2(N__28705),
            .in3(N__28441),
            .lcout(n11954),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_5_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_5_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_5_24_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i9_3_lut_LC_5_24_0 (
            .in0(N__38499),
            .in1(N__46182),
            .in2(_gnd_net_),
            .in3(N__36666),
            .lcout(n311),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_5_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_5_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_5_24_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1728_3_lut_LC_5_24_1 (
            .in0(_gnd_net_),
            .in1(N__28638),
            .in2(N__28605),
            .in3(N__33163),
            .lcout(n2632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_5_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_5_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_5_24_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_5_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36665),
            .lcout(n25_adj_646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_5_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_5_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_5_24_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1727_3_lut_LC_5_24_3 (
            .in0(_gnd_net_),
            .in1(N__28590),
            .in2(N__28566),
            .in3(N__33164),
            .lcout(n2631),
            .ltout(n2631_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10076_4_lut_LC_5_24_4.C_ON=1'b0;
    defparam i10076_4_lut_LC_5_24_4.SEQ_MODE=4'b0000;
    defparam i10076_4_lut_LC_5_24_4.LUT_INIT=16'b1111111011110000;
    LogicCell40 i10076_4_lut_LC_5_24_4 (
            .in0(N__40121),
            .in1(N__28536),
            .in2(N__28506),
            .in3(N__28498),
            .lcout(n12044),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_5_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_5_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_5_24_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1525_3_lut_LC_5_24_6 (
            .in0(N__32037),
            .in1(_gnd_net_),
            .in2(N__28470),
            .in3(N__32672),
            .lcout(n2333),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_5_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_5_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_5_24_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_5_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36570),
            .lcout(n20_adj_641),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_5_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_5_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_5_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_2_lut_LC_5_25_0 (
            .in0(_gnd_net_),
            .in1(N__40054),
            .in2(_gnd_net_),
            .in3(N__28791),
            .lcout(n3201),
            .ltout(),
            .carryin(bfn_5_25_0_),
            .carryout(n12878),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_5_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_5_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_5_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_3_lut_LC_5_25_1 (
            .in0(_gnd_net_),
            .in1(N__53251),
            .in2(N__36933),
            .in3(N__28788),
            .lcout(n3200),
            .ltout(),
            .carryin(n12878),
            .carryout(n12879),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_5_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_5_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_5_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_4_lut_LC_5_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36906),
            .in3(N__28785),
            .lcout(n3199),
            .ltout(),
            .carryin(n12879),
            .carryout(n12880),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_5_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_5_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_5_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_5_lut_LC_5_25_3 (
            .in0(_gnd_net_),
            .in1(N__53252),
            .in2(N__36798),
            .in3(N__28782),
            .lcout(n3198),
            .ltout(),
            .carryin(n12880),
            .carryout(n12881),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_5_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_5_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_5_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_6_lut_LC_5_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36836),
            .in3(N__28779),
            .lcout(n3197),
            .ltout(),
            .carryin(n12881),
            .carryout(n12882),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_5_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_5_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_5_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_7_lut_LC_5_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36876),
            .in3(N__28776),
            .lcout(n3196),
            .ltout(),
            .carryin(n12882),
            .carryout(n12883),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_5_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_5_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_5_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_8_lut_LC_5_25_6 (
            .in0(_gnd_net_),
            .in1(N__53254),
            .in2(N__34545),
            .in3(N__28773),
            .lcout(n3195),
            .ltout(),
            .carryin(n12883),
            .carryout(n12884),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_5_25_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_5_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_5_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_9_lut_LC_5_25_7 (
            .in0(_gnd_net_),
            .in1(N__53253),
            .in2(N__34361),
            .in3(N__28770),
            .lcout(n3194),
            .ltout(),
            .carryin(n12884),
            .carryout(n12885),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_5_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_5_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_5_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_10_lut_LC_5_26_0 (
            .in0(_gnd_net_),
            .in1(N__53003),
            .in2(N__34243),
            .in3(N__28767),
            .lcout(n3193),
            .ltout(),
            .carryin(bfn_5_26_0_),
            .carryout(n12886),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_5_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_5_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_5_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_11_lut_LC_5_26_1 (
            .in0(_gnd_net_),
            .in1(N__53008),
            .in2(N__34920),
            .in3(N__28818),
            .lcout(n3192),
            .ltout(),
            .carryin(n12886),
            .carryout(n12887),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_5_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_5_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_5_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_12_lut_LC_5_26_2 (
            .in0(_gnd_net_),
            .in1(N__30953),
            .in2(N__53386),
            .in3(N__28815),
            .lcout(n3191),
            .ltout(),
            .carryin(n12887),
            .carryout(n12888),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_5_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_5_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_5_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_13_lut_LC_5_26_3 (
            .in0(_gnd_net_),
            .in1(N__53012),
            .in2(N__37044),
            .in3(N__28812),
            .lcout(n3190),
            .ltout(),
            .carryin(n12888),
            .carryout(n12889),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_5_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_5_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_5_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_14_lut_LC_5_26_4 (
            .in0(_gnd_net_),
            .in1(N__31138),
            .in2(N__53387),
            .in3(N__28809),
            .lcout(n3189),
            .ltout(),
            .carryin(n12889),
            .carryout(n12890),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_5_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_5_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_5_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_15_lut_LC_5_26_5 (
            .in0(_gnd_net_),
            .in1(N__53016),
            .in2(N__31005),
            .in3(N__28806),
            .lcout(n3188),
            .ltout(),
            .carryin(n12890),
            .carryout(n12891),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_5_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_5_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_5_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_16_lut_LC_5_26_6 (
            .in0(_gnd_net_),
            .in1(N__53004),
            .in2(N__31458),
            .in3(N__28803),
            .lcout(n3187),
            .ltout(),
            .carryin(n12891),
            .carryout(n12892),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_5_26_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_5_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_5_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_17_lut_LC_5_26_7 (
            .in0(_gnd_net_),
            .in1(N__34457),
            .in2(N__53385),
            .in3(N__28800),
            .lcout(n3186),
            .ltout(),
            .carryin(n12892),
            .carryout(n12893),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_5_27_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_5_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_5_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_18_lut_LC_5_27_0 (
            .in0(_gnd_net_),
            .in1(N__34780),
            .in2(N__54286),
            .in3(N__28797),
            .lcout(n3185),
            .ltout(),
            .carryin(bfn_5_27_0_),
            .carryout(n12894),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_5_27_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_5_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_5_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_19_lut_LC_5_27_1 (
            .in0(_gnd_net_),
            .in1(N__54102),
            .in2(N__34496),
            .in3(N__28794),
            .lcout(n3184),
            .ltout(),
            .carryin(n12894),
            .carryout(n12895),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_5_27_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_5_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_5_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_20_lut_LC_5_27_2 (
            .in0(_gnd_net_),
            .in1(N__30755),
            .in2(N__54287),
            .in3(N__28845),
            .lcout(n3183),
            .ltout(),
            .carryin(n12895),
            .carryout(n12896),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_5_27_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_5_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_5_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_21_lut_LC_5_27_3 (
            .in0(_gnd_net_),
            .in1(N__31076),
            .in2(N__54290),
            .in3(N__28842),
            .lcout(n3182),
            .ltout(),
            .carryin(n12896),
            .carryout(n12897),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_5_27_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_5_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_5_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_22_lut_LC_5_27_4 (
            .in0(_gnd_net_),
            .in1(N__31050),
            .in2(N__54288),
            .in3(N__28839),
            .lcout(n3181),
            .ltout(),
            .carryin(n12897),
            .carryout(n12898),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_5_27_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_5_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_5_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_23_lut_LC_5_27_5 (
            .in0(_gnd_net_),
            .in1(N__30921),
            .in2(N__54291),
            .in3(N__28836),
            .lcout(n3180),
            .ltout(),
            .carryin(n12898),
            .carryout(n12899),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_5_27_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_5_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_5_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_24_lut_LC_5_27_6 (
            .in0(_gnd_net_),
            .in1(N__34956),
            .in2(N__54289),
            .in3(N__28833),
            .lcout(n3179),
            .ltout(),
            .carryin(n12899),
            .carryout(n12900),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_5_27_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_5_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_5_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_25_lut_LC_5_27_7 (
            .in0(_gnd_net_),
            .in1(N__31201),
            .in2(N__54292),
            .in3(N__28830),
            .lcout(n3178),
            .ltout(),
            .carryin(n12900),
            .carryout(n12901),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_5_28_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_5_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_5_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_26_lut_LC_5_28_0 (
            .in0(_gnd_net_),
            .in1(N__54121),
            .in2(N__34292),
            .in3(N__28827),
            .lcout(n3177),
            .ltout(),
            .carryin(bfn_5_28_0_),
            .carryout(n12902),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_5_28_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_5_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_5_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_27_lut_LC_5_28_1 (
            .in0(_gnd_net_),
            .in1(N__43226),
            .in2(N__54293),
            .in3(N__28824),
            .lcout(n3176),
            .ltout(),
            .carryin(n12902),
            .carryout(n12903),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_5_28_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_5_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_5_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_28_lut_LC_5_28_2 (
            .in0(_gnd_net_),
            .in1(N__30893),
            .in2(N__54295),
            .in3(N__28821),
            .lcout(n3175),
            .ltout(),
            .carryin(n12903),
            .carryout(n12904),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_5_28_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_5_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_5_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_29_lut_LC_5_28_3 (
            .in0(_gnd_net_),
            .in1(N__30816),
            .in2(N__54294),
            .in3(N__29007),
            .lcout(n3174),
            .ltout(),
            .carryin(n12904),
            .carryout(n12905),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_5_28_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_5_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_5_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_30_lut_LC_5_28_4 (
            .in0(_gnd_net_),
            .in1(N__30848),
            .in2(N__54296),
            .in3(N__29004),
            .lcout(n3173),
            .ltout(),
            .carryin(n12905),
            .carryout(n12906),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_5_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_5_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_5_28_5.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_2106_31_lut_LC_5_28_5 (
            .in0(N__30873),
            .in1(N__54134),
            .in2(N__32366),
            .in3(N__29001),
            .lcout(n3204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_5_28_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_5_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_5_28_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2116_3_lut_LC_5_28_6 (
            .in0(_gnd_net_),
            .in1(N__30919),
            .in2(N__28998),
            .in3(N__43146),
            .lcout(n3212),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_5_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_5_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_5_28_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1992_3_lut_LC_5_28_7 (
            .in0(_gnd_net_),
            .in1(N__28985),
            .in2(N__28959),
            .in3(N__33844),
            .lcout(n3024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_5_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_5_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_5_29_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2067_3_lut_LC_5_29_0 (
            .in0(N__29093),
            .in1(_gnd_net_),
            .in2(N__28944),
            .in3(N__37193),
            .lcout(n3131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_5_29_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_5_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_5_29_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i2044_3_lut_LC_5_29_1 (
            .in0(N__37195),
            .in1(_gnd_net_),
            .in2(N__28932),
            .in3(N__29673),
            .lcout(n3108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_5_29_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_5_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_5_29_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1993_3_lut_LC_5_29_2 (
            .in0(_gnd_net_),
            .in1(N__28913),
            .in2(N__28893),
            .in3(N__33865),
            .lcout(n3025),
            .ltout(n3025_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_67_LC_5_29_3.C_ON=1'b0;
    defparam i1_4_lut_adj_67_LC_5_29_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_67_LC_5_29_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_67_LC_5_29_3 (
            .in0(N__37255),
            .in1(N__28870),
            .in2(N__28854),
            .in3(N__29058),
            .lcout(n14736),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_5_29_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_5_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_5_29_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2049_3_lut_LC_5_29_4 (
            .in0(_gnd_net_),
            .in1(N__29175),
            .in2(N__29154),
            .in3(N__37194),
            .lcout(n3113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_5_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_5_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_5_29_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2068_3_lut_LC_5_29_5 (
            .in0(_gnd_net_),
            .in1(N__29114),
            .in2(N__37217),
            .in3(N__29139),
            .lcout(n3132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_5_29_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_5_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_5_29_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2001_3_lut_LC_5_29_6 (
            .in0(N__32425),
            .in1(_gnd_net_),
            .in2(N__29130),
            .in3(N__33866),
            .lcout(n3033),
            .ltout(n3033_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9964_3_lut_LC_5_29_7.C_ON=1'b0;
    defparam i9964_3_lut_LC_5_29_7.SEQ_MODE=4'b0000;
    defparam i9964_3_lut_LC_5_29_7.LUT_INIT=16'b1111101000000000;
    LogicCell40 i9964_3_lut_LC_5_29_7 (
            .in0(N__42220),
            .in1(_gnd_net_),
            .in2(N__29100),
            .in3(N__29092),
            .lcout(n11932),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_5_30_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_5_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_5_30_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1990_3_lut_LC_5_30_0 (
            .in0(_gnd_net_),
            .in1(N__30672),
            .in2(N__29073),
            .in3(N__33862),
            .lcout(n3022),
            .ltout(n3022_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_66_LC_5_30_1.C_ON=1'b0;
    defparam i1_4_lut_adj_66_LC_5_30_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_66_LC_5_30_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_66_LC_5_30_1 (
            .in0(N__29233),
            .in1(N__31489),
            .in2(N__29061),
            .in3(N__31384),
            .lcout(n14732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_69_LC_5_30_2.C_ON=1'b0;
    defparam i1_4_lut_adj_69_LC_5_30_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_69_LC_5_30_2.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_69_LC_5_30_2 (
            .in0(N__29048),
            .in1(N__29033),
            .in2(N__29396),
            .in3(N__29022),
            .lcout(),
            .ltout(n13859_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_70_LC_5_30_3.C_ON=1'b0;
    defparam i1_4_lut_adj_70_LC_5_30_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_70_LC_5_30_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_70_LC_5_30_3 (
            .in0(N__29306),
            .in1(N__29503),
            .in2(N__29016),
            .in3(N__29013),
            .lcout(n14744),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_5_30_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_5_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_5_30_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1999_3_lut_LC_5_30_4 (
            .in0(_gnd_net_),
            .in1(N__29436),
            .in2(N__29424),
            .in3(N__33863),
            .lcout(n3031),
            .ltout(n3031_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_5_30_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_5_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_5_30_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2066_3_lut_LC_5_30_5 (
            .in0(_gnd_net_),
            .in1(N__29376),
            .in2(N__29364),
            .in3(N__37155),
            .lcout(n3130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_5_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_5_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_5_30_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1983_3_lut_LC_5_30_6 (
            .in0(_gnd_net_),
            .in1(N__29361),
            .in2(N__29328),
            .in3(N__33864),
            .lcout(n3015),
            .ltout(n3015_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_5_30_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_5_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_5_30_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2050_3_lut_LC_5_30_7 (
            .in0(_gnd_net_),
            .in1(N__29295),
            .in2(N__29283),
            .in3(N__37156),
            .lcout(n3114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_5_31_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_5_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_5_31_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2057_3_lut_LC_5_31_1 (
            .in0(_gnd_net_),
            .in1(N__29280),
            .in2(N__29268),
            .in3(N__37158),
            .lcout(n3121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_5_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_5_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_5_31_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2063_3_lut_LC_5_31_2 (
            .in0(_gnd_net_),
            .in1(N__29247),
            .in2(N__37204),
            .in3(N__29234),
            .lcout(n3127),
            .ltout(n3127_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_32_LC_5_31_3.C_ON=1'b0;
    defparam i1_4_lut_adj_32_LC_5_31_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_32_LC_5_31_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_32_LC_5_31_3 (
            .in0(N__34444),
            .in1(N__34534),
            .in2(N__29211),
            .in3(N__34245),
            .lcout(n14196),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_101_LC_5_31_4.C_ON=1'b0;
    defparam i1_4_lut_adj_101_LC_5_31_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_101_LC_5_31_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_101_LC_5_31_4 (
            .in0(N__29206),
            .in1(N__34330),
            .in2(N__29571),
            .in3(N__29190),
            .lcout(),
            .ltout(n14750_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_165_LC_5_31_5.C_ON=1'b0;
    defparam i1_4_lut_adj_165_LC_5_31_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_165_LC_5_31_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_165_LC_5_31_5 (
            .in0(N__29184),
            .in1(N__29752),
            .in2(N__29178),
            .in3(N__29665),
            .lcout(),
            .ltout(n14754_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12690_4_lut_LC_5_31_6.C_ON=1'b0;
    defparam i12690_4_lut_LC_5_31_6.SEQ_MODE=4'b0000;
    defparam i12690_4_lut_LC_5_31_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12690_4_lut_LC_5_31_6 (
            .in0(N__29648),
            .in1(N__29633),
            .in2(N__29604),
            .in3(N__29601),
            .lcout(n3039),
            .ltout(n3039_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_5_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_5_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_5_31_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2047_3_lut_LC_5_31_7 (
            .in0(_gnd_net_),
            .in1(N__29583),
            .in2(N__29574),
            .in3(N__29569),
            .lcout(n3111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_30_LC_5_32_0.C_ON=1'b0;
    defparam i1_4_lut_adj_30_LC_5_32_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_30_LC_5_32_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_30_LC_5_32_0 (
            .in0(N__30946),
            .in1(N__34906),
            .in2(N__34782),
            .in3(N__31140),
            .lcout(),
            .ltout(n14194_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_33_LC_5_32_1.C_ON=1'b0;
    defparam i1_4_lut_adj_33_LC_5_32_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_33_LC_5_32_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_33_LC_5_32_1 (
            .in0(N__29514),
            .in1(N__30748),
            .in2(N__29553),
            .in3(N__29550),
            .lcout(n14204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_5_32_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_5_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_5_32_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i2053_3_lut_LC_5_32_2 (
            .in0(N__29544),
            .in1(_gnd_net_),
            .in2(N__37205),
            .in3(N__29529),
            .lcout(n3117),
            .ltout(n3117_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_31_LC_5_32_3.C_ON=1'b0;
    defparam i1_4_lut_adj_31_LC_5_32_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_31_LC_5_32_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_31_LC_5_32_3 (
            .in0(N__30988),
            .in1(N__31441),
            .in2(N__29517),
            .in3(N__37039),
            .lcout(n14198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_5_32_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_5_32_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_5_32_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2052_3_lut_LC_5_32_4 (
            .in0(_gnd_net_),
            .in1(N__29508),
            .in2(N__37206),
            .in3(N__29487),
            .lcout(n3116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_5_32_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_5_32_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_5_32_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2060_3_lut_LC_5_32_5 (
            .in0(_gnd_net_),
            .in1(N__29474),
            .in2(N__29451),
            .in3(N__37162),
            .lcout(n3124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_5_32_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_5_32_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_5_32_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2045_3_lut_LC_5_32_7 (
            .in0(N__29757),
            .in1(_gnd_net_),
            .in2(N__29736),
            .in3(N__37169),
            .lcout(n3109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_6_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_6_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_6_17_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1385_3_lut_LC_6_17_0 (
            .in0(_gnd_net_),
            .in1(N__31410),
            .in2(N__37974),
            .in3(N__34024),
            .lcout(n2129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12989_1_lut_LC_6_17_3.C_ON=1'b0;
    defparam i12989_1_lut_LC_6_17_3.SEQ_MODE=4'b0000;
    defparam i12989_1_lut_LC_6_17_3.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12989_1_lut_LC_6_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34169),
            .in3(_gnd_net_),
            .lcout(n15714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_6_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_6_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_6_17_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1387_3_lut_LC_6_17_6 (
            .in0(_gnd_net_),
            .in1(N__31422),
            .in2(N__38118),
            .in3(N__34025),
            .lcout(n2131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_6_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_6_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_6_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_6_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36608),
            .lcout(n21_adj_642),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_6_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_6_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_6_18_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1384_3_lut_LC_6_18_1 (
            .in0(_gnd_net_),
            .in1(N__31401),
            .in2(N__36174),
            .in3(N__33985),
            .lcout(n2128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_6_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_6_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_6_18_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1448_3_lut_LC_6_18_2 (
            .in0(N__31847),
            .in1(_gnd_net_),
            .in2(N__29724),
            .in3(N__34154),
            .lcout(n2224),
            .ltout(n2224_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_6_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_6_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_6_18_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1515_3_lut_LC_6_18_3 (
            .in0(_gnd_net_),
            .in1(N__29715),
            .in2(N__29706),
            .in3(N__32653),
            .lcout(n2323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_6_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_6_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_6_18_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1382_3_lut_LC_6_18_5 (
            .in0(_gnd_net_),
            .in1(N__31569),
            .in2(N__37677),
            .in3(N__33984),
            .lcout(n2126),
            .ltout(n2126_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1449_3_lut_LC_6_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1449_3_lut_LC_6_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1449_3_lut_LC_6_18_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1449_3_lut_LC_6_18_6 (
            .in0(_gnd_net_),
            .in1(N__29838),
            .in2(N__29832),
            .in3(N__34155),
            .lcout(n2225),
            .ltout(n2225_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1516_3_lut_LC_6_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1516_3_lut_LC_6_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1516_3_lut_LC_6_18_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1516_3_lut_LC_6_18_7 (
            .in0(_gnd_net_),
            .in1(N__29829),
            .in2(N__29820),
            .in3(N__32654),
            .lcout(n2324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_6_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_6_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_6_19_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1381_3_lut_LC_6_19_0 (
            .in0(_gnd_net_),
            .in1(N__31560),
            .in2(N__36372),
            .in3(N__34002),
            .lcout(n2125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_6_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_6_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_6_19_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1372_3_lut_LC_6_19_1 (
            .in0(N__36317),
            .in1(_gnd_net_),
            .in2(N__34027),
            .in3(N__31710),
            .lcout(n2116),
            .ltout(n2116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_6_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_6_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_6_19_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1439_3_lut_LC_6_19_2 (
            .in0(N__34153),
            .in1(_gnd_net_),
            .in2(N__29781),
            .in3(N__29778),
            .lcout(n2215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12967_4_lut_LC_6_19_3.C_ON=1'b0;
    defparam i12967_4_lut_LC_6_19_3.SEQ_MODE=4'b0000;
    defparam i12967_4_lut_LC_6_19_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12967_4_lut_LC_6_19_3 (
            .in0(N__36316),
            .in1(N__36092),
            .in2(N__31629),
            .in3(N__36435),
            .lcout(n2049),
            .ltout(n2049_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_6_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_6_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_6_19_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1379_3_lut_LC_6_19_4 (
            .in0(_gnd_net_),
            .in1(N__36203),
            .in2(N__29769),
            .in3(N__31548),
            .lcout(n2123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_6_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_6_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_6_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1442_3_lut_LC_6_19_5 (
            .in0(_gnd_net_),
            .in1(N__31905),
            .in2(N__29766),
            .in3(N__34152),
            .lcout(n2218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_6_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_6_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_6_19_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1376_3_lut_LC_6_19_6 (
            .in0(_gnd_net_),
            .in1(N__31533),
            .in2(N__38028),
            .in3(N__34003),
            .lcout(n2120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_6_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_6_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_6_19_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1375_3_lut_LC_6_19_7 (
            .in0(_gnd_net_),
            .in1(N__31524),
            .in2(N__34026),
            .in3(N__37886),
            .lcout(n2119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_6_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_6_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_6_20_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1514_3_lut_LC_6_20_0 (
            .in0(_gnd_net_),
            .in1(N__30403),
            .in2(N__30066),
            .in3(N__32613),
            .lcout(n2322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_6_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_6_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_6_20_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1373_3_lut_LC_6_20_1 (
            .in0(_gnd_net_),
            .in1(N__31628),
            .in2(N__31722),
            .in3(N__34015),
            .lcout(n2117),
            .ltout(n2117_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12992_4_lut_LC_6_20_2.C_ON=1'b0;
    defparam i12992_4_lut_LC_6_20_2.SEQ_MODE=4'b0000;
    defparam i12992_4_lut_LC_6_20_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12992_4_lut_LC_6_20_2 (
            .in0(N__31691),
            .in1(N__30029),
            .in2(N__30018),
            .in3(N__31884),
            .lcout(n2148),
            .ltout(n2148_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_6_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_6_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_6_20_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1453_3_lut_LC_6_20_3 (
            .in0(_gnd_net_),
            .in1(N__31991),
            .in2(N__30015),
            .in3(N__30012),
            .lcout(n2229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_6_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_6_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_6_20_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1445_3_lut_LC_6_20_4 (
            .in0(_gnd_net_),
            .in1(N__31862),
            .in2(N__29976),
            .in3(N__34148),
            .lcout(n2221),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_6_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_6_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_6_20_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1440_3_lut_LC_6_20_5 (
            .in0(N__29964),
            .in1(_gnd_net_),
            .in2(N__34168),
            .in3(N__29958),
            .lcout(n2216),
            .ltout(n2216_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13017_4_lut_LC_6_20_6.C_ON=1'b0;
    defparam i13017_4_lut_LC_6_20_6.SEQ_MODE=4'b0000;
    defparam i13017_4_lut_LC_6_20_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13017_4_lut_LC_6_20_6 (
            .in0(N__29923),
            .in1(N__29897),
            .in2(N__29886),
            .in3(N__30126),
            .lcout(n2247),
            .ltout(n2247_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_6_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_6_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_6_20_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1522_3_lut_LC_6_20_7 (
            .in0(N__29883),
            .in1(_gnd_net_),
            .in2(N__29877),
            .in3(N__32124),
            .lcout(n2330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_6_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_6_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_6_21_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1443_3_lut_LC_6_21_0 (
            .in0(N__30285),
            .in1(_gnd_net_),
            .in2(N__34162),
            .in3(N__31797),
            .lcout(n2219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_6_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_6_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_6_21_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1455_3_lut_LC_6_21_1 (
            .in0(_gnd_net_),
            .in1(N__32453),
            .in2(N__30276),
            .in3(N__34128),
            .lcout(n2231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_6_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_6_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_6_21_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1509_3_lut_LC_6_21_2 (
            .in0(N__30173),
            .in1(_gnd_net_),
            .in2(N__30261),
            .in3(N__32635),
            .lcout(n2317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_6_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_6_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_6_21_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1456_3_lut_LC_6_21_3 (
            .in0(_gnd_net_),
            .in1(N__32207),
            .in2(N__30216),
            .in3(N__34129),
            .lcout(n2232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_6_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_6_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_6_21_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1447_3_lut_LC_6_21_4 (
            .in0(_gnd_net_),
            .in1(N__31595),
            .in2(N__34161),
            .in3(N__30201),
            .lcout(n2223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_6_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_6_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_6_21_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1441_3_lut_LC_6_21_5 (
            .in0(_gnd_net_),
            .in1(N__32057),
            .in2(N__30192),
            .in3(N__34137),
            .lcout(n2217),
            .ltout(n2217_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_105_LC_6_21_6.C_ON=1'b0;
    defparam i1_4_lut_adj_105_LC_6_21_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_105_LC_6_21_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_105_LC_6_21_6 (
            .in0(N__30172),
            .in1(N__30145),
            .in2(N__30129),
            .in3(N__30291),
            .lcout(n14598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_6_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_6_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_6_21_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1444_3_lut_LC_6_21_7 (
            .in0(_gnd_net_),
            .in1(N__30120),
            .in2(N__31751),
            .in3(N__34133),
            .lcout(n2220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_6_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_6_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_6_22_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1524_3_lut_LC_6_22_0 (
            .in0(_gnd_net_),
            .in1(N__32138),
            .in2(N__30111),
            .in3(N__32636),
            .lcout(n2332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_6_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_6_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_6_22_1.LUT_INIT=16'b1101100011011000;
    LogicCell40 encoder0_position_31__I_0_i1446_3_lut_LC_6_22_1 (
            .in0(N__34163),
            .in1(N__31671),
            .in2(N__30522),
            .in3(_gnd_net_),
            .lcout(n2222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_99_LC_6_22_2.C_ON=1'b0;
    defparam i1_2_lut_adj_99_LC_6_22_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_99_LC_6_22_2.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_99_LC_6_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30499),
            .in3(N__30467),
            .lcout(),
            .ltout(n14578_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_100_LC_6_22_3.C_ON=1'b0;
    defparam i1_4_lut_adj_100_LC_6_22_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_100_LC_6_22_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_100_LC_6_22_3 (
            .in0(N__30452),
            .in1(N__32236),
            .in2(N__30429),
            .in3(N__30422),
            .lcout(),
            .ltout(n14582_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_102_LC_6_22_4.C_ON=1'b0;
    defparam i1_4_lut_adj_102_LC_6_22_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_102_LC_6_22_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_102_LC_6_22_4 (
            .in0(N__30404),
            .in1(N__30376),
            .in2(N__30360),
            .in3(N__30352),
            .lcout(),
            .ltout(n14588_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_104_LC_6_22_5.C_ON=1'b0;
    defparam i1_4_lut_adj_104_LC_6_22_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_104_LC_6_22_5.LUT_INIT=16'b1111111011111100;
    LogicCell40 i1_4_lut_adj_104_LC_6_22_5 (
            .in0(N__32076),
            .in1(N__30319),
            .in2(N__30303),
            .in3(N__30300),
            .lcout(n14592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13014_1_lut_LC_6_22_6.C_ON=1'b0;
    defparam i13014_1_lut_LC_6_22_6.SEQ_MODE=4'b0000;
    defparam i13014_1_lut_LC_6_22_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 i13014_1_lut_LC_6_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32637),
            .lcout(n15739),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_23_0.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41919),
            .in3(_gnd_net_),
            .lcout(n17_adj_638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12759_1_lut_LC_6_23_2.C_ON=1'b0;
    defparam i12759_1_lut_LC_6_23_2.SEQ_MODE=4'b0000;
    defparam i12759_1_lut_LC_6_23_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12759_1_lut_LC_6_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32390),
            .lcout(n15484),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_23_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36718),
            .lcout(n19_adj_640),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_6_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_6_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_6_23_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i14_3_lut_LC_6_23_4 (
            .in0(N__38661),
            .in1(N__46158),
            .in2(_gnd_net_),
            .in3(N__36569),
            .lcout(n306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_6_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_6_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_6_23_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i11_3_lut_LC_6_23_5 (
            .in0(N__46159),
            .in1(N__38754),
            .in2(_gnd_net_),
            .in3(N__40007),
            .lcout(n309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12762_4_lut_LC_6_24_0.C_ON=1'b0;
    defparam i12762_4_lut_LC_6_24_0.SEQ_MODE=4'b0000;
    defparam i12762_4_lut_LC_6_24_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12762_4_lut_LC_6_24_0 (
            .in0(N__35754),
            .in1(N__30528),
            .in2(N__31347),
            .in3(N__30603),
            .lcout(n12034),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_6_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_6_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_6_24_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2198_3_lut_LC_6_24_2 (
            .in0(_gnd_net_),
            .in1(N__35016),
            .in2(N__34992),
            .in3(N__34632),
            .lcout(),
            .ltout(n17_adj_710_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_117_LC_6_24_3.C_ON=1'b0;
    defparam i1_4_lut_adj_117_LC_6_24_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_117_LC_6_24_3.LUT_INIT=16'b1111110111111000;
    LogicCell40 i1_4_lut_adj_117_LC_6_24_3 (
            .in0(N__34633),
            .in1(N__35231),
            .in2(N__30543),
            .in3(N__35205),
            .lcout(n14236),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2197_3_lut_LC_6_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2197_3_lut_LC_6_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2197_3_lut_LC_6_24_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2197_3_lut_LC_6_24_4 (
            .in0(_gnd_net_),
            .in1(N__35481),
            .in2(N__35457),
            .in3(N__34634),
            .lcout(),
            .ltout(n19_adj_711_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_118_LC_6_24_5.C_ON=1'b0;
    defparam i1_4_lut_adj_118_LC_6_24_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_118_LC_6_24_5.LUT_INIT=16'b1111110111111000;
    LogicCell40 i1_4_lut_adj_118_LC_6_24_5 (
            .in0(N__34635),
            .in1(N__35435),
            .in2(N__30540),
            .in3(N__35415),
            .lcout(),
            .ltout(n14230_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_122_LC_6_24_6.C_ON=1'b0;
    defparam i1_4_lut_adj_122_LC_6_24_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_122_LC_6_24_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_122_LC_6_24_6 (
            .in0(N__30537),
            .in1(N__34254),
            .in2(N__30531),
            .in3(N__30615),
            .lcout(n14248),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2176_3_lut_LC_6_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2176_3_lut_LC_6_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2176_3_lut_LC_6_25_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i2176_3_lut_LC_6_25_0 (
            .in0(N__35820),
            .in1(N__35834),
            .in2(_gnd_net_),
            .in3(N__34656),
            .lcout(n61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_152_LC_6_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_152_LC_6_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_152_LC_6_25_1.LUT_INIT=16'b1111111111001010;
    LogicCell40 i1_4_lut_adj_152_LC_6_25_1 (
            .in0(N__35955),
            .in1(N__35969),
            .in2(N__34699),
            .in3(N__31296),
            .lcout(),
            .ltout(n14268_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_153_LC_6_25_2.C_ON=1'b0;
    defparam i1_4_lut_adj_153_LC_6_25_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_153_LC_6_25_2.LUT_INIT=16'b1111110011111010;
    LogicCell40 i1_4_lut_adj_153_LC_6_25_2 (
            .in0(N__35940),
            .in1(N__43006),
            .in2(N__30624),
            .in3(N__34655),
            .lcout(n14270),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_163_LC_6_25_3.C_ON=1'b0;
    defparam i1_4_lut_adj_163_LC_6_25_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_163_LC_6_25_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_163_LC_6_25_3 (
            .in0(N__35917),
            .in1(N__35968),
            .in2(N__43010),
            .in3(N__30726),
            .lcout(),
            .ltout(n14806_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12758_4_lut_LC_6_25_4.C_ON=1'b0;
    defparam i12758_4_lut_LC_6_25_4.SEQ_MODE=4'b0000;
    defparam i12758_4_lut_LC_6_25_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12758_4_lut_LC_6_25_4 (
            .in0(N__35875),
            .in1(N__35833),
            .in2(N__30621),
            .in3(N__35774),
            .lcout(n3237),
            .ltout(n3237_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_115_LC_6_25_5.C_ON=1'b0;
    defparam i1_4_lut_adj_115_LC_6_25_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_115_LC_6_25_5.LUT_INIT=16'b1111111110101100;
    LogicCell40 i1_4_lut_adj_115_LC_6_25_5 (
            .in0(N__35400),
            .in1(N__35376),
            .in2(N__30618),
            .in3(N__30774),
            .lcout(n14228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9894_4_lut_LC_6_25_6.C_ON=1'b0;
    defparam i9894_4_lut_LC_6_25_6.SEQ_MODE=4'b0000;
    defparam i9894_4_lut_LC_6_25_6.LUT_INIT=16'b1111101011101110;
    LogicCell40 i9894_4_lut_LC_6_25_6 (
            .in0(N__34565),
            .in1(N__35190),
            .in2(N__40563),
            .in3(N__34651),
            .lcout(n11861),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_154_LC_6_25_7.C_ON=1'b0;
    defparam i1_4_lut_adj_154_LC_6_25_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_154_LC_6_25_7.LUT_INIT=16'b1111111110101100;
    LogicCell40 i1_4_lut_adj_154_LC_6_25_7 (
            .in0(N__35918),
            .in1(N__35898),
            .in2(N__34700),
            .in3(N__30609),
            .lcout(n14272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_6_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_6_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_6_26_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2109_3_lut_LC_6_26_0 (
            .in0(N__30852),
            .in1(N__30597),
            .in2(N__43173),
            .in3(_gnd_net_),
            .lcout(n3205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_6_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_6_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_6_26_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2118_3_lut_LC_6_26_1 (
            .in0(_gnd_net_),
            .in1(N__31077),
            .in2(N__30588),
            .in3(N__43152),
            .lcout(n3214),
            .ltout(n3214_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_161_LC_6_26_2.C_ON=1'b0;
    defparam i1_4_lut_adj_161_LC_6_26_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_161_LC_6_26_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_161_LC_6_26_2 (
            .in0(N__35560),
            .in1(N__35618),
            .in2(N__30789),
            .in3(N__34389),
            .lcout(n14794),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_6_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_6_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_6_26_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2126_3_lut_LC_6_26_3 (
            .in0(_gnd_net_),
            .in1(N__37043),
            .in2(N__30786),
            .in3(N__43150),
            .lcout(n3222),
            .ltout(n3222_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_6_26_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_6_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_6_26_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i2193_3_lut_LC_6_26_4 (
            .in0(N__35310),
            .in1(_gnd_net_),
            .in2(N__30777),
            .in3(N__34629),
            .lcout(n27_adj_713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_6_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_6_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_6_26_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2119_3_lut_LC_6_26_5 (
            .in0(_gnd_net_),
            .in1(N__30768),
            .in2(N__30762),
            .in3(N__43151),
            .lcout(n3215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_162_LC_6_26_6.C_ON=1'b0;
    defparam i1_4_lut_adj_162_LC_6_26_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_162_LC_6_26_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_162_LC_6_26_6 (
            .in0(N__35524),
            .in1(N__36035),
            .in2(N__36013),
            .in3(N__30732),
            .lcout(n14800),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_6_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_6_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_6_27_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1923_3_lut_LC_6_27_0 (
            .in0(_gnd_net_),
            .in1(N__30720),
            .in2(N__30711),
            .in3(N__33696),
            .lcout(n2923),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_6_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_6_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_6_27_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2123_3_lut_LC_6_27_1 (
            .in0(_gnd_net_),
            .in1(N__30639),
            .in2(N__31457),
            .in3(N__43085),
            .lcout(n3219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_6_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_6_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_6_27_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2125_3_lut_LC_6_27_2 (
            .in0(_gnd_net_),
            .in1(N__30633),
            .in2(N__43147),
            .in3(N__31139),
            .lcout(n3221),
            .ltout(n3221_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_155_LC_6_27_3.C_ON=1'b0;
    defparam i1_2_lut_adj_155_LC_6_27_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_155_LC_6_27_3.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_155_LC_6_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30627),
            .in3(N__35221),
            .lcout(n14764),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_6_27_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_6_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_6_27_4.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2111_3_lut_LC_6_27_4 (
            .in0(N__31011),
            .in1(_gnd_net_),
            .in2(N__43149),
            .in3(N__30897),
            .lcout(n3207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_6_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_6_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_6_27_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2124_3_lut_LC_6_27_5 (
            .in0(_gnd_net_),
            .in1(N__31004),
            .in2(N__30972),
            .in3(N__43086),
            .lcout(n3220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_6_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_6_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_6_27_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2127_3_lut_LC_6_27_6 (
            .in0(_gnd_net_),
            .in1(N__30963),
            .in2(N__43148),
            .in3(N__30957),
            .lcout(n3223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_6_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_6_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_6_27_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2115_3_lut_LC_6_27_7 (
            .in0(_gnd_net_),
            .in1(N__34952),
            .in2(N__30930),
            .in3(N__43093),
            .lcout(n3211),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_36_LC_6_28_0.C_ON=1'b0;
    defparam i1_4_lut_adj_36_LC_6_28_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_36_LC_6_28_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_36_LC_6_28_0 (
            .in0(N__31202),
            .in1(N__34948),
            .in2(N__30920),
            .in3(N__31017),
            .lcout(),
            .ltout(n14216_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_37_LC_6_28_1.C_ON=1'b0;
    defparam i1_4_lut_adj_37_LC_6_28_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_37_LC_6_28_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_37_LC_6_28_1 (
            .in0(N__30892),
            .in1(N__34285),
            .in2(N__30876),
            .in3(N__43225),
            .lcout(),
            .ltout(n14222_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12724_4_lut_LC_6_28_2.C_ON=1'b0;
    defparam i12724_4_lut_LC_6_28_2.SEQ_MODE=4'b0000;
    defparam i12724_4_lut_LC_6_28_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12724_4_lut_LC_6_28_2 (
            .in0(N__30814),
            .in1(N__30872),
            .in2(N__30855),
            .in3(N__30847),
            .lcout(n3138),
            .ltout(n3138_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12720_1_lut_LC_6_28_3.C_ON=1'b0;
    defparam i12720_1_lut_LC_6_28_3.SEQ_MODE=4'b0000;
    defparam i12720_1_lut_LC_6_28_3.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12720_1_lut_LC_6_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30819),
            .in3(_gnd_net_),
            .lcout(n15445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_6_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_6_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_6_28_4.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2110_3_lut_LC_6_28_4 (
            .in0(N__30815),
            .in1(N__30795),
            .in2(N__43170),
            .in3(_gnd_net_),
            .lcout(n3206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_6_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_6_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_6_28_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i2137_3_lut_LC_6_28_5 (
            .in0(N__31230),
            .in1(N__40055),
            .in2(_gnd_net_),
            .in3(N__43133),
            .lcout(n3233),
            .ltout(n3233_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9958_4_lut_LC_6_28_6.C_ON=1'b0;
    defparam i9958_4_lut_LC_6_28_6.SEQ_MODE=4'b0000;
    defparam i9958_4_lut_LC_6_28_6.LUT_INIT=16'b1010000010001000;
    LogicCell40 i9958_4_lut_LC_6_28_6 (
            .in0(N__31215),
            .in1(N__35163),
            .in2(N__31206),
            .in3(N__34726),
            .lcout(n11926),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_6_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_6_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_6_28_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2114_3_lut_LC_6_28_7 (
            .in0(_gnd_net_),
            .in1(N__31203),
            .in2(N__31179),
            .in3(N__43134),
            .lcout(n3210),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_6_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_6_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_6_29_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2058_3_lut_LC_6_29_0 (
            .in0(_gnd_net_),
            .in1(N__31170),
            .in2(N__37218),
            .in3(N__31152),
            .lcout(n3122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_6_29_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_6_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_6_29_1.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2117_3_lut_LC_6_29_1 (
            .in0(N__31113),
            .in1(_gnd_net_),
            .in2(N__43172),
            .in3(N__31046),
            .lcout(n3213),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_6_29_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_6_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_6_29_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2135_3_lut_LC_6_29_2 (
            .in0(_gnd_net_),
            .in1(N__36898),
            .in2(N__31104),
            .in3(N__43138),
            .lcout(n3231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_6_29_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_6_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_6_29_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2134_3_lut_LC_6_29_3 (
            .in0(_gnd_net_),
            .in1(N__36787),
            .in2(N__43171),
            .in3(N__31089),
            .lcout(n3230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_35_LC_6_29_4.C_ON=1'b0;
    defparam i1_4_lut_adj_35_LC_6_29_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_35_LC_6_29_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_35_LC_6_29_4 (
            .in0(N__31072),
            .in1(N__31042),
            .in2(N__36768),
            .in3(N__31026),
            .lcout(n14210),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_6_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_6_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_6_29_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i2069_3_lut_LC_6_29_5 (
            .in0(N__31284),
            .in1(N__42224),
            .in2(_gnd_net_),
            .in3(N__37196),
            .lcout(n3133),
            .ltout(n3133_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_6_29_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_6_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_6_29_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2136_3_lut_LC_6_29_6 (
            .in0(_gnd_net_),
            .in1(N__31275),
            .in2(N__31263),
            .in3(N__43139),
            .lcout(n3232),
            .ltout(n3232_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10062_4_lut_LC_6_29_7.C_ON=1'b0;
    defparam i10062_4_lut_LC_6_29_7.SEQ_MODE=4'b0000;
    defparam i10062_4_lut_LC_6_29_7.LUT_INIT=16'b1111111111100000;
    LogicCell40 i10062_4_lut_LC_6_29_7 (
            .in0(N__40558),
            .in1(N__35174),
            .in2(N__31260),
            .in3(N__35125),
            .lcout(n12030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_119_LC_6_30_1.C_ON=1'b0;
    defparam i1_4_lut_adj_119_LC_6_30_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_119_LC_6_30_1.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_119_LC_6_30_1 (
            .in0(N__35739),
            .in1(N__35718),
            .in2(N__34578),
            .in3(N__34703),
            .lcout(n14234),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16_4_lut_LC_6_30_2.C_ON=1'b0;
    defparam i16_4_lut_LC_6_30_2.SEQ_MODE=4'b0000;
    defparam i16_4_lut_LC_6_30_2.LUT_INIT=16'b1010110000001100;
    LogicCell40 i16_4_lut_LC_6_30_2 (
            .in0(N__35127),
            .in1(N__35079),
            .in2(N__34728),
            .in3(N__35099),
            .lcout(n5_adj_703),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2188_3_lut_LC_6_30_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2188_3_lut_LC_6_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2188_3_lut_LC_6_30_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2188_3_lut_LC_6_30_3 (
            .in0(_gnd_net_),
            .in1(N__35679),
            .in2(N__35709),
            .in3(N__34702),
            .lcout(n37_adj_715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2194_3_lut_LC_6_30_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2194_3_lut_LC_6_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2194_3_lut_LC_6_30_4.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2194_3_lut_LC_6_30_4 (
            .in0(N__35358),
            .in1(N__35337),
            .in2(N__34727),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n25_adj_712_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_120_LC_6_30_5.C_ON=1'b0;
    defparam i1_4_lut_adj_120_LC_6_30_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_120_LC_6_30_5.LUT_INIT=16'b1111110011111010;
    LogicCell40 i1_4_lut_adj_120_LC_6_30_5 (
            .in0(N__35025),
            .in1(N__35046),
            .in2(N__31257),
            .in3(N__34707),
            .lcout(),
            .ltout(n14238_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_124_LC_6_30_6.C_ON=1'b0;
    defparam i1_4_lut_adj_124_LC_6_30_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_124_LC_6_30_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_124_LC_6_30_6 (
            .in0(N__31254),
            .in1(N__31248),
            .in2(N__31242),
            .in3(N__31239),
            .lcout(),
            .ltout(n14250_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_126_LC_6_30_7.C_ON=1'b0;
    defparam i1_4_lut_adj_126_LC_6_30_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_126_LC_6_30_7.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_126_LC_6_30_7 (
            .in0(N__35670),
            .in1(N__35643),
            .in2(N__31392),
            .in3(N__34708),
            .lcout(n14252),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_6_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_6_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_6_31_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2061_3_lut_LC_6_31_2 (
            .in0(_gnd_net_),
            .in1(N__31389),
            .in2(N__31362),
            .in3(N__37170),
            .lcout(n3125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2177_3_lut_LC_6_31_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2177_3_lut_LC_6_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2177_3_lut_LC_6_31_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2177_3_lut_LC_6_31_3 (
            .in0(_gnd_net_),
            .in1(N__35879),
            .in2(N__34730),
            .in3(N__35850),
            .lcout(n59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_132_LC_6_31_4.C_ON=1'b0;
    defparam i1_4_lut_adj_132_LC_6_31_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_132_LC_6_31_4.LUT_INIT=16'b1111111111100010;
    LogicCell40 i1_4_lut_adj_132_LC_6_31_4 (
            .in0(N__35607),
            .in1(N__34715),
            .in2(N__35634),
            .in3(N__31332),
            .lcout(),
            .ltout(n14254_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_133_LC_6_31_5.C_ON=1'b0;
    defparam i1_4_lut_adj_133_LC_6_31_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_133_LC_6_31_5.LUT_INIT=16'b1111110011111000;
    LogicCell40 i1_4_lut_adj_133_LC_6_31_5 (
            .in0(N__31305),
            .in1(N__31326),
            .in2(N__31320),
            .in3(N__31317),
            .lcout(),
            .ltout(n14256_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_134_LC_6_31_6.C_ON=1'b0;
    defparam i1_4_lut_adj_134_LC_6_31_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_134_LC_6_31_6.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_134_LC_6_31_6 (
            .in0(N__35597),
            .in1(N__35577),
            .in2(N__31308),
            .in3(N__34716),
            .lcout(n14258),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2203_3_lut_LC_6_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2203_3_lut_LC_6_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2203_3_lut_LC_6_31_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i2203_3_lut_LC_6_31_7 (
            .in0(N__35154),
            .in1(_gnd_net_),
            .in2(N__34729),
            .in3(N__35139),
            .lcout(n7_adj_708),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_150_LC_6_32_0.C_ON=1'b0;
    defparam i1_4_lut_adj_150_LC_6_32_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_150_LC_6_32_0.LUT_INIT=16'b1111111111001010;
    LogicCell40 i1_4_lut_adj_150_LC_6_32_0 (
            .in0(N__36024),
            .in1(N__36051),
            .in2(N__34731),
            .in3(N__31506),
            .lcout(),
            .ltout(n14264_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_151_LC_6_32_1.C_ON=1'b0;
    defparam i1_4_lut_adj_151_LC_6_32_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_151_LC_6_32_1.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_151_LC_6_32_1 (
            .in0(N__36014),
            .in1(N__35982),
            .in2(N__31299),
            .in3(N__34725),
            .lcout(n14266),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_136_LC_6_32_3.C_ON=1'b0;
    defparam i1_4_lut_adj_136_LC_6_32_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_136_LC_6_32_3.LUT_INIT=16'b1111111110111000;
    LogicCell40 i1_4_lut_adj_136_LC_6_32_3 (
            .in0(N__35568),
            .in1(N__34720),
            .in2(N__35538),
            .in3(N__31515),
            .lcout(),
            .ltout(n14260_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_144_LC_6_32_4.C_ON=1'b0;
    defparam i1_4_lut_adj_144_LC_6_32_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_144_LC_6_32_4.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_144_LC_6_32_4 (
            .in0(N__34721),
            .in1(N__35490),
            .in2(N__31509),
            .in3(N__35526),
            .lcout(n14262),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_6_32_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_6_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_6_32_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2056_3_lut_LC_6_32_6 (
            .in0(_gnd_net_),
            .in1(N__31500),
            .in2(N__31473),
            .in3(N__37157),
            .lcout(n3120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_7_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_7_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_7_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_2_lut_LC_7_17_0 (
            .in0(_gnd_net_),
            .in1(N__38402),
            .in2(_gnd_net_),
            .in3(N__31428),
            .lcout(n2101),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(n12625),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_7_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_7_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_7_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_3_lut_LC_7_17_1 (
            .in0(_gnd_net_),
            .in1(N__54399),
            .in2(N__38321),
            .in3(N__31425),
            .lcout(n2100),
            .ltout(),
            .carryin(n12625),
            .carryout(n12626),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_7_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_7_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_7_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_4_lut_LC_7_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38117),
            .in3(N__31416),
            .lcout(n2099),
            .ltout(),
            .carryin(n12626),
            .carryout(n12627),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_7_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_7_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_7_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_5_lut_LC_7_17_3 (
            .in0(_gnd_net_),
            .in1(N__54400),
            .in2(N__38427),
            .in3(N__31413),
            .lcout(n2098),
            .ltout(),
            .carryin(n12627),
            .carryout(n12628),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_7_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_7_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_7_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_6_lut_LC_7_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37973),
            .in3(N__31404),
            .lcout(n2097),
            .ltout(),
            .carryin(n12628),
            .carryout(n12629),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_7_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_7_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_7_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_7_lut_LC_7_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36173),
            .in3(N__31395),
            .lcout(n2096),
            .ltout(),
            .carryin(n12629),
            .carryout(n12630),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_7_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_7_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_7_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_8_lut_LC_7_17_6 (
            .in0(_gnd_net_),
            .in1(N__54402),
            .in2(N__38280),
            .in3(N__31572),
            .lcout(n2095),
            .ltout(),
            .carryin(n12630),
            .carryout(n12631),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_7_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_7_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_7_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_9_lut_LC_7_17_7 (
            .in0(_gnd_net_),
            .in1(N__54401),
            .in2(N__37676),
            .in3(N__31563),
            .lcout(n2094),
            .ltout(),
            .carryin(n12631),
            .carryout(n12632),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_7_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_7_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_7_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_10_lut_LC_7_18_0 (
            .in0(_gnd_net_),
            .in1(N__54389),
            .in2(N__36371),
            .in3(N__31554),
            .lcout(n2093),
            .ltout(),
            .carryin(bfn_7_18_0_),
            .carryout(n12633),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_7_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_7_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_7_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_11_lut_LC_7_18_1 (
            .in0(_gnd_net_),
            .in1(N__53560),
            .in2(N__36273),
            .in3(N__31551),
            .lcout(n2092),
            .ltout(),
            .carryin(n12633),
            .carryout(n12634),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_7_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_7_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_7_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_12_lut_LC_7_18_2 (
            .in0(_gnd_net_),
            .in1(N__54390),
            .in2(N__36207),
            .in3(N__31542),
            .lcout(n2091),
            .ltout(),
            .carryin(n12634),
            .carryout(n12635),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_7_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_7_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_7_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_13_lut_LC_7_18_3 (
            .in0(_gnd_net_),
            .in1(N__53561),
            .in2(N__36414),
            .in3(N__31539),
            .lcout(n2090),
            .ltout(),
            .carryin(n12635),
            .carryout(n12636),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_7_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_7_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_7_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_14_lut_LC_7_18_4 (
            .in0(_gnd_net_),
            .in1(N__54391),
            .in2(N__36242),
            .in3(N__31536),
            .lcout(n2089),
            .ltout(),
            .carryin(n12636),
            .carryout(n12637),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_7_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_7_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_7_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_15_lut_LC_7_18_5 (
            .in0(_gnd_net_),
            .in1(N__38024),
            .in2(N__54503),
            .in3(N__31527),
            .lcout(n2088),
            .ltout(),
            .carryin(n12637),
            .carryout(n12638),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_7_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_7_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_7_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_16_lut_LC_7_18_6 (
            .in0(_gnd_net_),
            .in1(N__54395),
            .in2(N__37887),
            .in3(N__31518),
            .lcout(n2087),
            .ltout(),
            .carryin(n12638),
            .carryout(n12639),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_7_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_7_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_7_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_17_lut_LC_7_18_7 (
            .in0(_gnd_net_),
            .in1(N__36464),
            .in2(N__54504),
            .in3(N__31725),
            .lcout(n2086),
            .ltout(),
            .carryin(n12639),
            .carryout(n12640),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_7_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_7_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_7_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_18_lut_LC_7_19_0 (
            .in0(_gnd_net_),
            .in1(N__31627),
            .in2(N__54459),
            .in3(N__31713),
            .lcout(n2085),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(n12641),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_7_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_7_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_7_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_19_lut_LC_7_19_1 (
            .in0(_gnd_net_),
            .in1(N__36318),
            .in2(N__54502),
            .in3(N__31704),
            .lcout(n2084),
            .ltout(),
            .carryin(n12641),
            .carryout(n12642),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_7_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_7_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_7_19_2.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1369_20_lut_LC_7_19_2 (
            .in0(N__54365),
            .in1(N__36093),
            .in2(N__34046),
            .in3(N__31701),
            .lcout(n2115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_7_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_7_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_7_19_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1383_3_lut_LC_7_19_3 (
            .in0(_gnd_net_),
            .in1(N__38279),
            .in2(N__34016),
            .in3(N__31680),
            .lcout(n2127),
            .ltout(n2127_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_94_LC_7_19_4.C_ON=1'b0;
    defparam i1_4_lut_adj_94_LC_7_19_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_94_LC_7_19_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_94_LC_7_19_4 (
            .in0(N__31663),
            .in1(N__31585),
            .in2(N__31647),
            .in3(N__31640),
            .lcout(n14384),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_7_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_7_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_7_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1306_3_lut_LC_7_19_5 (
            .in0(_gnd_net_),
            .in1(N__39717),
            .in2(N__36117),
            .in3(N__38210),
            .lcout(n2018),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_7_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_7_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_7_19_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1380_3_lut_LC_7_19_6 (
            .in0(_gnd_net_),
            .in1(N__36269),
            .in2(N__31608),
            .in3(N__33977),
            .lcout(n2124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12964_1_lut_LC_7_19_7.C_ON=1'b0;
    defparam i12964_1_lut_LC_7_19_7.SEQ_MODE=4'b0000;
    defparam i12964_1_lut_LC_7_19_7.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12964_1_lut_LC_7_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34017),
            .in3(_gnd_net_),
            .lcout(n15689),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_7_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_7_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_7_20_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1386_3_lut_LC_7_20_0 (
            .in0(N__38423),
            .in1(N__32007),
            .in2(N__34028),
            .in3(_gnd_net_),
            .lcout(n2130),
            .ltout(n2130_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_97_LC_7_20_1.C_ON=1'b0;
    defparam i1_4_lut_adj_97_LC_7_20_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_97_LC_7_20_1.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_97_LC_7_20_1 (
            .in0(N__31969),
            .in1(N__31940),
            .in2(N__31908),
            .in3(N__32190),
            .lcout(),
            .ltout(n13775_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_98_LC_7_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_98_LC_7_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_98_LC_7_20_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_98_LC_7_20_2 (
            .in0(N__31903),
            .in1(N__32053),
            .in2(N__31887),
            .in3(N__31767),
            .lcout(n14398),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_7_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_7_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_7_20_4.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1378_3_lut_LC_7_20_4 (
            .in0(N__34011),
            .in1(N__31878),
            .in2(N__36413),
            .in3(_gnd_net_),
            .lcout(n2122),
            .ltout(n2122_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_95_LC_7_20_5.C_ON=1'b0;
    defparam i1_3_lut_adj_95_LC_7_20_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_95_LC_7_20_5.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_95_LC_7_20_5 (
            .in0(_gnd_net_),
            .in1(N__31843),
            .in2(N__31827),
            .in3(N__31822),
            .lcout(),
            .ltout(n14386_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_96_LC_7_20_6.C_ON=1'b0;
    defparam i1_4_lut_adj_96_LC_7_20_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_96_LC_7_20_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_96_LC_7_20_6 (
            .in0(N__31792),
            .in1(N__31741),
            .in2(N__31776),
            .in3(N__31773),
            .lcout(n14392),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_7_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_7_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_7_20_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1377_3_lut_LC_7_20_7 (
            .in0(_gnd_net_),
            .in1(N__31761),
            .in2(N__36243),
            .in3(N__34010),
            .lcout(n2121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_7_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_7_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_7_21_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1450_3_lut_LC_7_21_0 (
            .in0(_gnd_net_),
            .in1(N__32285),
            .in2(N__32265),
            .in3(N__34144),
            .lcout(n2226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_7_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_7_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_7_21_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1389_3_lut_LC_7_21_1 (
            .in0(N__32223),
            .in1(N__38398),
            .in2(_gnd_net_),
            .in3(N__34019),
            .lcout(n2133),
            .ltout(n2133_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9925_3_lut_LC_7_21_2.C_ON=1'b0;
    defparam i9925_3_lut_LC_7_21_2.SEQ_MODE=4'b0000;
    defparam i9925_3_lut_LC_7_21_2.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9925_3_lut_LC_7_21_2 (
            .in0(_gnd_net_),
            .in1(N__32182),
            .in2(N__32193),
            .in3(N__32449),
            .lcout(n11892),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_7_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_7_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_7_21_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1457_3_lut_LC_7_21_5 (
            .in0(N__32183),
            .in1(_gnd_net_),
            .in2(N__34167),
            .in3(N__32157),
            .lcout(n2233),
            .ltout(n2233_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9982_4_lut_LC_7_21_6.C_ON=1'b0;
    defparam i9982_4_lut_LC_7_21_6.SEQ_MODE=4'b0000;
    defparam i9982_4_lut_LC_7_21_6.LUT_INIT=16'b1111111011001100;
    LogicCell40 i9982_4_lut_LC_7_21_6 (
            .in0(N__32023),
            .in1(N__32116),
            .in2(N__32100),
            .in3(N__32092),
            .lcout(n11950),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_7_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_7_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_7_21_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1374_3_lut_LC_7_21_7 (
            .in0(_gnd_net_),
            .in1(N__32070),
            .in2(N__36468),
            .in3(N__34020),
            .lcout(n2118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_7_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_7_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_7_22_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_7_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37847),
            .lcout(n24_adj_645),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_22_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_22_2 (
            .in0(N__36633),
            .in1(N__38727),
            .in2(_gnd_net_),
            .in3(N__46160),
            .lcout(n308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_7_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_7_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_7_22_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_7_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36632),
            .lcout(n22_adj_643),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_7_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_7_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_7_22_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1508_3_lut_LC_7_22_4 (
            .in0(_gnd_net_),
            .in1(N__32535),
            .in2(N__32526),
            .in3(N__32652),
            .lcout(n2316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_22_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_22_5 (
            .in0(N__46164),
            .in1(N__36537),
            .in2(_gnd_net_),
            .in3(N__38079),
            .lcout(n319),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_7_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_7_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_7_22_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1388_3_lut_LC_7_22_6 (
            .in0(_gnd_net_),
            .in1(N__32469),
            .in2(N__38322),
            .in3(N__34018),
            .lcout(n2132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_22_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_22_7 (
            .in0(N__36504),
            .in1(_gnd_net_),
            .in2(N__46195),
            .in3(N__38568),
            .lcout(n315),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i0_LC_7_23_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i0_LC_7_23_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i0_LC_7_23_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i0_LC_7_23_0 (
            .in0(N__32397),
            .in1(N__42115),
            .in2(N__32391),
            .in3(N__32376),
            .lcout(encoder0_position_scaled_0),
            .ltout(),
            .carryin(bfn_7_23_0_),
            .carryout(n12938),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i1_LC_7_23_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i1_LC_7_23_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i1_LC_7_23_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i1_LC_7_23_1 (
            .in0(N__35801),
            .in1(N__34701),
            .in2(N__42175),
            .in3(N__32373),
            .lcout(encoder0_position_scaled_1),
            .ltout(),
            .carryin(n12938),
            .carryout(n12939),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i2_LC_7_23_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i2_LC_7_23_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i2_LC_7_23_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i2_LC_7_23_2 (
            .in0(N__32370),
            .in1(N__43178),
            .in2(N__42178),
            .in3(N__32349),
            .lcout(encoder0_position_scaled_2),
            .ltout(),
            .carryin(n12939),
            .carryout(n12940),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i3_LC_7_23_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i3_LC_7_23_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i3_LC_7_23_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i3_LC_7_23_3 (
            .in0(N__32346),
            .in1(N__42128),
            .in2(N__37224),
            .in3(N__32319),
            .lcout(encoder0_position_scaled_3),
            .ltout(),
            .carryin(n12940),
            .carryout(n12941),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i4_LC_7_23_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i4_LC_7_23_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i4_LC_7_23_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i4_LC_7_23_4 (
            .in0(N__32316),
            .in1(N__33897),
            .in2(N__42179),
            .in3(N__33741),
            .lcout(encoder0_position_scaled_4),
            .ltout(),
            .carryin(n12941),
            .carryout(n12942),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i5_LC_7_23_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i5_LC_7_23_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i5_LC_7_23_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i5_LC_7_23_5 (
            .in0(N__33738),
            .in1(N__33714),
            .in2(N__42176),
            .in3(N__33555),
            .lcout(encoder0_position_scaled_5),
            .ltout(),
            .carryin(n12942),
            .carryout(n12943),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i6_LC_7_23_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i6_LC_7_23_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i6_LC_7_23_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i6_LC_7_23_6 (
            .in0(N__33552),
            .in1(N__33528),
            .in2(N__42180),
            .in3(N__33372),
            .lcout(encoder0_position_scaled_6),
            .ltout(),
            .carryin(n12943),
            .carryout(n12944),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i7_LC_7_23_7.C_ON=1'b1;
    defparam encoder0_position_scaled_i7_LC_7_23_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i7_LC_7_23_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i7_LC_7_23_7 (
            .in0(N__33369),
            .in1(N__33350),
            .in2(N__42177),
            .in3(N__33198),
            .lcout(encoder0_position_scaled_7),
            .ltout(),
            .carryin(n12944),
            .carryout(n12945),
            .clk(N__55778),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i8_LC_7_24_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i8_LC_7_24_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i8_LC_7_24_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i8_LC_7_24_0 (
            .in0(N__33195),
            .in1(N__33171),
            .in2(N__42185),
            .in3(N__33027),
            .lcout(encoder0_position_scaled_8),
            .ltout(),
            .carryin(bfn_7_24_0_),
            .carryout(n12946),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i9_LC_7_24_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i9_LC_7_24_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i9_LC_7_24_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i9_LC_7_24_1 (
            .in0(N__33020),
            .in1(N__32999),
            .in2(N__42181),
            .in3(N__32853),
            .lcout(encoder0_position_scaled_9),
            .ltout(),
            .carryin(n12946),
            .carryout(n12947),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i10_LC_7_24_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i10_LC_7_24_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i10_LC_7_24_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i10_LC_7_24_2 (
            .in0(N__32850),
            .in1(N__32829),
            .in2(N__42186),
            .in3(N__32706),
            .lcout(encoder0_position_scaled_10),
            .ltout(),
            .carryin(n12947),
            .carryout(n12948),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i11_LC_7_24_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i11_LC_7_24_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i11_LC_7_24_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i11_LC_7_24_3 (
            .in0(N__32703),
            .in1(N__32683),
            .in2(N__42182),
            .in3(N__32538),
            .lcout(encoder0_position_scaled_11),
            .ltout(),
            .carryin(n12948),
            .carryout(n12949),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i12_LC_7_24_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i12_LC_7_24_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i12_LC_7_24_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i12_LC_7_24_4 (
            .in0(N__34191),
            .in1(N__34170),
            .in2(N__42187),
            .in3(N__34053),
            .lcout(encoder0_position_scaled_12),
            .ltout(),
            .carryin(n12949),
            .carryout(n12950),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i13_LC_7_24_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i13_LC_7_24_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i13_LC_7_24_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i13_LC_7_24_5 (
            .in0(N__34050),
            .in1(N__34029),
            .in2(N__42183),
            .in3(N__33921),
            .lcout(encoder0_position_scaled_13),
            .ltout(),
            .carryin(n12950),
            .carryout(n12951),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i14_LC_7_24_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i14_LC_7_24_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i14_LC_7_24_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i14_LC_7_24_6 (
            .in0(N__37944),
            .in1(N__38217),
            .in2(N__42188),
            .in3(N__33918),
            .lcout(encoder0_position_scaled_14),
            .ltout(),
            .carryin(n12951),
            .carryout(n12952),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i15_LC_7_24_7.C_ON=1'b1;
    defparam encoder0_position_scaled_i15_LC_7_24_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i15_LC_7_24_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i15_LC_7_24_7 (
            .in0(N__39780),
            .in1(N__39888),
            .in2(N__42184),
            .in3(N__33915),
            .lcout(encoder0_position_scaled_15),
            .ltout(),
            .carryin(n12952),
            .carryout(n12953),
            .clk(N__55779),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i16_LC_7_25_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i16_LC_7_25_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i16_LC_7_25_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i16_LC_7_25_0 (
            .in0(N__44550),
            .in1(N__41805),
            .in2(N__42171),
            .in3(N__33912),
            .lcout(encoder0_position_scaled_16),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(n12954),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i17_LC_7_25_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i17_LC_7_25_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i17_LC_7_25_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i17_LC_7_25_1 (
            .in0(N__47988),
            .in1(N__50202),
            .in2(N__42189),
            .in3(N__33909),
            .lcout(encoder0_position_scaled_17),
            .ltout(),
            .carryin(n12954),
            .carryout(n12955),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i18_LC_7_25_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i18_LC_7_25_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i18_LC_7_25_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i18_LC_7_25_2 (
            .in0(N__45738),
            .in1(N__50676),
            .in2(N__42172),
            .in3(N__33906),
            .lcout(encoder0_position_scaled_18),
            .ltout(),
            .carryin(n12955),
            .carryout(n12956),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i19_LC_7_25_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i19_LC_7_25_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i19_LC_7_25_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i19_LC_7_25_3 (
            .in0(N__51324),
            .in1(N__51405),
            .in2(N__42190),
            .in3(N__33903),
            .lcout(encoder0_position_scaled_19),
            .ltout(),
            .carryin(n12956),
            .carryout(n12957),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i20_LC_7_25_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i20_LC_7_25_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i20_LC_7_25_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i20_LC_7_25_4 (
            .in0(N__48513),
            .in1(N__51300),
            .in2(N__42173),
            .in3(N__33900),
            .lcout(encoder0_position_scaled_20),
            .ltout(),
            .carryin(n12957),
            .carryout(n12958),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i21_LC_7_25_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i21_LC_7_25_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i21_LC_7_25_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i21_LC_7_25_5 (
            .in0(N__51531),
            .in1(N__51603),
            .in2(N__42191),
            .in3(N__34314),
            .lcout(encoder0_position_scaled_21),
            .ltout(),
            .carryin(n12958),
            .carryout(n12959),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i22_LC_7_25_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i22_LC_7_25_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i22_LC_7_25_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i22_LC_7_25_6 (
            .in0(N__52365),
            .in1(N__52275),
            .in2(N__42174),
            .in3(N__34311),
            .lcout(encoder0_position_scaled_22),
            .ltout(),
            .carryin(n12959),
            .carryout(n12960),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i23_LC_7_25_7.C_ON=1'b0;
    defparam encoder0_position_scaled_i23_LC_7_25_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i23_LC_7_25_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i23_LC_7_25_7 (
            .in0(N__46356),
            .in1(N__46425),
            .in2(N__42192),
            .in3(N__34308),
            .lcout(encoder0_position_scaled_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55783),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_7_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_7_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_7_26_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2113_3_lut_LC_7_26_0 (
            .in0(_gnd_net_),
            .in1(N__34305),
            .in2(N__43174),
            .in3(N__34293),
            .lcout(n3209),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2191_3_lut_LC_7_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2191_3_lut_LC_7_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2191_3_lut_LC_7_26_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2191_3_lut_LC_7_26_1 (
            .in0(N__35261),
            .in1(_gnd_net_),
            .in2(N__35247),
            .in3(N__34630),
            .lcout(),
            .ltout(n31_adj_714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_116_LC_7_26_2.C_ON=1'b0;
    defparam i1_4_lut_adj_116_LC_7_26_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_116_LC_7_26_2.LUT_INIT=16'b1111110111111000;
    LogicCell40 i1_4_lut_adj_116_LC_7_26_2 (
            .in0(N__34631),
            .in1(N__35291),
            .in2(N__34257),
            .in3(N__35277),
            .lcout(n14232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_7_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_7_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_7_26_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2129_3_lut_LC_7_26_3 (
            .in0(_gnd_net_),
            .in1(N__34244),
            .in2(N__34215),
            .in3(N__43156),
            .lcout(n3225),
            .ltout(n3225_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_156_LC_7_26_4.C_ON=1'b0;
    defparam i1_4_lut_adj_156_LC_7_26_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_156_LC_7_26_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_156_LC_7_26_4 (
            .in0(N__35008),
            .in1(N__35260),
            .in2(N__34203),
            .in3(N__35321),
            .lcout(),
            .ltout(n14776_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_158_LC_7_26_5.C_ON=1'b0;
    defparam i1_4_lut_adj_158_LC_7_26_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_158_LC_7_26_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_158_LC_7_26_5 (
            .in0(N__35470),
            .in1(N__35350),
            .in2(N__34200),
            .in3(N__34197),
            .lcout(),
            .ltout(n14780_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_159_LC_7_26_6.C_ON=1'b0;
    defparam i1_4_lut_adj_159_LC_7_26_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_159_LC_7_26_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_159_LC_7_26_6 (
            .in0(N__34410),
            .in1(N__35659),
            .in2(N__34548),
            .in3(N__35704),
            .lcout(n14786),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_7_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_7_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_7_27_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2131_3_lut_LC_7_27_0 (
            .in0(_gnd_net_),
            .in1(N__34544),
            .in2(N__34512),
            .in3(N__43125),
            .lcout(n3227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_7_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_7_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_7_27_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2120_3_lut_LC_7_27_1 (
            .in0(_gnd_net_),
            .in1(N__34497),
            .in2(N__43169),
            .in3(N__34467),
            .lcout(n3216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_7_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_7_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_7_27_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2122_3_lut_LC_7_27_2 (
            .in0(_gnd_net_),
            .in1(N__34458),
            .in2(N__34428),
            .in3(N__43129),
            .lcout(n3218),
            .ltout(n3218_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_157_LC_7_27_3.C_ON=1'b0;
    defparam i1_3_lut_adj_157_LC_7_27_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_157_LC_7_27_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_157_LC_7_27_3 (
            .in0(_gnd_net_),
            .in1(N__35392),
            .in2(N__34413),
            .in3(N__35041),
            .lcout(n14778),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_160_LC_7_27_4.C_ON=1'b0;
    defparam i1_4_lut_adj_160_LC_7_27_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_160_LC_7_27_4.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_160_LC_7_27_4 (
            .in0(N__35100),
            .in1(N__34404),
            .in2(N__35070),
            .in3(N__34395),
            .lcout(n14788),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_7_27_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_7_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_7_27_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_7_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34383),
            .lcout(n13_adj_570),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_7_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_7_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_7_27_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2130_3_lut_LC_7_27_7 (
            .in0(_gnd_net_),
            .in1(N__34374),
            .in2(N__43168),
            .in3(N__34362),
            .lcout(n3226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_7_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_7_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_7_28_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2048_3_lut_LC_7_28_0 (
            .in0(_gnd_net_),
            .in1(N__34338),
            .in2(N__34971),
            .in3(N__37216),
            .lcout(n3112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_7_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_7_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_7_28_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2128_3_lut_LC_7_28_1 (
            .in0(_gnd_net_),
            .in1(N__34932),
            .in2(N__43166),
            .in3(N__34916),
            .lcout(n3224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_7_28_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_7_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_7_28_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2132_3_lut_LC_7_28_2 (
            .in0(_gnd_net_),
            .in1(N__36874),
            .in2(N__34890),
            .in3(N__43117),
            .lcout(n3228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12725_1_lut_LC_7_28_3.C_ON=1'b0;
    defparam i12725_1_lut_LC_7_28_3.SEQ_MODE=4'b0000;
    defparam i12725_1_lut_LC_7_28_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12725_1_lut_LC_7_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34664),
            .lcout(n15450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i2_4_lut_LC_7_28_4 .C_ON=1'b0;
    defparam \debounce.i2_4_lut_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \debounce.i2_4_lut_LC_7_28_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \debounce.i2_4_lut_LC_7_28_4  (
            .in0(N__34875),
            .in1(N__39426),
            .in2(N__34853),
            .in3(N__34824),
            .lcout(\debounce.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_7_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_7_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_7_28_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2121_3_lut_LC_7_28_5 (
            .in0(_gnd_net_),
            .in1(N__34794),
            .in2(N__43167),
            .in3(N__34781),
            .lcout(n3217),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_7_28_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_7_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_7_28_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2133_3_lut_LC_7_28_6 (
            .in0(_gnd_net_),
            .in1(N__36837),
            .in2(N__34749),
            .in3(N__43124),
            .lcout(n3229),
            .ltout(n3229_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2200_3_lut_LC_7_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2200_3_lut_LC_7_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2200_3_lut_LC_7_28_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2200_3_lut_LC_7_28_7 (
            .in0(_gnd_net_),
            .in1(N__35055),
            .in2(N__34734),
            .in3(N__34663),
            .lcout(n13_adj_709),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_2_LC_7_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_2_LC_7_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_2_LC_7_29_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 encoder0_position_31__I_0_add_2173_2_LC_7_29_0 (
            .in0(_gnd_net_),
            .in1(N__34566),
            .in2(N__53636),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_29_0_),
            .carryout(n12907),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1 (
            .in0(_gnd_net_),
            .in1(N__40559),
            .in2(_gnd_net_),
            .in3(N__35178),
            .lcout(n3301),
            .ltout(),
            .carryin(n12907),
            .carryout(n12908),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2 (
            .in0(_gnd_net_),
            .in1(N__35175),
            .in2(N__53637),
            .in3(N__35157),
            .lcout(n3300),
            .ltout(),
            .carryin(n12908),
            .carryout(n12909),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3 (
            .in0(_gnd_net_),
            .in1(N__35150),
            .in2(_gnd_net_),
            .in3(N__35130),
            .lcout(n3299),
            .ltout(),
            .carryin(n12909),
            .carryout(n12910),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4 (
            .in0(_gnd_net_),
            .in1(N__35126),
            .in2(N__53638),
            .in3(N__35109),
            .lcout(n3298),
            .ltout(),
            .carryin(n12910),
            .carryout(n12911),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5 (
            .in0(N__35106),
            .in1(N__35098),
            .in2(_gnd_net_),
            .in3(N__35073),
            .lcout(n15097),
            .ltout(),
            .carryin(n12911),
            .carryout(n12912),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6 (
            .in0(_gnd_net_),
            .in1(N__35069),
            .in2(_gnd_net_),
            .in3(N__35049),
            .lcout(n3296),
            .ltout(),
            .carryin(n12912),
            .carryout(n12913),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7 (
            .in0(_gnd_net_),
            .in1(N__35042),
            .in2(N__53639),
            .in3(N__35019),
            .lcout(n3295),
            .ltout(),
            .carryin(n12913),
            .carryout(n12914),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0 (
            .in0(_gnd_net_),
            .in1(N__35015),
            .in2(N__53987),
            .in3(N__34974),
            .lcout(n3294),
            .ltout(),
            .carryin(bfn_7_30_0_),
            .carryout(n12915),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1 (
            .in0(_gnd_net_),
            .in1(N__35477),
            .in2(N__54002),
            .in3(N__35439),
            .lcout(n3293),
            .ltout(),
            .carryin(n12915),
            .carryout(n12916),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2 (
            .in0(_gnd_net_),
            .in1(N__35436),
            .in2(N__53988),
            .in3(N__35403),
            .lcout(n3292),
            .ltout(),
            .carryin(n12916),
            .carryout(n12917),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3 (
            .in0(_gnd_net_),
            .in1(N__35399),
            .in2(N__54003),
            .in3(N__35361),
            .lcout(n3291),
            .ltout(),
            .carryin(n12917),
            .carryout(n12918),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4 (
            .in0(_gnd_net_),
            .in1(N__35357),
            .in2(N__53989),
            .in3(N__35331),
            .lcout(n3290),
            .ltout(),
            .carryin(n12918),
            .carryout(n12919),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5 (
            .in0(_gnd_net_),
            .in1(N__35328),
            .in2(N__54004),
            .in3(N__35298),
            .lcout(n3289),
            .ltout(),
            .carryin(n12919),
            .carryout(n12920),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6 (
            .in0(_gnd_net_),
            .in1(N__53694),
            .in2(N__35295),
            .in3(N__35268),
            .lcout(n3288),
            .ltout(),
            .carryin(n12920),
            .carryout(n12921),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7 (
            .in0(_gnd_net_),
            .in1(N__35265),
            .in2(N__54005),
            .in3(N__35235),
            .lcout(n3287),
            .ltout(),
            .carryin(n12921),
            .carryout(n12922),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0 (
            .in0(_gnd_net_),
            .in1(N__35232),
            .in2(N__53990),
            .in3(N__35193),
            .lcout(n3286),
            .ltout(),
            .carryin(bfn_7_31_0_),
            .carryout(n12923),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1 (
            .in0(_gnd_net_),
            .in1(N__35735),
            .in2(N__53994),
            .in3(N__35712),
            .lcout(n3285),
            .ltout(),
            .carryin(n12923),
            .carryout(n12924),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2 (
            .in0(_gnd_net_),
            .in1(N__35705),
            .in2(N__53991),
            .in3(N__35673),
            .lcout(n3284),
            .ltout(),
            .carryin(n12924),
            .carryout(n12925),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3 (
            .in0(_gnd_net_),
            .in1(N__35666),
            .in2(N__53995),
            .in3(N__35637),
            .lcout(n3283),
            .ltout(),
            .carryin(n12925),
            .carryout(n12926),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4 (
            .in0(_gnd_net_),
            .in1(N__35630),
            .in2(N__53992),
            .in3(N__35601),
            .lcout(n3282),
            .ltout(),
            .carryin(n12926),
            .carryout(n12927),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5 (
            .in0(_gnd_net_),
            .in1(N__35598),
            .in2(N__53996),
            .in3(N__35571),
            .lcout(n3281),
            .ltout(),
            .carryin(n12927),
            .carryout(n12928),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6 (
            .in0(_gnd_net_),
            .in1(N__35567),
            .in2(N__53993),
            .in3(N__35529),
            .lcout(n3280),
            .ltout(),
            .carryin(n12928),
            .carryout(n12929),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7 (
            .in0(_gnd_net_),
            .in1(N__35525),
            .in2(N__53997),
            .in3(N__35484),
            .lcout(n3279),
            .ltout(),
            .carryin(n12929),
            .carryout(n12930),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0 (
            .in0(_gnd_net_),
            .in1(N__36047),
            .in2(N__53998),
            .in3(N__36018),
            .lcout(n3278),
            .ltout(),
            .carryin(bfn_7_32_0_),
            .carryout(n12931),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1 (
            .in0(_gnd_net_),
            .in1(N__36015),
            .in2(N__54006),
            .in3(N__35976),
            .lcout(n3277),
            .ltout(),
            .carryin(n12931),
            .carryout(n12932),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2 (
            .in0(_gnd_net_),
            .in1(N__35973),
            .in2(N__53999),
            .in3(N__35943),
            .lcout(n3276),
            .ltout(),
            .carryin(n12932),
            .carryout(n12933),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3 (
            .in0(_gnd_net_),
            .in1(N__43011),
            .in2(N__54007),
            .in3(N__35928),
            .lcout(n3275),
            .ltout(),
            .carryin(n12933),
            .carryout(n12934),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4 (
            .in0(_gnd_net_),
            .in1(N__35925),
            .in2(N__54000),
            .in3(N__35883),
            .lcout(n3274),
            .ltout(),
            .carryin(n12934),
            .carryout(n12935),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5 (
            .in0(_gnd_net_),
            .in1(N__35880),
            .in2(N__54008),
            .in3(N__35844),
            .lcout(n3273),
            .ltout(),
            .carryin(n12935),
            .carryout(n12936),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6 (
            .in0(_gnd_net_),
            .in1(N__35841),
            .in2(N__54001),
            .in3(N__35805),
            .lcout(n3272),
            .ltout(),
            .carryin(n12936),
            .carryout(n12937),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7 (
            .in0(N__53707),
            .in1(N__35802),
            .in2(N__35781),
            .in3(N__35757),
            .lcout(n14873),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_9_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_9_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_9_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_2_lut_LC_9_17_0 (
            .in0(_gnd_net_),
            .in1(N__38359),
            .in2(_gnd_net_),
            .in3(N__36078),
            .lcout(n2001),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(n12608),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_9_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_9_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_9_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_3_lut_LC_9_17_1 (
            .in0(_gnd_net_),
            .in1(N__38233),
            .in2(N__54360),
            .in3(N__36075),
            .lcout(n2000),
            .ltout(),
            .carryin(n12608),
            .carryout(n12609),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_9_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_9_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_4_lut_LC_9_17_2 (
            .in0(_gnd_net_),
            .in1(N__38456),
            .in2(_gnd_net_),
            .in3(N__36072),
            .lcout(n1999),
            .ltout(),
            .carryin(n12609),
            .carryout(n12610),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_9_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_9_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_9_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_5_lut_LC_9_17_3 (
            .in0(_gnd_net_),
            .in1(N__54201),
            .in2(N__39954),
            .in3(N__36069),
            .lcout(n1998),
            .ltout(),
            .carryin(n12610),
            .carryout(n12611),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_9_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_9_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_9_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_6_lut_LC_9_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39690),
            .in3(N__36066),
            .lcout(n1997),
            .ltout(),
            .carryin(n12611),
            .carryout(n12612),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_9_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_9_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_9_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_7_lut_LC_9_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39662),
            .in3(N__36063),
            .lcout(n1996),
            .ltout(),
            .carryin(n12612),
            .carryout(n12613),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_9_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_9_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_8_lut_LC_9_17_6 (
            .in0(_gnd_net_),
            .in1(N__54197),
            .in2(N__39618),
            .in3(N__36060),
            .lcout(n1995),
            .ltout(),
            .carryin(n12613),
            .carryout(n12614),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_9_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_9_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_9_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_9_lut_LC_9_17_7 (
            .in0(_gnd_net_),
            .in1(N__37787),
            .in2(N__54361),
            .in3(N__36057),
            .lcout(n1994),
            .ltout(),
            .carryin(n12614),
            .carryout(n12615),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_9_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_9_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_9_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_10_lut_LC_9_18_0 (
            .in0(_gnd_net_),
            .in1(N__53152),
            .in2(N__37748),
            .in3(N__36054),
            .lcout(n1993),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(n12616),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_9_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_9_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_9_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_11_lut_LC_9_18_1 (
            .in0(_gnd_net_),
            .in1(N__53158),
            .in2(N__37641),
            .in3(N__36135),
            .lcout(n1992),
            .ltout(),
            .carryin(n12616),
            .carryout(n12617),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_9_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_9_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_9_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_12_lut_LC_9_18_2 (
            .in0(_gnd_net_),
            .in1(N__53153),
            .in2(N__37721),
            .in3(N__36132),
            .lcout(n1991),
            .ltout(),
            .carryin(n12617),
            .carryout(n12618),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_9_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_9_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_9_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_13_lut_LC_9_18_3 (
            .in0(_gnd_net_),
            .in1(N__53159),
            .in2(N__37769),
            .in3(N__36129),
            .lcout(n1990),
            .ltout(),
            .carryin(n12618),
            .carryout(n12619),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_9_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_9_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_9_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_14_lut_LC_9_18_4 (
            .in0(_gnd_net_),
            .in1(N__53154),
            .in2(N__38052),
            .in3(N__36126),
            .lcout(n1989),
            .ltout(),
            .carryin(n12619),
            .carryout(n12620),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_9_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_9_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_9_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_15_lut_LC_9_18_5 (
            .in0(_gnd_net_),
            .in1(N__53160),
            .in2(N__37904),
            .in3(N__36123),
            .lcout(n1988),
            .ltout(),
            .carryin(n12620),
            .carryout(n12621),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_9_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_9_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_9_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_16_lut_LC_9_18_6 (
            .in0(_gnd_net_),
            .in1(N__39737),
            .in2(N__53559),
            .in3(N__36120),
            .lcout(n1987),
            .ltout(),
            .carryin(n12621),
            .carryout(n12622),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_9_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_9_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_9_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_17_lut_LC_9_18_7 (
            .in0(_gnd_net_),
            .in1(N__39716),
            .in2(N__53558),
            .in3(N__36102),
            .lcout(n1986),
            .ltout(),
            .carryin(n12622),
            .carryout(n12623),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_9_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_9_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_9_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_18_lut_LC_9_19_0 (
            .in0(_gnd_net_),
            .in1(N__53452),
            .in2(N__39926),
            .in3(N__36099),
            .lcout(n1985),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(n12624),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_9_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_9_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_9_19_1.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1302_19_lut_LC_9_19_1 (
            .in0(N__53453),
            .in1(N__37937),
            .in2(N__37926),
            .in3(N__36096),
            .lcout(n2016),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_9_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_9_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_9_19_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1313_3_lut_LC_9_19_2 (
            .in0(_gnd_net_),
            .in1(N__36336),
            .in2(N__37752),
            .in3(N__38184),
            .lcout(n2025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_9_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_9_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_9_19_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1310_3_lut_LC_9_19_3 (
            .in0(_gnd_net_),
            .in1(N__37770),
            .in2(N__38208),
            .in3(N__36330),
            .lcout(n2022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_9_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_9_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_9_19_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1305_3_lut_LC_9_19_4 (
            .in0(_gnd_net_),
            .in1(N__36324),
            .in2(N__39927),
            .in3(N__38195),
            .lcout(n2017),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_9_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_9_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_9_19_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1312_3_lut_LC_9_19_5 (
            .in0(_gnd_net_),
            .in1(N__37639),
            .in2(N__38207),
            .in3(N__36297),
            .lcout(n2024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_9_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_9_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_9_19_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1317_3_lut_LC_9_19_6 (
            .in0(_gnd_net_),
            .in1(N__39686),
            .in2(N__36291),
            .in3(N__38191),
            .lcout(n2029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_9_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_9_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_9_19_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1307_3_lut_LC_9_19_7 (
            .in0(_gnd_net_),
            .in1(N__36279),
            .in2(N__38209),
            .in3(N__39741),
            .lcout(n2019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_90_LC_9_20_0.C_ON=1'b0;
    defparam i1_4_lut_adj_90_LC_9_20_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_90_LC_9_20_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_90_LC_9_20_0 (
            .in0(N__36352),
            .in1(N__36259),
            .in2(N__38269),
            .in3(N__37663),
            .lcout(),
            .ltout(n14550_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_91_LC_9_20_1.C_ON=1'b0;
    defparam i1_4_lut_adj_91_LC_9_20_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_91_LC_9_20_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_91_LC_9_20_1 (
            .in0(N__36223),
            .in1(N__36199),
            .in2(N__36177),
            .in3(N__36397),
            .lcout(),
            .ltout(n14556_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_92_LC_9_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_92_LC_9_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_92_LC_9_20_2.LUT_INIT=16'b1111100011110000;
    LogicCell40 i1_4_lut_adj_92_LC_9_20_2 (
            .in0(N__36154),
            .in1(N__37966),
            .in2(N__36138),
            .in3(N__38367),
            .lcout(),
            .ltout(n14558_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_93_LC_9_20_3.C_ON=1'b0;
    defparam i1_4_lut_adj_93_LC_9_20_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_93_LC_9_20_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_93_LC_9_20_3 (
            .in0(N__37870),
            .in1(N__38011),
            .in2(N__36471),
            .in3(N__36451),
            .lcout(n14564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_9_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_9_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_9_20_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1311_3_lut_LC_9_20_4 (
            .in0(N__37722),
            .in1(_gnd_net_),
            .in2(N__38206),
            .in3(N__36423),
            .lcout(n2023),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_9_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_9_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_9_20_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1314_3_lut_LC_9_20_5 (
            .in0(_gnd_net_),
            .in1(N__36381),
            .in2(N__37797),
            .in3(N__38180),
            .lcout(n2026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_9_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_9_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_9_21_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_9_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42374),
            .lcout(n15_adj_636),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_9_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_9_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_9_21_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_9_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40579),
            .lcout(n32_adj_653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_21_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40072),
            .lcout(n31_adj_652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_21_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38977),
            .lcout(n28_adj_649),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_21_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36532),
            .lcout(n33_adj_654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44887),
            .lcout(n27_adj_648),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36499),
            .lcout(n29_adj_650),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40141),
            .lcout(n26_adj_647),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i0_LC_9_22_0 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i0_LC_9_22_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i0_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i0_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__36536),
            .in2(_gnd_net_),
            .in3(N__36516),
            .lcout(encoder0_position_0),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\quad_counter0.n13025 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i1_LC_9_22_1 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i1_LC_9_22_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i1_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i1_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__37367),
            .in2(N__40589),
            .in3(N__36513),
            .lcout(encoder0_position_1),
            .ltout(),
            .carryin(\quad_counter0.n13025 ),
            .carryout(\quad_counter0.n13026 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i2_LC_9_22_2 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i2_LC_9_22_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i2_LC_9_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i2_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__40076),
            .in2(N__37415),
            .in3(N__36510),
            .lcout(encoder0_position_2),
            .ltout(),
            .carryin(\quad_counter0.n13026 ),
            .carryout(\quad_counter0.n13027 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i3_LC_9_22_3 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i3_LC_9_22_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i3_LC_9_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i3_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__37371),
            .in2(N__42250),
            .in3(N__36507),
            .lcout(encoder0_position_3),
            .ltout(),
            .carryin(\quad_counter0.n13027 ),
            .carryout(\quad_counter0.n13028 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i4_LC_9_22_4 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i4_LC_9_22_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i4_LC_9_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i4_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__36503),
            .in2(N__37416),
            .in3(N__36483),
            .lcout(encoder0_position_4),
            .ltout(),
            .carryin(\quad_counter0.n13028 ),
            .carryout(\quad_counter0.n13029 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i5_LC_9_22_5 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i5_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i5_LC_9_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i5_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__37375),
            .in2(N__38987),
            .in3(N__36480),
            .lcout(encoder0_position_5),
            .ltout(),
            .carryin(\quad_counter0.n13029 ),
            .carryout(\quad_counter0.n13030 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i6_LC_9_22_6 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i6_LC_9_22_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i6_LC_9_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i6_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__44891),
            .in2(N__37417),
            .in3(N__36477),
            .lcout(encoder0_position_6),
            .ltout(),
            .carryin(\quad_counter0.n13030 ),
            .carryout(\quad_counter0.n13031 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i7_LC_9_22_7 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i7_LC_9_22_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i7_LC_9_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i7_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(N__37379),
            .in2(N__40151),
            .in3(N__36474),
            .lcout(encoder0_position_7),
            .ltout(),
            .carryin(\quad_counter0.n13031 ),
            .carryout(\quad_counter0.n13032 ),
            .clk(N__55780),
            .ce(N__39117),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i8_LC_9_23_0 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i8_LC_9_23_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i8_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i8_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__37380),
            .in2(N__36664),
            .in3(N__36642),
            .lcout(encoder0_position_8),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\quad_counter0.n13033 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i9_LC_9_23_1 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i9_LC_9_23_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i9_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i9_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__37840),
            .in2(N__37418),
            .in3(N__36639),
            .lcout(encoder0_position_9),
            .ltout(),
            .carryin(\quad_counter0.n13033 ),
            .carryout(\quad_counter0.n13034 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i10_LC_9_23_2 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i10_LC_9_23_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i10_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i10_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__37384),
            .in2(N__40008),
            .in3(N__36636),
            .lcout(encoder0_position_10),
            .ltout(),
            .carryin(\quad_counter0.n13034 ),
            .carryout(\quad_counter0.n13035 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i11_LC_9_23_3 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i11_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i11_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i11_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__36626),
            .in2(N__37419),
            .in3(N__36612),
            .lcout(encoder0_position_11),
            .ltout(),
            .carryin(\quad_counter0.n13035 ),
            .carryout(\quad_counter0.n13036 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i12_LC_9_23_4 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i12_LC_9_23_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i12_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i12_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__37388),
            .in2(N__36601),
            .in3(N__36573),
            .lcout(encoder0_position_12),
            .ltout(),
            .carryin(\quad_counter0.n13036 ),
            .carryout(\quad_counter0.n13037 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i13_LC_9_23_5 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i13_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i13_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i13_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__36565),
            .in2(N__37420),
            .in3(N__36546),
            .lcout(encoder0_position_13),
            .ltout(),
            .carryin(\quad_counter0.n13037 ),
            .carryout(\quad_counter0.n13038 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i14_LC_9_23_6 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i14_LC_9_23_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i14_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i14_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__37392),
            .in2(N__36720),
            .in3(N__36543),
            .lcout(encoder0_position_14),
            .ltout(),
            .carryin(\quad_counter0.n13038 ),
            .carryout(\quad_counter0.n13039 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i15_LC_9_23_7 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i15_LC_9_23_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i15_LC_9_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i15_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__42437),
            .in2(N__37421),
            .in3(N__36540),
            .lcout(encoder0_position_15),
            .ltout(),
            .carryin(\quad_counter0.n13039 ),
            .carryout(\quad_counter0.n13040 ),
            .clk(N__55784),
            .ce(N__39113),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i16_LC_9_24_0 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i16_LC_9_24_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i16_LC_9_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i16_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__41908),
            .in2(N__37422),
            .in3(N__36693),
            .lcout(encoder0_position_16),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\quad_counter0.n13041 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i17_LC_9_24_1 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i17_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i17_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i17_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__37399),
            .in2(N__42289),
            .in3(N__36690),
            .lcout(encoder0_position_17),
            .ltout(),
            .carryin(\quad_counter0.n13041 ),
            .carryout(\quad_counter0.n13042 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i18_LC_9_24_2 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i18_LC_9_24_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i18_LC_9_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i18_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__42373),
            .in2(N__37423),
            .in3(N__36687),
            .lcout(encoder0_position_18),
            .ltout(),
            .carryin(\quad_counter0.n13042 ),
            .carryout(\quad_counter0.n13043 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i19_LC_9_24_3 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i19_LC_9_24_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i19_LC_9_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i19_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__37403),
            .in2(N__45809),
            .in3(N__36684),
            .lcout(encoder0_position_19),
            .ltout(),
            .carryin(\quad_counter0.n13043 ),
            .carryout(\quad_counter0.n13044 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i20_LC_9_24_4 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i20_LC_9_24_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i20_LC_9_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i20_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(N__44605),
            .in2(N__37424),
            .in3(N__36681),
            .lcout(encoder0_position_20),
            .ltout(),
            .carryin(\quad_counter0.n13044 ),
            .carryout(\quad_counter0.n13045 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i21_LC_9_24_5 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i21_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i21_LC_9_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i21_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__37407),
            .in2(N__46331),
            .in3(N__36678),
            .lcout(encoder0_position_21),
            .ltout(),
            .carryin(\quad_counter0.n13045 ),
            .carryout(\quad_counter0.n13046 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i22_LC_9_24_6 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i22_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i22_LC_9_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i22_LC_9_24_6  (
            .in0(_gnd_net_),
            .in1(N__44798),
            .in2(N__37425),
            .in3(N__36675),
            .lcout(encoder0_position_22),
            .ltout(),
            .carryin(\quad_counter0.n13046 ),
            .carryout(\quad_counter0.n13047 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i23_LC_9_24_7 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i23_LC_9_24_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i23_LC_9_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i23_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__37411),
            .in2(N__41992),
            .in3(N__36672),
            .lcout(encoder0_position_23),
            .ltout(),
            .carryin(\quad_counter0.n13047 ),
            .carryout(\quad_counter0.n13048 ),
            .clk(N__55786),
            .ce(N__39111),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i24_LC_9_25_0 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i24_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i24_LC_9_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i24_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(N__37353),
            .in2(N__44728),
            .in3(N__36669),
            .lcout(encoder0_position_24),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\quad_counter0.n13049 ),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i25_LC_9_25_1 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i25_LC_9_25_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i25_LC_9_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i25_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__40355),
            .in2(N__37412),
            .in3(N__36753),
            .lcout(encoder0_position_25),
            .ltout(),
            .carryin(\quad_counter0.n13049 ),
            .carryout(\quad_counter0.n13050 ),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i26_LC_9_25_2 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i26_LC_9_25_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i26_LC_9_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i26_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__37357),
            .in2(N__42724),
            .in3(N__36750),
            .lcout(encoder0_position_26),
            .ltout(),
            .carryin(\quad_counter0.n13050 ),
            .carryout(\quad_counter0.n13051 ),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i27_LC_9_25_3 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i27_LC_9_25_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i27_LC_9_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i27_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(N__42813),
            .in2(N__37413),
            .in3(N__36747),
            .lcout(encoder0_position_27),
            .ltout(),
            .carryin(\quad_counter0.n13051 ),
            .carryout(\quad_counter0.n13052 ),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i28_LC_9_25_4 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i28_LC_9_25_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i28_LC_9_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i28_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__37361),
            .in2(N__40428),
            .in3(N__36744),
            .lcout(encoder0_position_28),
            .ltout(),
            .carryin(\quad_counter0.n13052 ),
            .carryout(\quad_counter0.n13053 ),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i29_LC_9_25_5 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i29_LC_9_25_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i29_LC_9_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i29_LC_9_25_5  (
            .in0(_gnd_net_),
            .in1(N__40735),
            .in2(N__37414),
            .in3(N__36741),
            .lcout(encoder0_position_29),
            .ltout(),
            .carryin(\quad_counter0.n13053 ),
            .carryout(\quad_counter0.n13054 ),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i30_LC_9_25_6 .C_ON=1'b1;
    defparam \quad_counter0.position_656__i30_LC_9_25_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i30_LC_9_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_656__i30_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__37365),
            .in2(N__40665),
            .in3(N__36738),
            .lcout(encoder0_position_30),
            .ltout(),
            .carryin(\quad_counter0.n13054 ),
            .carryout(\quad_counter0.n13055 ),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_656__i31_LC_9_25_7 .C_ON=1'b0;
    defparam \quad_counter0.position_656__i31_LC_9_25_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_656__i31_LC_9_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter0.position_656__i31_LC_9_25_7  (
            .in0(N__37366),
            .in1(N__46061),
            .in2(_gnd_net_),
            .in3(N__36735),
            .lcout(encoder0_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55787),
            .ce(N__39112),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_26_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_26_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36732),
            .lcout(n8_adj_575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_9_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_9_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_9_26_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_9_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44606),
            .lcout(n13_adj_634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_26_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_26_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_26_2 (
            .in0(N__38628),
            .in1(N__36719),
            .in2(_gnd_net_),
            .in3(N__46053),
            .lcout(n305),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i1_LC_9_26_3.C_ON=1'b0;
    defparam pwm_setpoint_i1_LC_9_26_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i1_LC_9_26_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i1_LC_9_26_3 (
            .in0(N__42932),
            .in1(N__55331),
            .in2(_gnd_net_),
            .in3(N__37530),
            .lcout(pwm_setpoint_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55789),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_9_26_5.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_9_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_9_26_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_9_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36969),
            .lcout(n21_adj_556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i0_LC_9_26_6.C_ON=1'b0;
    defparam pwm_setpoint_i0_LC_9_26_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i0_LC_9_26_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i0_LC_9_26_6 (
            .in0(N__55330),
            .in1(N__37440),
            .in2(_gnd_net_),
            .in3(N__42968),
            .lcout(pwm_setpoint_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55789),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_9_26_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_9_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_9_26_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_9_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36957),
            .lcout(n20_adj_557),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.debounce_cnt_50_LC_9_27_0 .C_ON=1'b0;
    defparam \quad_counter0.debounce_cnt_50_LC_9_27_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.debounce_cnt_50_LC_9_27_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \quad_counter0.debounce_cnt_50_LC_9_27_0  (
            .in0(N__39162),
            .in1(N__36992),
            .in2(N__39080),
            .in3(N__38927),
            .lcout(\quad_counter0.debounce_cnt ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55791),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_9_27_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_9_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_9_27_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_9_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36945),
            .lcout(n3_adj_580),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_new_i1_LC_9_27_2 .C_ON=1'b0;
    defparam \quad_counter0.a_new_i1_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_new_i1_LC_9_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.a_new_i1_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36993),
            .lcout(a_new_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55791),
            .ce(),
            .sr(_gnd_net_));
    defparam i9962_3_lut_LC_9_27_3.C_ON=1'b0;
    defparam i9962_3_lut_LC_9_27_3.SEQ_MODE=4'b0000;
    defparam i9962_3_lut_LC_9_27_3.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9962_3_lut_LC_9_27_3 (
            .in0(_gnd_net_),
            .in1(N__40056),
            .in2(N__36932),
            .in3(N__36905),
            .lcout(),
            .ltout(n11930_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_34_LC_9_27_4.C_ON=1'b0;
    defparam i1_4_lut_adj_34_LC_9_27_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_34_LC_9_27_4.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_34_LC_9_27_4 (
            .in0(N__36875),
            .in1(N__36835),
            .in2(N__36801),
            .in3(N__36794),
            .lcout(n13819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12559_4_lut_LC_9_27_5 .C_ON=1'b0;
    defparam \quad_counter0.i12559_4_lut_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12559_4_lut_LC_9_27_5 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \quad_counter0.i12559_4_lut_LC_9_27_5  (
            .in0(N__36991),
            .in1(N__39160),
            .in2(N__39081),
            .in3(N__38926),
            .lcout(\quad_counter0.a_prev_N_543 ),
            .ltout(\quad_counter0.a_prev_N_543_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_52_LC_9_27_6 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_52_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_prev_52_LC_9_27_6 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \quad_counter0.b_prev_52_LC_9_27_6  (
            .in0(N__39161),
            .in1(N__39045),
            .in2(N__37428),
            .in3(N__39135),
            .lcout(b_prev),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55791),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_9_27_7 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_9_27_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter0.b_prev_I_0_63_2_lut_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__39070),
            .in2(_gnd_net_),
            .in3(N__39042),
            .lcout(\quad_counter0.direction_N_536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_9_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_9_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_9_28_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2059_3_lut_LC_9_28_0 (
            .in0(_gnd_net_),
            .in1(N__37265),
            .in2(N__37239),
            .in3(N__37215),
            .lcout(n3123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i8_1_lut_LC_9_28_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i8_1_lut_LC_9_28_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i8_1_lut_LC_9_28_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i8_1_lut_LC_9_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43392),
            .lcout(n18_adj_598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_new_i0_LC_9_28_2 .C_ON=1'b0;
    defparam \quad_counter0.a_new_i0_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_new_i0_LC_9_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.a_new_i0_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37011),
            .lcout(\quad_counter0.a_new_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55793),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i3_1_lut_LC_9_28_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i3_1_lut_LC_9_28_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i3_1_lut_LC_9_28_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i3_1_lut_LC_9_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42896),
            .lcout(n23_adj_603),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i2_1_lut_LC_9_28_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i2_1_lut_LC_9_28_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i2_1_lut_LC_9_28_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i2_1_lut_LC_9_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42933),
            .lcout(n24_adj_604),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_9_28_5.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_9_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_9_28_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_9_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36981),
            .lcout(n4_adj_579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_9_28_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_9_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_9_28_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_9_28_6 (
            .in0(N__37461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n6_adj_577),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i1_1_lut_LC_9_28_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i1_1_lut_LC_9_28_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i1_1_lut_LC_9_28_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i1_1_lut_LC_9_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42969),
            .lcout(n25_adj_605),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i13_1_lut_LC_9_29_0.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i13_1_lut_LC_9_29_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i13_1_lut_LC_9_29_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i13_1_lut_LC_9_29_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44094),
            .lcout(n13_adj_593),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i20_1_lut_LC_9_29_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i20_1_lut_LC_9_29_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i20_1_lut_LC_9_29_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i20_1_lut_LC_9_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43907),
            .lcout(n6_adj_586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i9_1_lut_LC_9_29_2.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i9_1_lut_LC_9_29_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i9_1_lut_LC_9_29_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i9_1_lut_LC_9_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46908),
            .lcout(n17_adj_597),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i4_1_lut_LC_9_29_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i4_1_lut_LC_9_29_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i4_1_lut_LC_9_29_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i4_1_lut_LC_9_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43518),
            .lcout(n22_adj_602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i16_1_lut_LC_9_29_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i16_1_lut_LC_9_29_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i16_1_lut_LC_9_29_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i16_1_lut_LC_9_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43634),
            .lcout(n10_adj_590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i12_1_lut_LC_9_29_6.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i12_1_lut_LC_9_29_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i12_1_lut_LC_9_29_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i12_1_lut_LC_9_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44007),
            .lcout(n14_adj_594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_2_lut_LC_9_30_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_2_lut_LC_9_30_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_2_lut_LC_9_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_2_lut_LC_9_30_0 (
            .in0(_gnd_net_),
            .in1(N__37449),
            .in2(_gnd_net_),
            .in3(N__37431),
            .lcout(pwm_setpoint_23_N_171_0),
            .ltout(),
            .carryin(bfn_9_30_0_),
            .carryout(n12412),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_3_lut_LC_9_30_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_3_lut_LC_9_30_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_3_lut_LC_9_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_3_lut_LC_9_30_1 (
            .in0(_gnd_net_),
            .in1(N__37539),
            .in2(_gnd_net_),
            .in3(N__37521),
            .lcout(pwm_setpoint_23_N_171_1),
            .ltout(),
            .carryin(n12412),
            .carryout(n12413),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_4_lut_LC_9_30_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_4_lut_LC_9_30_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_4_lut_LC_9_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_4_lut_LC_9_30_2 (
            .in0(_gnd_net_),
            .in1(N__37518),
            .in2(_gnd_net_),
            .in3(N__37509),
            .lcout(pwm_setpoint_23_N_171_2),
            .ltout(),
            .carryin(n12413),
            .carryout(n12414),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_5_lut_LC_9_30_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_5_lut_LC_9_30_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_5_lut_LC_9_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_5_lut_LC_9_30_3 (
            .in0(_gnd_net_),
            .in1(N__37506),
            .in2(_gnd_net_),
            .in3(N__37500),
            .lcout(pwm_setpoint_23_N_171_3),
            .ltout(),
            .carryin(n12414),
            .carryout(n12415),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_6_lut_LC_9_30_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_6_lut_LC_9_30_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_6_lut_LC_9_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_6_lut_LC_9_30_4 (
            .in0(_gnd_net_),
            .in1(N__39303),
            .in2(_gnd_net_),
            .in3(N__37497),
            .lcout(pwm_setpoint_23_N_171_4),
            .ltout(),
            .carryin(n12415),
            .carryout(n12416),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_7_lut_LC_9_30_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_7_lut_LC_9_30_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_7_lut_LC_9_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_7_lut_LC_9_30_5 (
            .in0(_gnd_net_),
            .in1(N__39321),
            .in2(_gnd_net_),
            .in3(N__37494),
            .lcout(pwm_setpoint_23_N_171_5),
            .ltout(),
            .carryin(n12416),
            .carryout(n12417),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_8_lut_LC_9_30_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_8_lut_LC_9_30_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_8_lut_LC_9_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_8_lut_LC_9_30_6 (
            .in0(_gnd_net_),
            .in1(N__39468),
            .in2(_gnd_net_),
            .in3(N__37491),
            .lcout(pwm_setpoint_23_N_171_6),
            .ltout(),
            .carryin(n12417),
            .carryout(n12418),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_9_lut_LC_9_30_7.C_ON=1'b1;
    defparam unary_minus_13_add_3_9_lut_LC_9_30_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_9_lut_LC_9_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_9_lut_LC_9_30_7 (
            .in0(_gnd_net_),
            .in1(N__37488),
            .in2(_gnd_net_),
            .in3(N__37479),
            .lcout(pwm_setpoint_23_N_171_7),
            .ltout(),
            .carryin(n12418),
            .carryout(n12419),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_10_lut_LC_9_31_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_10_lut_LC_9_31_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_10_lut_LC_9_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_10_lut_LC_9_31_0 (
            .in0(_gnd_net_),
            .in1(N__37476),
            .in2(_gnd_net_),
            .in3(N__37467),
            .lcout(pwm_setpoint_23_N_171_8),
            .ltout(),
            .carryin(bfn_9_31_0_),
            .carryout(n12420),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_11_lut_LC_9_31_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_11_lut_LC_9_31_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_11_lut_LC_9_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_11_lut_LC_9_31_1 (
            .in0(_gnd_net_),
            .in1(N__39315),
            .in2(_gnd_net_),
            .in3(N__37464),
            .lcout(pwm_setpoint_23_N_171_9),
            .ltout(),
            .carryin(n12420),
            .carryout(n12421),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_12_lut_LC_9_31_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_12_lut_LC_9_31_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_12_lut_LC_9_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_12_lut_LC_9_31_2 (
            .in0(_gnd_net_),
            .in1(N__39309),
            .in2(_gnd_net_),
            .in3(N__37593),
            .lcout(pwm_setpoint_23_N_171_10),
            .ltout(),
            .carryin(n12421),
            .carryout(n12422),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_13_lut_LC_9_31_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_13_lut_LC_9_31_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_13_lut_LC_9_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_13_lut_LC_9_31_3 (
            .in0(_gnd_net_),
            .in1(N__37590),
            .in2(_gnd_net_),
            .in3(N__37581),
            .lcout(pwm_setpoint_23_N_171_11),
            .ltout(),
            .carryin(n12422),
            .carryout(n12423),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_14_lut_LC_9_31_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_14_lut_LC_9_31_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_14_lut_LC_9_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_14_lut_LC_9_31_4 (
            .in0(_gnd_net_),
            .in1(N__37578),
            .in2(_gnd_net_),
            .in3(N__37569),
            .lcout(pwm_setpoint_23_N_171_12),
            .ltout(),
            .carryin(n12423),
            .carryout(n12424),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_15_lut_LC_9_31_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_15_lut_LC_9_31_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_15_lut_LC_9_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_15_lut_LC_9_31_5 (
            .in0(_gnd_net_),
            .in1(N__39261),
            .in2(_gnd_net_),
            .in3(N__37566),
            .lcout(pwm_setpoint_23_N_171_13),
            .ltout(),
            .carryin(n12424),
            .carryout(n12425),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_16_lut_LC_9_31_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_16_lut_LC_9_31_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_16_lut_LC_9_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_16_lut_LC_9_31_6 (
            .in0(_gnd_net_),
            .in1(N__39582),
            .in2(_gnd_net_),
            .in3(N__37563),
            .lcout(pwm_setpoint_23_N_171_14),
            .ltout(),
            .carryin(n12425),
            .carryout(n12426),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_17_lut_LC_9_31_7.C_ON=1'b1;
    defparam unary_minus_13_add_3_17_lut_LC_9_31_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_17_lut_LC_9_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_17_lut_LC_9_31_7 (
            .in0(_gnd_net_),
            .in1(N__37560),
            .in2(_gnd_net_),
            .in3(N__37551),
            .lcout(pwm_setpoint_23_N_171_15),
            .ltout(),
            .carryin(n12426),
            .carryout(n12427),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_18_lut_LC_9_32_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_18_lut_LC_9_32_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_18_lut_LC_9_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_18_lut_LC_9_32_0 (
            .in0(_gnd_net_),
            .in1(N__39564),
            .in2(_gnd_net_),
            .in3(N__37548),
            .lcout(pwm_setpoint_23_N_171_16),
            .ltout(),
            .carryin(bfn_9_32_0_),
            .carryout(n12428),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_19_lut_LC_9_32_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_19_lut_LC_9_32_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_19_lut_LC_9_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_19_lut_LC_9_32_1 (
            .in0(_gnd_net_),
            .in1(N__41100),
            .in2(_gnd_net_),
            .in3(N__37545),
            .lcout(pwm_setpoint_23_N_171_17),
            .ltout(),
            .carryin(n12428),
            .carryout(n12429),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_20_lut_LC_9_32_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_20_lut_LC_9_32_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_20_lut_LC_9_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_20_lut_LC_9_32_2 (
            .in0(_gnd_net_),
            .in1(N__39438),
            .in2(_gnd_net_),
            .in3(N__37542),
            .lcout(pwm_setpoint_23_N_171_18),
            .ltout(),
            .carryin(n12429),
            .carryout(n12430),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_21_lut_LC_9_32_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_21_lut_LC_9_32_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_21_lut_LC_9_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_21_lut_LC_9_32_3 (
            .in0(_gnd_net_),
            .in1(N__37617),
            .in2(_gnd_net_),
            .in3(N__37608),
            .lcout(pwm_setpoint_23_N_171_19),
            .ltout(),
            .carryin(n12430),
            .carryout(n12431),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_22_lut_LC_9_32_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_22_lut_LC_9_32_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_22_lut_LC_9_32_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_22_lut_LC_9_32_4 (
            .in0(_gnd_net_),
            .in1(N__41091),
            .in2(_gnd_net_),
            .in3(N__37605),
            .lcout(pwm_setpoint_23_N_171_20),
            .ltout(),
            .carryin(n12431),
            .carryout(n12432),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_23_lut_LC_9_32_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_23_lut_LC_9_32_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_23_lut_LC_9_32_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_23_lut_LC_9_32_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44112),
            .in3(N__37602),
            .lcout(pwm_setpoint_23_N_171_21),
            .ltout(),
            .carryin(n12432),
            .carryout(n12433),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_24_lut_LC_9_32_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_24_lut_LC_9_32_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_24_lut_LC_9_32_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_24_lut_LC_9_32_6 (
            .in0(_gnd_net_),
            .in1(N__39570),
            .in2(_gnd_net_),
            .in3(N__37599),
            .lcout(pwm_setpoint_23_N_171_22),
            .ltout(),
            .carryin(n12433),
            .carryout(n12434),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i23_LC_9_32_7.C_ON=1'b0;
    defparam pwm_setpoint_i23_LC_9_32_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i23_LC_9_32_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 pwm_setpoint_i23_LC_9_32_7 (
            .in0(_gnd_net_),
            .in1(N__44339),
            .in2(_gnd_net_),
            .in3(N__37596),
            .lcout(pwm_setpoint_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55812),
            .ce(),
            .sr(N__44340));
    defparam i1_3_lut_adj_85_LC_10_17_0.C_ON=1'b0;
    defparam i1_3_lut_adj_85_LC_10_17_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_85_LC_10_17_0.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_85_LC_10_17_0 (
            .in0(_gnd_net_),
            .in1(N__39607),
            .in2(N__37640),
            .in3(N__37786),
            .lcout(n14408),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_10_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_10_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_10_17_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1246_3_lut_LC_10_17_1 (
            .in0(_gnd_net_),
            .in1(N__41226),
            .in2(N__41838),
            .in3(N__39839),
            .lcout(n1926),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_10_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_10_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_10_17_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1182_3_lut_LC_10_17_2 (
            .in0(_gnd_net_),
            .in1(N__44250),
            .in2(N__41803),
            .in3(N__45690),
            .lcout(n1830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_10_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_10_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_10_17_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1253_3_lut_LC_10_17_3 (
            .in0(N__41448),
            .in1(N__42423),
            .in2(_gnd_net_),
            .in3(N__39840),
            .lcout(n1933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_17_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_17_6 (
            .in0(N__38469),
            .in1(N__46181),
            .in2(_gnd_net_),
            .in3(N__37848),
            .lcout(n310),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_10_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_10_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_10_17_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1247_3_lut_LC_10_17_7 (
            .in0(_gnd_net_),
            .in1(N__41261),
            .in2(N__41241),
            .in3(N__39838),
            .lcout(n1927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_10_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_10_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_10_18_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1243_3_lut_LC_10_18_0 (
            .in0(_gnd_net_),
            .in1(N__41626),
            .in2(N__39874),
            .in3(N__41604),
            .lcout(n1923),
            .ltout(n1923_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_86_LC_10_18_1.C_ON=1'b0;
    defparam i1_3_lut_adj_86_LC_10_18_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_86_LC_10_18_1.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_86_LC_10_18_1 (
            .in0(_gnd_net_),
            .in1(N__37741),
            .in2(N__37725),
            .in3(N__37714),
            .lcout(n14410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_10_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_10_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_10_18_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1244_3_lut_LC_10_18_2 (
            .in0(_gnd_net_),
            .in1(N__41660),
            .in2(N__39873),
            .in3(N__41640),
            .lcout(n1924),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_10_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_10_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_10_18_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i1241_3_lut_LC_10_18_4 (
            .in0(N__39852),
            .in1(_gnd_net_),
            .in2(N__41523),
            .in3(N__41553),
            .lcout(n1921),
            .ltout(n1921_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_87_LC_10_18_5.C_ON=1'b0;
    defparam i1_4_lut_adj_87_LC_10_18_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_87_LC_10_18_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_87_LC_10_18_5 (
            .in0(N__38048),
            .in1(N__37698),
            .in2(N__37692),
            .in3(N__37689),
            .lcout(n14416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_10_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_10_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_10_18_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1315_3_lut_LC_10_18_6 (
            .in0(_gnd_net_),
            .in1(N__37683),
            .in2(N__39617),
            .in3(N__38173),
            .lcout(n2027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_10_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_10_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_10_18_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1245_3_lut_LC_10_18_7 (
            .in0(_gnd_net_),
            .in1(N__41676),
            .in2(N__41694),
            .in3(N__39845),
            .lcout(n1925),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_10_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_10_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_10_19_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1242_3_lut_LC_10_19_0 (
            .in0(_gnd_net_),
            .in1(N__41591),
            .in2(N__41571),
            .in3(N__39867),
            .lcout(n1922),
            .ltout(n1922_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_10_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_10_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_10_19_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1309_3_lut_LC_10_19_1 (
            .in0(_gnd_net_),
            .in1(N__38037),
            .in2(N__38031),
            .in3(N__38197),
            .lcout(n2021),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_89_LC_10_19_2.C_ON=1'b0;
    defparam i1_4_lut_adj_89_LC_10_19_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_89_LC_10_19_2.LUT_INIT=16'b1111111111101010;
    LogicCell40 i1_4_lut_adj_89_LC_10_19_2 (
            .in0(N__39730),
            .in1(N__37854),
            .in2(N__39630),
            .in3(N__37998),
            .lcout(),
            .ltout(n14420_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12944_4_lut_LC_10_19_3.C_ON=1'b0;
    defparam i12944_4_lut_LC_10_19_3.SEQ_MODE=4'b0000;
    defparam i12944_4_lut_LC_10_19_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12944_4_lut_LC_10_19_3 (
            .in0(N__39914),
            .in1(N__39703),
            .in2(N__37992),
            .in3(N__37922),
            .lcout(n1950),
            .ltout(n1950_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_10_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_10_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_10_19_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1318_3_lut_LC_10_19_4 (
            .in0(_gnd_net_),
            .in1(N__39950),
            .in2(N__37989),
            .in3(N__37986),
            .lcout(n2030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12941_1_lut_LC_10_19_5.C_ON=1'b0;
    defparam i12941_1_lut_LC_10_19_5.SEQ_MODE=4'b0000;
    defparam i12941_1_lut_LC_10_19_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12941_1_lut_LC_10_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38198),
            .lcout(n15666),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_10_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_10_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_10_19_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1237_3_lut_LC_10_19_6 (
            .in0(_gnd_net_),
            .in1(N__44523),
            .in2(N__41871),
            .in3(N__39868),
            .lcout(n1917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_10_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_10_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_10_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1308_3_lut_LC_10_19_7 (
            .in0(_gnd_net_),
            .in1(N__37911),
            .in2(N__37905),
            .in3(N__38196),
            .lcout(n2020),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9998_4_lut_LC_10_20_0.C_ON=1'b0;
    defparam i9998_4_lut_LC_10_20_0.SEQ_MODE=4'b0000;
    defparam i9998_4_lut_LC_10_20_0.LUT_INIT=16'b1111110011101100;
    LogicCell40 i9998_4_lut_LC_10_20_0 (
            .in0(N__38360),
            .in1(N__39946),
            .in2(N__38457),
            .in3(N__38234),
            .lcout(n11966),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_10_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_10_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_10_20_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1252_3_lut_LC_10_20_1 (
            .in0(_gnd_net_),
            .in1(N__41412),
            .in2(N__39884),
            .in3(N__41432),
            .lcout(n1932),
            .ltout(n1932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_10_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_10_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_10_20_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1319_3_lut_LC_10_20_2 (
            .in0(N__38179),
            .in1(_gnd_net_),
            .in2(N__38439),
            .in3(N__38436),
            .lcout(n2031),
            .ltout(n2031_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9996_4_lut_LC_10_20_3.C_ON=1'b0;
    defparam i9996_4_lut_LC_10_20_3.SEQ_MODE=4'b0000;
    defparam i9996_4_lut_LC_10_20_3.LUT_INIT=16'b1111110011111000;
    LogicCell40 i9996_4_lut_LC_10_20_3 (
            .in0(N__38403),
            .in1(N__38099),
            .in2(N__38370),
            .in3(N__38302),
            .lcout(n11964),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_10_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_10_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_10_20_4.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1321_3_lut_LC_10_20_4 (
            .in0(N__38361),
            .in1(N__38334),
            .in2(N__38205),
            .in3(_gnd_net_),
            .lcout(n2033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_10_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_10_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_10_20_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1316_3_lut_LC_10_20_5 (
            .in0(_gnd_net_),
            .in1(N__38289),
            .in2(N__39663),
            .in3(N__38178),
            .lcout(n2028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_10_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_10_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_10_20_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1320_3_lut_LC_10_20_7 (
            .in0(_gnd_net_),
            .in1(N__38250),
            .in2(N__38238),
            .in3(N__38174),
            .lcout(n2032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_10_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_10_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_10_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_10_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38088),
            .in3(N__38067),
            .lcout(n33),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(n12968),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_10_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_10_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_10_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_10_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38064),
            .in3(N__38055),
            .lcout(n32),
            .ltout(),
            .carryin(n12968),
            .carryout(n12969),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_10_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_10_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_10_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_10_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38592),
            .in3(N__38583),
            .lcout(n31),
            .ltout(),
            .carryin(n12969),
            .carryout(n12970),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_10_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_10_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_10_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_10_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40167),
            .in3(N__38580),
            .lcout(n30),
            .ltout(),
            .carryin(n12970),
            .carryout(n12971),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_10_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_10_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_10_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_10_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38577),
            .in3(N__38556),
            .lcout(n29),
            .ltout(),
            .carryin(n12971),
            .carryout(n12972),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_10_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_10_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_10_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_10_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38553),
            .in3(N__38544),
            .lcout(n28),
            .ltout(),
            .carryin(n12972),
            .carryout(n12973),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_10_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_10_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_10_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_10_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38541),
            .in3(N__38532),
            .lcout(n27),
            .ltout(),
            .carryin(n12973),
            .carryout(n12974),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_10_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_10_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_10_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_10_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38529),
            .in3(N__38520),
            .lcout(n26),
            .ltout(),
            .carryin(n12974),
            .carryout(n12975),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_10_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_10_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_10_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_10_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38517),
            .in3(N__38484),
            .lcout(n25_adj_551),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(n12976),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_10_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_10_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_10_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_10_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38481),
            .in3(N__38460),
            .lcout(n24),
            .ltout(),
            .carryin(n12976),
            .carryout(n12977),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_10_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_10_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_10_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_10_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39978),
            .in3(N__38739),
            .lcout(n23),
            .ltout(),
            .carryin(n12977),
            .carryout(n12978),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_10_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_10_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_10_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_10_22_3 (
            .in0(_gnd_net_),
            .in1(N__38736),
            .in2(_gnd_net_),
            .in3(N__38718),
            .lcout(n22),
            .ltout(),
            .carryin(n12978),
            .carryout(n12979),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_10_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_10_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_10_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_10_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38715),
            .in3(N__38682),
            .lcout(n21),
            .ltout(),
            .carryin(n12979),
            .carryout(n12980),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_10_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_10_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_10_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_10_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38679),
            .in3(N__38646),
            .lcout(n20),
            .ltout(),
            .carryin(n12980),
            .carryout(n12981),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_10_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_10_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_10_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_10_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38643),
            .in3(N__38616),
            .lcout(n19),
            .ltout(),
            .carryin(n12981),
            .carryout(n12982),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_10_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_10_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_10_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_10_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41946),
            .in3(N__38613),
            .lcout(n18),
            .ltout(),
            .carryin(n12982),
            .carryout(n12983),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_10_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_10_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_10_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_10_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38610),
            .in3(N__38598),
            .lcout(n17),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(n12984),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_10_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_10_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_10_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_10_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41709),
            .in3(N__38595),
            .lcout(n16),
            .ltout(),
            .carryin(n12984),
            .carryout(n12985),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_10_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_10_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_10_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_10_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38805),
            .in3(N__38793),
            .lcout(n15),
            .ltout(),
            .carryin(n12985),
            .carryout(n12986),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_10_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_10_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_10_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_10_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45789),
            .in3(N__38790),
            .lcout(n14),
            .ltout(),
            .carryin(n12986),
            .carryout(n12987),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_10_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_10_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_10_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_10_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38787),
            .in3(N__38775),
            .lcout(n13),
            .ltout(),
            .carryin(n12987),
            .carryout(n12988),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_10_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_10_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_10_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_10_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46305),
            .in3(N__38772),
            .lcout(n12),
            .ltout(),
            .carryin(n12988),
            .carryout(n12989),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_10_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_10_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_10_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_10_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44784),
            .in3(N__38769),
            .lcout(n11),
            .ltout(),
            .carryin(n12989),
            .carryout(n12990),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_10_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_10_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_10_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_10_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41961),
            .in3(N__38766),
            .lcout(n10),
            .ltout(),
            .carryin(n12990),
            .carryout(n12991),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_10_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_10_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_10_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_10_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44706),
            .in3(N__38763),
            .lcout(n9),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(n12992),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_10_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_10_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_10_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_10_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38823),
            .in3(N__38760),
            .lcout(n8),
            .ltout(),
            .carryin(n12992),
            .carryout(n12993),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_10_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_10_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_10_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_10_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38814),
            .in3(N__38757),
            .lcout(n7),
            .ltout(),
            .carryin(n12993),
            .carryout(n12994),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_10_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_10_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_10_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_10_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38832),
            .in3(N__38856),
            .lcout(n6),
            .ltout(),
            .carryin(n12994),
            .carryout(n12995),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_10_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_10_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_10_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_10_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38841),
            .in3(N__38853),
            .lcout(n5),
            .ltout(),
            .carryin(n12995),
            .carryout(n12996),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_10_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_10_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_10_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_10_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39018),
            .in3(N__38850),
            .lcout(n4),
            .ltout(),
            .carryin(n12996),
            .carryout(n12997),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_10_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_10_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_10_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_10_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39201),
            .in3(N__38847),
            .lcout(n3),
            .ltout(),
            .carryin(n12997),
            .carryout(n12998),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_10_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_10_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_10_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_10_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42102),
            .in3(N__38844),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40416),
            .lcout(n5_adj_626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_25_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_25_1.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42814),
            .in3(_gnd_net_),
            .lcout(n6_adj_627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_166_LC_10_25_2.C_ON=1'b0;
    defparam i1_3_lut_adj_166_LC_10_25_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_166_LC_10_25_2.LUT_INIT=16'b1010000000000000;
    LogicCell40 i1_3_lut_adj_166_LC_10_25_2 (
            .in0(N__46031),
            .in1(_gnd_net_),
            .in2(N__40689),
            .in3(N__40464),
            .lcout(n14574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40351),
            .lcout(n8_adj_629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_10_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_10_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_10_25_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_10_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42709),
            .lcout(n7_adj_628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_25_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_25_5 (
            .in0(_gnd_net_),
            .in1(N__46029),
            .in2(N__42815),
            .in3(N__42865),
            .lcout(n292),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_10_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_10_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_10_25_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_10_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40728),
            .lcout(n4_adj_625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_25_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_25_7 (
            .in0(_gnd_net_),
            .in1(N__46030),
            .in2(N__40663),
            .in3(N__40684),
            .lcout(n403),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i4_4_lut_LC_10_26_0.C_ON=1'b0;
    defparam LessThan_299_i4_4_lut_LC_10_26_0.SEQ_MODE=4'b0000;
    defparam LessThan_299_i4_4_lut_LC_10_26_0.LUT_INIT=16'b0100110101000100;
    LogicCell40 LessThan_299_i4_4_lut_LC_10_26_0 (
            .in0(N__45180),
            .in1(N__39009),
            .in2(N__45201),
            .in3(N__39003),
            .lcout(n4_adj_655),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_10_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_10_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_10_26_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i6_3_lut_LC_10_26_1 (
            .in0(N__38997),
            .in1(N__46060),
            .in2(_gnd_net_),
            .in3(N__38988),
            .lcout(n314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_new_i1_LC_10_26_2 .C_ON=1'b0;
    defparam \quad_counter0.b_new_i1_LC_10_26_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_new_i1_LC_10_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.b_new_i1_LC_10_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38928),
            .lcout(\quad_counter0.b_new_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55790),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_10_26_3.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_10_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_10_26_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_10_26_3 (
            .in0(N__38892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n25_adj_552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_10_26_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_10_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_10_26_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_10_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38880),
            .lcout(n10_adj_573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_10_26_5.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_10_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_10_26_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_10_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38868),
            .lcout(n12_adj_571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_10_26_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_10_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_10_26_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_10_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40653),
            .lcout(n3_adj_624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_10_26_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_10_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_10_26_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_10_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39189),
            .lcout(n23_adj_554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12508_3_lut_LC_10_27_0.C_ON=1'b0;
    defparam i12508_3_lut_LC_10_27_0.SEQ_MODE=4'b0000;
    defparam i12508_3_lut_LC_10_27_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12508_3_lut_LC_10_27_0 (
            .in0(N__43781),
            .in1(N__43762),
            .in2(_gnd_net_),
            .in3(N__39177),
            .lcout(n15233),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_prev_51_LC_10_27_1 .C_ON=1'b0;
    defparam \quad_counter0.a_prev_51_LC_10_27_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_prev_51_LC_10_27_1 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \quad_counter0.a_prev_51_LC_10_27_1  (
            .in0(N__39144),
            .in1(N__39134),
            .in2(N__39171),
            .in3(N__39076),
            .lcout(\quad_counter0.a_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55792),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_10_27_2 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_10_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter0.b_prev_I_0_65_2_lut_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(N__39159),
            .in2(_gnd_net_),
            .in3(N__39043),
            .lcout(),
            .ltout(\quad_counter0.direction_N_540_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_27_3 .C_ON=1'b0;
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_27_3 .LUT_INIT=16'b1100010011001000;
    LogicCell40 \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_27_3  (
            .in0(N__39143),
            .in1(N__39133),
            .in2(N__39120),
            .in3(N__39074),
            .lcout(direction_N_537),
            .ltout(direction_N_537_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.direction_57_LC_10_27_4 .C_ON=1'b0;
    defparam \quad_counter0.direction_57_LC_10_27_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.direction_57_LC_10_27_4 .LUT_INIT=16'b0101110010101100;
    LogicCell40 \quad_counter0.direction_57_LC_10_27_4  (
            .in0(N__39075),
            .in1(N__39024),
            .in2(N__39048),
            .in3(N__39044),
            .lcout(n1302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55792),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i29_2_lut_LC_10_27_6.C_ON=1'b0;
    defparam LessThan_299_i29_2_lut_LC_10_27_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i29_2_lut_LC_10_27_6.LUT_INIT=16'b0110011001100110;
    LogicCell40 LessThan_299_i29_2_lut_LC_10_27_6 (
            .in0(N__39212),
            .in1(N__46637),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n29_adj_672),
            .ltout(n29_adj_672_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12509_3_lut_LC_10_27_7.C_ON=1'b0;
    defparam i12509_3_lut_LC_10_27_7.SEQ_MODE=4'b0000;
    defparam i12509_3_lut_LC_10_27_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 i12509_3_lut_LC_10_27_7 (
            .in0(_gnd_net_),
            .in1(N__39213),
            .in2(N__39291),
            .in3(N__39288),
            .lcout(n15234),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12457_3_lut_LC_10_28_0.C_ON=1'b0;
    defparam i12457_3_lut_LC_10_28_0.SEQ_MODE=4'b0000;
    defparam i12457_3_lut_LC_10_28_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12457_3_lut_LC_10_28_0 (
            .in0(N__39399),
            .in1(N__39382),
            .in2(_gnd_net_),
            .in3(N__39282),
            .lcout(n15182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_10_28_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_10_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_10_28_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_10_28_2 (
            .in0(N__39276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n9_adj_574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i33_2_lut_LC_10_28_3.C_ON=1'b0;
    defparam LessThan_299_i33_2_lut_LC_10_28_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i33_2_lut_LC_10_28_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i33_2_lut_LC_10_28_3 (
            .in0(_gnd_net_),
            .in1(N__46593),
            .in2(_gnd_net_),
            .in3(N__40911),
            .lcout(n33_adj_675),
            .ltout(n33_adj_675_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12396_4_lut_LC_10_28_4.C_ON=1'b0;
    defparam i12396_4_lut_LC_10_28_4.SEQ_MODE=4'b0000;
    defparam i12396_4_lut_LC_10_28_4.LUT_INIT=16'b1111000011110001;
    LogicCell40 i12396_4_lut_LC_10_28_4 (
            .in0(N__39350),
            .in1(N__39383),
            .in2(N__39264),
            .in3(N__40782),
            .lcout(n15121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i14_1_lut_LC_10_28_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i14_1_lut_LC_10_28_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i14_1_lut_LC_10_28_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i14_1_lut_LC_10_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43701),
            .lcout(n12_adj_592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i16_LC_10_28_6.C_ON=1'b0;
    defparam pwm_setpoint_i16_LC_10_28_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i16_LC_10_28_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i16_LC_10_28_6 (
            .in0(N__43599),
            .in1(N__55307),
            .in2(_gnd_net_),
            .in3(N__39252),
            .lcout(pwm_setpoint_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55794),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i2_LC_10_28_7.C_ON=1'b0;
    defparam pwm_setpoint_i2_LC_10_28_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i2_LC_10_28_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 pwm_setpoint_i2_LC_10_28_7 (
            .in0(N__55306),
            .in1(_gnd_net_),
            .in2(N__39240),
            .in3(N__42897),
            .lcout(pwm_setpoint_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55794),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i14_LC_10_29_0.C_ON=1'b0;
    defparam pwm_setpoint_i14_LC_10_29_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i14_LC_10_29_0.LUT_INIT=16'b1111000010101010;
    LogicCell40 pwm_setpoint_i14_LC_10_29_0 (
            .in0(N__43674),
            .in1(_gnd_net_),
            .in2(N__39228),
            .in3(N__55329),
            .lcout(pwm_setpoint_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55797),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i10_3_lut_3_lut_LC_10_29_3.C_ON=1'b0;
    defparam LessThan_299_i10_3_lut_3_lut_LC_10_29_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i10_3_lut_3_lut_LC_10_29_3.LUT_INIT=16'b1000100011101110;
    LogicCell40 LessThan_299_i10_3_lut_3_lut_LC_10_29_3 (
            .in0(N__45306),
            .in1(N__45284),
            .in2(_gnd_net_),
            .in3(N__46713),
            .lcout(n10_adj_659),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12552_4_lut_LC_10_29_4.C_ON=1'b0;
    defparam i12552_4_lut_LC_10_29_4.SEQ_MODE=4'b0000;
    defparam i12552_4_lut_LC_10_29_4.LUT_INIT=16'b1111000111100000;
    LogicCell40 i12552_4_lut_LC_10_29_4 (
            .in0(N__39366),
            .in1(N__43821),
            .in2(N__39330),
            .in3(N__39360),
            .lcout(n15277),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12500_4_lut_LC_10_29_5.C_ON=1'b0;
    defparam i12500_4_lut_LC_10_29_5.SEQ_MODE=4'b0000;
    defparam i12500_4_lut_LC_10_29_5.LUT_INIT=16'b1111111011111111;
    LogicCell40 i12500_4_lut_LC_10_29_5 (
            .in0(N__39384),
            .in1(N__39354),
            .in2(N__43767),
            .in3(N__47379),
            .lcout(n15225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i30_3_lut_LC_10_29_6.C_ON=1'b0;
    defparam LessThan_299_i30_3_lut_LC_10_29_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i30_3_lut_LC_10_29_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 LessThan_299_i30_3_lut_LC_10_29_6 (
            .in0(N__43941),
            .in1(N__40929),
            .in2(_gnd_net_),
            .in3(N__43819),
            .lcout(),
            .ltout(n30_adj_673_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12542_4_lut_LC_10_29_7.C_ON=1'b0;
    defparam i12542_4_lut_LC_10_29_7.SEQ_MODE=4'b0000;
    defparam i12542_4_lut_LC_10_29_7.LUT_INIT=16'b1111000111100000;
    LogicCell40 i12542_4_lut_LC_10_29_7 (
            .in0(N__43820),
            .in1(N__40881),
            .in2(N__39339),
            .in3(N__39336),
            .lcout(n15267),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i6_1_lut_LC_10_30_0.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i6_1_lut_LC_10_30_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i6_1_lut_LC_10_30_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i6_1_lut_LC_10_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43448),
            .lcout(n20_adj_600),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i10_1_lut_LC_10_30_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i10_1_lut_LC_10_30_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i10_1_lut_LC_10_30_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i10_1_lut_LC_10_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43352),
            .lcout(n16_adj_596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i11_1_lut_LC_10_30_2.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i11_1_lut_LC_10_30_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i11_1_lut_LC_10_30_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i11_1_lut_LC_10_30_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43325),
            .lcout(n15_adj_595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i5_1_lut_LC_10_30_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i5_1_lut_LC_10_30_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i5_1_lut_LC_10_30_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i5_1_lut_LC_10_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43478),
            .lcout(n21_adj_601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i5_LC_10_30_4.C_ON=1'b0;
    defparam pwm_setpoint_i5_LC_10_30_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i5_LC_10_30_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i5_LC_10_30_4 (
            .in0(N__55323),
            .in1(N__39297),
            .in2(_gnd_net_),
            .in3(N__43449),
            .lcout(pwm_setpoint_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55801),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i7_1_lut_LC_10_30_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i7_1_lut_LC_10_30_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i7_1_lut_LC_10_30_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i7_1_lut_LC_10_30_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43421),
            .lcout(n19_adj_599),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i6_LC_10_30_6.C_ON=1'b0;
    defparam pwm_setpoint_i6_LC_10_30_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i6_LC_10_30_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 pwm_setpoint_i6_LC_10_30_6 (
            .in0(N__55324),
            .in1(_gnd_net_),
            .in2(N__43425),
            .in3(N__39462),
            .lcout(pwm_setpoint_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55801),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i10_LC_10_30_7.C_ON=1'b0;
    defparam pwm_setpoint_i10_LC_10_30_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i10_LC_10_30_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i10_LC_10_30_7 (
            .in0(N__43326),
            .in1(N__55325),
            .in2(_gnd_net_),
            .in3(N__39456),
            .lcout(pwm_setpoint_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55801),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i9_LC_10_31_0.C_ON=1'b0;
    defparam pwm_setpoint_i9_LC_10_31_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i9_LC_10_31_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i9_LC_10_31_0 (
            .in0(N__55326),
            .in1(N__39450),
            .in2(_gnd_net_),
            .in3(N__43353),
            .lcout(pwm_setpoint_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55806),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i4_LC_10_31_1.C_ON=1'b0;
    defparam pwm_setpoint_i4_LC_10_31_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i4_LC_10_31_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i4_LC_10_31_1 (
            .in0(N__43485),
            .in1(N__55328),
            .in2(_gnd_net_),
            .in3(N__39444),
            .lcout(pwm_setpoint_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55806),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i19_1_lut_LC_10_31_2.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i19_1_lut_LC_10_31_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i19_1_lut_LC_10_31_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i19_1_lut_LC_10_31_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43553),
            .lcout(n7_adj_587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i15_LC_10_31_3.C_ON=1'b0;
    defparam pwm_setpoint_i15_LC_10_31_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i15_LC_10_31_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i15_LC_10_31_3 (
            .in0(N__43635),
            .in1(N__55327),
            .in2(_gnd_net_),
            .in3(N__39432),
            .lcout(pwm_setpoint_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55806),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i1_LC_10_31_4 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i1_LC_10_31_4 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i1_LC_10_31_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \debounce.reg_out_i0_i1_LC_10_31_4  (
            .in0(N__47581),
            .in1(N__39425),
            .in2(_gnd_net_),
            .in3(N__39539),
            .lcout(h2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55806),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i31_2_lut_LC_10_31_6.C_ON=1'b0;
    defparam LessThan_299_i31_2_lut_LC_10_31_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i31_2_lut_LC_10_31_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i31_2_lut_LC_10_31_6 (
            .in0(_gnd_net_),
            .in1(N__39395),
            .in2(_gnd_net_),
            .in3(N__46454),
            .lcout(n31_adj_674),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i15_1_lut_LC_10_31_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i15_1_lut_LC_10_31_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i15_1_lut_LC_10_31_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i15_1_lut_LC_10_31_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43673),
            .lcout(n11_adj_591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i18_LC_10_32_0.C_ON=1'b0;
    defparam pwm_setpoint_i18_LC_10_32_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i18_LC_10_32_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i18_LC_10_32_0 (
            .in0(N__55332),
            .in1(N__43554),
            .in2(_gnd_net_),
            .in3(N__39576),
            .lcout(pwm_setpoint_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55813),
            .ce(),
            .sr(_gnd_net_));
    defparam i12212_4_lut_LC_10_32_1.C_ON=1'b0;
    defparam i12212_4_lut_LC_10_32_1.SEQ_MODE=4'b0000;
    defparam i12212_4_lut_LC_10_32_1.LUT_INIT=16'b1111110111100000;
    LogicCell40 i12212_4_lut_LC_10_32_1 (
            .in0(N__41181),
            .in1(N__41145),
            .in2(N__41205),
            .in3(N__41163),
            .lcout(n14937),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i23_1_lut_LC_10_32_2.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i23_1_lut_LC_10_32_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i23_1_lut_LC_10_32_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i23_1_lut_LC_10_32_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43847),
            .lcout(n3_adj_583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i17_1_lut_LC_10_32_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i17_1_lut_LC_10_32_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i17_1_lut_LC_10_32_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i17_1_lut_LC_10_32_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43598),
            .lcout(n9_adj_589),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i2_LC_10_32_4 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i2_LC_10_32_4 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i2_LC_10_32_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \debounce.reg_out_i0_i2_LC_10_32_4  (
            .in0(N__39558),
            .in1(N__39526),
            .in2(_gnd_net_),
            .in3(N__47621),
            .lcout(h1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55813),
            .ce(),
            .sr(_gnd_net_));
    defparam i12211_4_lut_LC_10_32_5.C_ON=1'b0;
    defparam i12211_4_lut_LC_10_32_5.SEQ_MODE=4'b0000;
    defparam i12211_4_lut_LC_10_32_5.LUT_INIT=16'b1011001010110000;
    LogicCell40 i12211_4_lut_LC_10_32_5 (
            .in0(N__41180),
            .in1(N__41144),
            .in2(N__41204),
            .in3(N__41162),
            .lcout(),
            .ltout(n14936_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12213_3_lut_LC_10_32_6.C_ON=1'b0;
    defparam i12213_3_lut_LC_10_32_6.SEQ_MODE=4'b0000;
    defparam i12213_3_lut_LC_10_32_6.LUT_INIT=16'b0101010100001111;
    LogicCell40 i12213_3_lut_LC_10_32_6 (
            .in0(N__39498),
            .in1(_gnd_net_),
            .in2(N__39492),
            .in3(N__41124),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i22_LC_10_32_7.C_ON=1'b0;
    defparam pwm_setpoint_i22_LC_10_32_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i22_LC_10_32_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i22_LC_10_32_7 (
            .in0(N__43848),
            .in1(N__55333),
            .in2(_gnd_net_),
            .in3(N__39474),
            .lcout(pwm_setpoint_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55813),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_11_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_11_17_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1181_3_lut_LC_11_17_0 (
            .in0(_gnd_net_),
            .in1(N__44238),
            .in2(N__41804),
            .in3(N__45535),
            .lcout(n1829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12513_3_lut_LC_11_17_1.C_ON=1'b0;
    defparam i12513_3_lut_LC_11_17_1.SEQ_MODE=4'b0000;
    defparam i12513_3_lut_LC_11_17_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12513_3_lut_LC_11_17_1 (
            .in0(_gnd_net_),
            .in1(N__49790),
            .in2(N__44466),
            .in3(N__41796),
            .lcout(n1826),
            .ltout(n1826_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_81_LC_11_17_2.C_ON=1'b0;
    defparam i1_4_lut_adj_81_LC_11_17_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_81_LC_11_17_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_81_LC_11_17_2 (
            .in0(N__41827),
            .in1(N__41257),
            .in2(N__39621),
            .in3(N__41656),
            .lcout(n14526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_11_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_11_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_11_17_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1248_3_lut_LC_11_17_3 (
            .in0(_gnd_net_),
            .in1(N__41291),
            .in2(N__41274),
            .in3(N__39841),
            .lcout(n1928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_82_LC_11_17_4.C_ON=1'b0;
    defparam i1_3_lut_adj_82_LC_11_17_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_82_LC_11_17_4.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_82_LC_11_17_4 (
            .in0(_gnd_net_),
            .in1(N__41587),
            .in2(N__41627),
            .in3(N__39591),
            .lcout(),
            .ltout(n14530_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_83_LC_11_17_5.C_ON=1'b0;
    defparam i1_4_lut_adj_83_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_83_LC_11_17_5.LUT_INIT=16'b1111100011110000;
    LogicCell40 i1_4_lut_adj_83_LC_11_17_5 (
            .in0(N__41320),
            .in1(N__41290),
            .in2(N__39585),
            .in3(N__39762),
            .lcout(n14532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_11_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_11_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_11_17_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1249_3_lut_LC_11_17_6 (
            .in0(_gnd_net_),
            .in1(N__41321),
            .in2(N__39872),
            .in3(N__41301),
            .lcout(n1929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_79_LC_11_18_0.C_ON=1'b0;
    defparam i1_2_lut_adj_79_LC_11_18_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_79_LC_11_18_0.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_79_LC_11_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45495),
            .in3(N__45537),
            .lcout(n14520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_11_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_11_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_11_18_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1180_3_lut_LC_11_18_1 (
            .in0(_gnd_net_),
            .in1(N__45493),
            .in2(N__44226),
            .in3(N__41760),
            .lcout(n1828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_11_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_11_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_11_18_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1175_3_lut_LC_11_18_2 (
            .in0(_gnd_net_),
            .in1(N__44424),
            .in2(N__41790),
            .in3(N__50313),
            .lcout(n1823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_11_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_11_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_11_18_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1176_3_lut_LC_11_18_3 (
            .in0(_gnd_net_),
            .in1(N__50286),
            .in2(N__44439),
            .in3(N__41767),
            .lcout(n1824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12443_3_lut_LC_11_18_4.C_ON=1'b0;
    defparam i12443_3_lut_LC_11_18_4.SEQ_MODE=4'b0000;
    defparam i12443_3_lut_LC_11_18_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 i12443_3_lut_LC_11_18_4 (
            .in0(_gnd_net_),
            .in1(N__50343),
            .in2(N__41789),
            .in3(N__44451),
            .lcout(n1825),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_11_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_11_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_11_18_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1171_3_lut_LC_11_18_5 (
            .in0(_gnd_net_),
            .in1(N__44562),
            .in2(N__44583),
            .in3(N__41768),
            .lcout(n1819),
            .ltout(n1819_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12922_4_lut_LC_11_18_6.C_ON=1'b0;
    defparam i12922_4_lut_LC_11_18_6.SEQ_MODE=4'b0000;
    defparam i12922_4_lut_LC_11_18_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12922_4_lut_LC_11_18_6 (
            .in0(N__40176),
            .in1(N__44519),
            .in2(N__39753),
            .in3(N__39750),
            .lcout(n1851),
            .ltout(n1851_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_11_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_11_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_11_18_7.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1240_3_lut_LC_11_18_7 (
            .in0(N__41856),
            .in1(N__41508),
            .in2(N__39744),
            .in3(_gnd_net_),
            .lcout(n1920),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_11_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_11_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_11_19_0.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1239_3_lut_LC_11_19_0 (
            .in0(N__41495),
            .in1(_gnd_net_),
            .in2(N__39882),
            .in3(N__41481),
            .lcout(n1919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_11_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_11_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_11_19_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1250_3_lut_LC_11_19_1 (
            .in0(N__41337),
            .in1(_gnd_net_),
            .in2(N__41363),
            .in3(N__39860),
            .lcout(n1930),
            .ltout(n1930_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_88_LC_11_19_2.C_ON=1'b0;
    defparam i1_2_lut_adj_88_LC_11_19_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_88_LC_11_19_2.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_88_LC_11_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39666),
            .in3(N__39652),
            .lcout(n14540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_11_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_11_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_11_19_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1251_3_lut_LC_11_19_3 (
            .in0(_gnd_net_),
            .in1(N__41376),
            .in2(N__41396),
            .in3(N__39859),
            .lcout(n1931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_11_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_11_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_11_19_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1238_3_lut_LC_11_19_4 (
            .in0(_gnd_net_),
            .in1(N__41471),
            .in2(N__39881),
            .in3(N__41457),
            .lcout(n1918),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_80_LC_11_19_5.C_ON=1'b0;
    defparam i1_4_lut_adj_80_LC_11_19_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_80_LC_11_19_5.LUT_INIT=16'b1111111111101010;
    LogicCell40 i1_4_lut_adj_80_LC_11_19_5 (
            .in0(N__44393),
            .in1(N__45609),
            .in2(N__39903),
            .in3(N__50223),
            .lcout(),
            .ltout(n14176_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12901_4_lut_LC_11_19_6.C_ON=1'b0;
    defparam i12901_4_lut_LC_11_19_6.SEQ_MODE=4'b0000;
    defparam i12901_4_lut_LC_11_19_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12901_4_lut_LC_11_19_6 (
            .in0(N__44371),
            .in1(N__44578),
            .in2(N__39894),
            .in3(N__47942),
            .lcout(n1752),
            .ltout(n1752_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_11_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_11_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_11_19_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1183_3_lut_LC_11_19_7 (
            .in0(_gnd_net_),
            .in1(N__44265),
            .in2(N__39891),
            .in3(N__45597),
            .lcout(n1831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12919_1_lut_LC_11_20_0.C_ON=1'b0;
    defparam i12919_1_lut_LC_11_20_0.SEQ_MODE=4'b0000;
    defparam i12919_1_lut_LC_11_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12919_1_lut_LC_11_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39883),
            .lcout(n15644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_11_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_11_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_11_20_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1184_3_lut_LC_11_20_2 (
            .in0(_gnd_net_),
            .in1(N__45669),
            .in2(N__44283),
            .in3(N__41770),
            .lcout(n1832),
            .ltout(n1832_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10000_4_lut_LC_11_20_3.C_ON=1'b0;
    defparam i10000_4_lut_LC_11_20_3.SEQ_MODE=4'b0000;
    defparam i10000_4_lut_LC_11_20_3.LUT_INIT=16'b1111101011101010;
    LogicCell40 i10000_4_lut_LC_11_20_3 (
            .in0(N__41353),
            .in1(N__42406),
            .in2(N__39765),
            .in3(N__41431),
            .lcout(n11968),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_11_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_11_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_11_20_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1185_3_lut_LC_11_20_4 (
            .in0(N__44301),
            .in1(N__45634),
            .in2(_gnd_net_),
            .in3(N__41769),
            .lcout(n1833),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_11_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_11_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_11_20_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1172_3_lut_LC_11_20_5 (
            .in0(N__44373),
            .in1(_gnd_net_),
            .in2(N__41792),
            .in3(N__44355),
            .lcout(n1820),
            .ltout(n1820_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_84_LC_11_20_6.C_ON=1'b0;
    defparam i1_3_lut_adj_84_LC_11_20_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_84_LC_11_20_6.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_84_LC_11_20_6 (
            .in0(_gnd_net_),
            .in1(N__41539),
            .in2(N__40179),
            .in3(N__41854),
            .lcout(n14538),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_11_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_11_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_11_20_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1174_3_lut_LC_11_20_7 (
            .in0(_gnd_net_),
            .in1(N__44412),
            .in2(N__41791),
            .in3(N__50253),
            .lcout(n1822),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_11_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_11_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_11_21_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_11_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42251),
            .lcout(n30_adj_651),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_11_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_11_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_11_21_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i8_3_lut_LC_11_21_2 (
            .in0(N__40158),
            .in1(N__46192),
            .in2(_gnd_net_),
            .in3(N__40152),
            .lcout(n312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_11_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_11_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_11_21_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i3_3_lut_LC_11_21_3 (
            .in0(N__46193),
            .in1(N__40086),
            .in2(_gnd_net_),
            .in3(N__40080),
            .lcout(n317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_11_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_11_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_11_21_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_11_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40006),
            .lcout(n23_adj_644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_11_21_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_11_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_11_21_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_11_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39969),
            .lcout(n24_adj_553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_11_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_11_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_11_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_2_lut_LC_11_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40329),
            .in3(N__39957),
            .lcout(n901),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(n12487),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_11_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_11_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_11_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_3_lut_LC_11_22_1 (
            .in0(_gnd_net_),
            .in1(N__52980),
            .in2(N__42687),
            .in3(N__40230),
            .lcout(n900),
            .ltout(),
            .carryin(n12487),
            .carryout(n12488),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_11_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_11_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_11_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_4_lut_LC_11_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42786),
            .in3(N__40227),
            .lcout(n899),
            .ltout(),
            .carryin(n12488),
            .carryout(n12489),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_11_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_11_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_11_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_5_lut_LC_11_22_3 (
            .in0(_gnd_net_),
            .in1(N__52981),
            .in2(N__40449),
            .in3(N__40224),
            .lcout(n898),
            .ltout(),
            .carryin(n12489),
            .carryout(n12490),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_11_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_11_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_11_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_6_lut_LC_11_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40497),
            .in3(N__40221),
            .lcout(n897),
            .ltout(),
            .carryin(n12490),
            .carryout(n12491),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_11_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_11_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_11_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_7_lut_LC_11_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40629),
            .in3(N__40218),
            .lcout(n896),
            .ltout(),
            .carryin(n12491),
            .carryout(n12492),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_11_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_11_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_11_22_6.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_565_8_lut_LC_11_22_6 (
            .in0(N__52982),
            .in1(N__40275),
            .in2(N__40296),
            .in3(N__40215),
            .lcout(n927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i573_3_lut_LC_11_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i573_3_lut_LC_11_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i573_3_lut_LC_11_23_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i573_3_lut_LC_11_23_0 (
            .in0(_gnd_net_),
            .in1(N__40327),
            .in2(N__40212),
            .in3(N__40262),
            .lcout(n933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i568_3_lut_LC_11_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i568_3_lut_LC_11_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i568_3_lut_LC_11_23_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i568_3_lut_LC_11_23_1 (
            .in0(_gnd_net_),
            .in1(N__40628),
            .in2(N__40274),
            .in3(N__40200),
            .lcout(n928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i572_3_lut_LC_11_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i572_3_lut_LC_11_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i572_3_lut_LC_11_23_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i572_3_lut_LC_11_23_2 (
            .in0(_gnd_net_),
            .in1(N__42682),
            .in2(N__40194),
            .in3(N__40261),
            .lcout(n932),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i571_3_lut_LC_11_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i571_3_lut_LC_11_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i571_3_lut_LC_11_23_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i571_3_lut_LC_11_23_3 (
            .in0(_gnd_net_),
            .in1(N__42782),
            .in2(N__40273),
            .in3(N__40185),
            .lcout(n931),
            .ltout(n931_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9972_4_lut_LC_11_23_4.C_ON=1'b0;
    defparam i9972_4_lut_LC_11_23_4.SEQ_MODE=4'b0000;
    defparam i9972_4_lut_LC_11_23_4.LUT_INIT=16'b1111110011111000;
    LogicCell40 i9972_4_lut_LC_11_23_4 (
            .in0(N__44756),
            .in1(N__42745),
            .in2(N__40383),
            .in3(N__44680),
            .lcout(n11940),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_11_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_11_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_11_23_5.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i24_3_lut_LC_11_23_5 (
            .in0(_gnd_net_),
            .in1(N__46151),
            .in2(N__40380),
            .in3(N__41994),
            .lcout(n296),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i569_3_lut_LC_11_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i569_3_lut_LC_11_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i569_3_lut_LC_11_23_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i569_3_lut_LC_11_23_6 (
            .in0(_gnd_net_),
            .in1(N__40493),
            .in2(N__40371),
            .in3(N__40263),
            .lcout(n929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_11_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_11_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_11_23_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i26_3_lut_LC_11_23_7 (
            .in0(_gnd_net_),
            .in1(N__46150),
            .in2(N__40362),
            .in3(N__40335),
            .lcout(n294),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10044_4_lut_LC_11_24_0.C_ON=1'b0;
    defparam i10044_4_lut_LC_11_24_0.SEQ_MODE=4'b0000;
    defparam i10044_4_lut_LC_11_24_0.LUT_INIT=16'b1111111110101000;
    LogicCell40 i10044_4_lut_LC_11_24_0 (
            .in0(N__42778),
            .in1(N__40328),
            .in2(N__42683),
            .in3(N__40441),
            .lcout(n12012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i500_4_lut_LC_11_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i500_4_lut_LC_11_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i500_4_lut_LC_11_24_1.LUT_INIT=16'b1000110010000000;
    LogicCell40 encoder0_position_31__I_0_i500_4_lut_LC_11_24_1 (
            .in0(N__43254),
            .in1(N__42326),
            .in2(N__40305),
            .in3(N__46154),
            .lcout(n828),
            .ltout(n828_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10130_4_lut_LC_11_24_2.C_ON=1'b0;
    defparam i10130_4_lut_LC_11_24_2.SEQ_MODE=4'b0000;
    defparam i10130_4_lut_LC_11_24_2.LUT_INIT=16'b1111100011110000;
    LogicCell40 i10130_4_lut_LC_11_24_2 (
            .in0(N__40489),
            .in1(N__40618),
            .in2(N__40284),
            .in3(N__40281),
            .lcout(n861),
            .ltout(n861_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i570_3_lut_LC_11_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i570_3_lut_LC_11_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i570_3_lut_LC_11_24_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i570_3_lut_LC_11_24_3 (
            .in0(N__40442),
            .in1(_gnd_net_),
            .in2(N__40242),
            .in3(N__40239),
            .lcout(n930),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10980_3_lut_LC_11_24_4.C_ON=1'b0;
    defparam i10980_3_lut_LC_11_24_4.SEQ_MODE=4'b0000;
    defparam i10980_3_lut_LC_11_24_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 i10980_3_lut_LC_11_24_4 (
            .in0(_gnd_net_),
            .in1(N__40706),
            .in2(N__42849),
            .in3(N__43299),
            .lcout(),
            .ltout(n13644_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10981_3_lut_LC_11_24_5.C_ON=1'b0;
    defparam i10981_3_lut_LC_11_24_5.SEQ_MODE=4'b0000;
    defparam i10981_3_lut_LC_11_24_5.LUT_INIT=16'b1111001111000000;
    LogicCell40 i10981_3_lut_LC_11_24_5 (
            .in0(_gnd_net_),
            .in1(N__46153),
            .in2(N__40500),
            .in3(N__40740),
            .lcout(n830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10986_3_lut_LC_11_24_6.C_ON=1'b0;
    defparam i10986_3_lut_LC_11_24_6.SEQ_MODE=4'b0000;
    defparam i10986_3_lut_LC_11_24_6.LUT_INIT=16'b1111101000001010;
    LogicCell40 i10986_3_lut_LC_11_24_6 (
            .in0(N__40473),
            .in1(_gnd_net_),
            .in2(N__42848),
            .in3(N__42630),
            .lcout(n13650),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_11_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_11_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_11_24_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i27_3_lut_LC_11_24_7 (
            .in0(_gnd_net_),
            .in1(N__46152),
            .in2(N__42729),
            .in3(N__40472),
            .lcout(n293),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_64_LC_11_25_0.C_ON=1'b0;
    defparam i1_4_lut_adj_64_LC_11_25_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_64_LC_11_25_0.LUT_INIT=16'b1111101011111000;
    LogicCell40 i1_4_lut_adj_64_LC_11_25_0 (
            .in0(N__40393),
            .in1(N__42866),
            .in2(N__40707),
            .in3(N__42641),
            .lcout(n5_adj_676),
            .ltout(n5_adj_676_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_65_LC_11_25_1.C_ON=1'b0;
    defparam i1_3_lut_adj_65_LC_11_25_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_65_LC_11_25_1.LUT_INIT=16'b1100000000000000;
    LogicCell40 i1_3_lut_adj_65_LC_11_25_1 (
            .in0(_gnd_net_),
            .in1(N__40680),
            .in2(N__40458),
            .in3(N__42316),
            .lcout(n13641),
            .ltout(n13641_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10982_3_lut_LC_11_25_2.C_ON=1'b0;
    defparam i10982_3_lut_LC_11_25_2.SEQ_MODE=4'b0000;
    defparam i10982_3_lut_LC_11_25_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 i10982_3_lut_LC_11_25_2 (
            .in0(N__40397),
            .in1(_gnd_net_),
            .in2(N__40455),
            .in3(N__42588),
            .lcout(),
            .ltout(n13646_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10983_3_lut_LC_11_25_3.C_ON=1'b0;
    defparam i10983_3_lut_LC_11_25_3.SEQ_MODE=4'b0000;
    defparam i10983_3_lut_LC_11_25_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 i10983_3_lut_LC_11_25_3 (
            .in0(N__46102),
            .in1(_gnd_net_),
            .in2(N__40452),
            .in3(N__40427),
            .lcout(n831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_11_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_11_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_11_25_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i29_3_lut_LC_11_25_4 (
            .in0(_gnd_net_),
            .in1(N__40426),
            .in2(N__40398),
            .in3(N__46098),
            .lcout(n174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_25_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_25_5 (
            .in0(_gnd_net_),
            .in1(N__40736),
            .in2(N__46165),
            .in3(N__40705),
            .lcout(n404),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10978_3_lut_LC_11_25_6.C_ON=1'b0;
    defparam i10978_3_lut_LC_11_25_6.SEQ_MODE=4'b0000;
    defparam i10978_3_lut_LC_11_25_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 i10978_3_lut_LC_11_25_6 (
            .in0(_gnd_net_),
            .in1(N__42847),
            .in2(N__40688),
            .in3(N__43278),
            .lcout(),
            .ltout(n13642_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10979_3_lut_LC_11_25_7.C_ON=1'b0;
    defparam i10979_3_lut_LC_11_25_7.SEQ_MODE=4'b0000;
    defparam i10979_3_lut_LC_11_25_7.LUT_INIT=16'b1110010011100100;
    LogicCell40 i10979_3_lut_LC_11_25_7 (
            .in0(N__46103),
            .in1(N__40664),
            .in2(N__40632),
            .in3(_gnd_net_),
            .lcout(n829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_11_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_11_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_11_26_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i2_3_lut_LC_11_26_0 (
            .in0(N__46180),
            .in1(N__40602),
            .in2(_gnd_net_),
            .in3(N__40590),
            .lcout(n318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_11_26_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_11_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_11_26_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_11_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40524),
            .lcout(n11_adj_572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_50_LC_11_26_3.C_ON=1'b0;
    defparam i4_4_lut_adj_50_LC_11_26_3.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_50_LC_11_26_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 i4_4_lut_adj_50_LC_11_26_3 (
            .in0(N__49019),
            .in1(N__48940),
            .in2(N__49068),
            .in3(N__46866),
            .lcout(),
            .ltout(n10_adj_606_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_52_LC_11_26_4.C_ON=1'b0;
    defparam i1_4_lut_adj_52_LC_11_26_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_52_LC_11_26_4.LUT_INIT=16'b1110110011001100;
    LogicCell40 i1_4_lut_adj_52_LC_11_26_4 (
            .in0(N__48977),
            .in1(N__54806),
            .in2(N__40512),
            .in3(N__48896),
            .lcout(),
            .ltout(n15_adj_565_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_55_LC_11_26_5.C_ON=1'b0;
    defparam i11_4_lut_adj_55_LC_11_26_5.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_55_LC_11_26_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_55_LC_11_26_5 (
            .in0(N__49547),
            .in1(N__49380),
            .in2(N__40509),
            .in3(N__40506),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_51_LC_11_26_6.C_ON=1'b0;
    defparam i2_2_lut_adj_51_LC_11_26_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_51_LC_11_26_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_adj_51_LC_11_26_6 (
            .in0(_gnd_net_),
            .in1(N__49435),
            .in2(_gnd_net_),
            .in3(N__54848),
            .lcout(n16_adj_564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_11_27_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_11_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_11_27_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_11_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40833),
            .lcout(n15_adj_568),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i3_LC_11_27_1.C_ON=1'b0;
    defparam pwm_setpoint_i3_LC_11_27_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i3_LC_11_27_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 pwm_setpoint_i3_LC_11_27_1 (
            .in0(N__40821),
            .in1(N__43514),
            .in2(_gnd_net_),
            .in3(N__55263),
            .lcout(pwm_setpoint_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55795),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_11_27_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_11_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_11_27_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_11_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40809),
            .lcout(n14_adj_569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i13_LC_11_27_3.C_ON=1'b0;
    defparam pwm_setpoint_i13_LC_11_27_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i13_LC_11_27_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i13_LC_11_27_3 (
            .in0(N__43697),
            .in1(N__55262),
            .in2(_gnd_net_),
            .in3(N__40797),
            .lcout(pwm_setpoint_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55795),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i15_2_lut_LC_11_27_4.C_ON=1'b0;
    defparam LessThan_299_i15_2_lut_LC_11_27_4.SEQ_MODE=4'b0000;
    defparam LessThan_299_i15_2_lut_LC_11_27_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i15_2_lut_LC_11_27_4 (
            .in0(_gnd_net_),
            .in1(N__46748),
            .in2(_gnd_net_),
            .in3(N__40896),
            .lcout(n15_adj_663),
            .ltout(n15_adj_663_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12400_4_lut_LC_11_27_5.C_ON=1'b0;
    defparam i12400_4_lut_LC_11_27_5.SEQ_MODE=4'b0000;
    defparam i12400_4_lut_LC_11_27_5.LUT_INIT=16'b1111111100000001;
    LogicCell40 i12400_4_lut_LC_11_27_5 (
            .in0(N__47445),
            .in1(N__47421),
            .in2(N__40785),
            .in3(N__43763),
            .lcout(n15125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_11_27_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_11_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_11_27_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_11_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40776),
            .lcout(n7_adj_576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_11_27_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_11_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_11_27_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_11_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40764),
            .lcout(n5_adj_578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_11_28_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_11_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_11_28_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_11_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40752),
            .lcout(n2_adj_581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i12_3_lut_3_lut_LC_11_28_1.C_ON=1'b0;
    defparam LessThan_299_i12_3_lut_3_lut_LC_11_28_1.SEQ_MODE=4'b0000;
    defparam LessThan_299_i12_3_lut_3_lut_LC_11_28_1.LUT_INIT=16'b1101110101000100;
    LogicCell40 LessThan_299_i12_3_lut_3_lut_LC_11_28_1 (
            .in0(N__46591),
            .in1(N__40909),
            .in2(_gnd_net_),
            .in3(N__40894),
            .lcout(n12_adj_661),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i37_2_lut_LC_11_28_2.C_ON=1'b0;
    defparam LessThan_299_i37_2_lut_LC_11_28_2.SEQ_MODE=4'b0000;
    defparam LessThan_299_i37_2_lut_LC_11_28_2.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i37_2_lut_LC_11_28_2 (
            .in0(N__44054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46476),
            .lcout(n37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i7_LC_11_28_3.C_ON=1'b0;
    defparam pwm_setpoint_i7_LC_11_28_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i7_LC_11_28_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i7_LC_11_28_3 (
            .in0(N__43391),
            .in1(N__55261),
            .in2(_gnd_net_),
            .in3(N__40923),
            .lcout(pwm_setpoint_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55798),
            .ce(),
            .sr(_gnd_net_));
    defparam i12394_2_lut_4_lut_LC_11_28_5.C_ON=1'b0;
    defparam i12394_2_lut_4_lut_LC_11_28_5.SEQ_MODE=4'b0000;
    defparam i12394_2_lut_4_lut_LC_11_28_5.LUT_INIT=16'b0110111111110110;
    LogicCell40 i12394_2_lut_4_lut_LC_11_28_5 (
            .in0(N__46592),
            .in1(N__40910),
            .in2(N__46752),
            .in3(N__40895),
            .lcout(n15119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i6_3_lut_3_lut_LC_11_28_6.C_ON=1'b0;
    defparam LessThan_299_i6_3_lut_3_lut_LC_11_28_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i6_3_lut_3_lut_LC_11_28_6.LUT_INIT=16'b1000100011101110;
    LogicCell40 LessThan_299_i6_3_lut_3_lut_LC_11_28_6 (
            .in0(N__46841),
            .in1(N__46826),
            .in2(_gnd_net_),
            .in3(N__46797),
            .lcout(n6_adj_656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_11_28_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_11_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_11_28_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_11_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40875),
            .lcout(n16_adj_563),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i0_LC_11_29_0.C_ON=1'b1;
    defparam blink_counter_660__i0_LC_11_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i0_LC_11_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i0_LC_11_29_0 (
            .in0(_gnd_net_),
            .in1(N__40860),
            .in2(_gnd_net_),
            .in3(N__40854),
            .lcout(n26_adj_697),
            .ltout(),
            .carryin(bfn_11_29_0_),
            .carryout(n13087),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i1_LC_11_29_1.C_ON=1'b1;
    defparam blink_counter_660__i1_LC_11_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i1_LC_11_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i1_LC_11_29_1 (
            .in0(_gnd_net_),
            .in1(N__40851),
            .in2(_gnd_net_),
            .in3(N__40845),
            .lcout(n25_adj_696),
            .ltout(),
            .carryin(n13087),
            .carryout(n13088),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i2_LC_11_29_2.C_ON=1'b1;
    defparam blink_counter_660__i2_LC_11_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i2_LC_11_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i2_LC_11_29_2 (
            .in0(_gnd_net_),
            .in1(N__40842),
            .in2(_gnd_net_),
            .in3(N__40836),
            .lcout(n24_adj_695),
            .ltout(),
            .carryin(n13088),
            .carryout(n13089),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i3_LC_11_29_3.C_ON=1'b1;
    defparam blink_counter_660__i3_LC_11_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i3_LC_11_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i3_LC_11_29_3 (
            .in0(_gnd_net_),
            .in1(N__41010),
            .in2(_gnd_net_),
            .in3(N__41004),
            .lcout(n23_adj_694),
            .ltout(),
            .carryin(n13089),
            .carryout(n13090),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i4_LC_11_29_4.C_ON=1'b1;
    defparam blink_counter_660__i4_LC_11_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i4_LC_11_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i4_LC_11_29_4 (
            .in0(_gnd_net_),
            .in1(N__41001),
            .in2(_gnd_net_),
            .in3(N__40995),
            .lcout(n22_adj_693),
            .ltout(),
            .carryin(n13090),
            .carryout(n13091),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i5_LC_11_29_5.C_ON=1'b1;
    defparam blink_counter_660__i5_LC_11_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i5_LC_11_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i5_LC_11_29_5 (
            .in0(_gnd_net_),
            .in1(N__40992),
            .in2(_gnd_net_),
            .in3(N__40986),
            .lcout(n21_adj_692),
            .ltout(),
            .carryin(n13091),
            .carryout(n13092),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i6_LC_11_29_6.C_ON=1'b1;
    defparam blink_counter_660__i6_LC_11_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i6_LC_11_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i6_LC_11_29_6 (
            .in0(_gnd_net_),
            .in1(N__40983),
            .in2(_gnd_net_),
            .in3(N__40977),
            .lcout(n20_adj_691),
            .ltout(),
            .carryin(n13092),
            .carryout(n13093),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i7_LC_11_29_7.C_ON=1'b1;
    defparam blink_counter_660__i7_LC_11_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i7_LC_11_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i7_LC_11_29_7 (
            .in0(_gnd_net_),
            .in1(N__40974),
            .in2(_gnd_net_),
            .in3(N__40968),
            .lcout(n19_adj_690),
            .ltout(),
            .carryin(n13093),
            .carryout(n13094),
            .clk(N__55802),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i8_LC_11_30_0.C_ON=1'b1;
    defparam blink_counter_660__i8_LC_11_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i8_LC_11_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i8_LC_11_30_0 (
            .in0(_gnd_net_),
            .in1(N__40965),
            .in2(_gnd_net_),
            .in3(N__40959),
            .lcout(n18_adj_689),
            .ltout(),
            .carryin(bfn_11_30_0_),
            .carryout(n13095),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i9_LC_11_30_1.C_ON=1'b1;
    defparam blink_counter_660__i9_LC_11_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i9_LC_11_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i9_LC_11_30_1 (
            .in0(_gnd_net_),
            .in1(N__40956),
            .in2(_gnd_net_),
            .in3(N__40950),
            .lcout(n17_adj_688),
            .ltout(),
            .carryin(n13095),
            .carryout(n13096),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i10_LC_11_30_2.C_ON=1'b1;
    defparam blink_counter_660__i10_LC_11_30_2.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i10_LC_11_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i10_LC_11_30_2 (
            .in0(_gnd_net_),
            .in1(N__40947),
            .in2(_gnd_net_),
            .in3(N__40941),
            .lcout(n16_adj_687),
            .ltout(),
            .carryin(n13096),
            .carryout(n13097),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i11_LC_11_30_3.C_ON=1'b1;
    defparam blink_counter_660__i11_LC_11_30_3.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i11_LC_11_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i11_LC_11_30_3 (
            .in0(_gnd_net_),
            .in1(N__40938),
            .in2(_gnd_net_),
            .in3(N__40932),
            .lcout(n15_adj_686),
            .ltout(),
            .carryin(n13097),
            .carryout(n13098),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i12_LC_11_30_4.C_ON=1'b1;
    defparam blink_counter_660__i12_LC_11_30_4.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i12_LC_11_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i12_LC_11_30_4 (
            .in0(_gnd_net_),
            .in1(N__41082),
            .in2(_gnd_net_),
            .in3(N__41076),
            .lcout(n14_adj_685),
            .ltout(),
            .carryin(n13098),
            .carryout(n13099),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i13_LC_11_30_5.C_ON=1'b1;
    defparam blink_counter_660__i13_LC_11_30_5.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i13_LC_11_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i13_LC_11_30_5 (
            .in0(_gnd_net_),
            .in1(N__41073),
            .in2(_gnd_net_),
            .in3(N__41067),
            .lcout(n13_adj_684),
            .ltout(),
            .carryin(n13099),
            .carryout(n13100),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i14_LC_11_30_6.C_ON=1'b1;
    defparam blink_counter_660__i14_LC_11_30_6.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i14_LC_11_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i14_LC_11_30_6 (
            .in0(_gnd_net_),
            .in1(N__41064),
            .in2(_gnd_net_),
            .in3(N__41058),
            .lcout(n12_adj_683),
            .ltout(),
            .carryin(n13100),
            .carryout(n13101),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i15_LC_11_30_7.C_ON=1'b1;
    defparam blink_counter_660__i15_LC_11_30_7.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i15_LC_11_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i15_LC_11_30_7 (
            .in0(_gnd_net_),
            .in1(N__41055),
            .in2(_gnd_net_),
            .in3(N__41049),
            .lcout(n11_adj_682),
            .ltout(),
            .carryin(n13101),
            .carryout(n13102),
            .clk(N__55807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i16_LC_11_31_0.C_ON=1'b1;
    defparam blink_counter_660__i16_LC_11_31_0.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i16_LC_11_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i16_LC_11_31_0 (
            .in0(_gnd_net_),
            .in1(N__41046),
            .in2(_gnd_net_),
            .in3(N__41040),
            .lcout(n10_adj_681),
            .ltout(),
            .carryin(bfn_11_31_0_),
            .carryout(n13103),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i17_LC_11_31_1.C_ON=1'b1;
    defparam blink_counter_660__i17_LC_11_31_1.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i17_LC_11_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i17_LC_11_31_1 (
            .in0(_gnd_net_),
            .in1(N__41037),
            .in2(_gnd_net_),
            .in3(N__41031),
            .lcout(n9_adj_680),
            .ltout(),
            .carryin(n13103),
            .carryout(n13104),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i18_LC_11_31_2.C_ON=1'b1;
    defparam blink_counter_660__i18_LC_11_31_2.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i18_LC_11_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i18_LC_11_31_2 (
            .in0(_gnd_net_),
            .in1(N__41028),
            .in2(_gnd_net_),
            .in3(N__41022),
            .lcout(n8_adj_679),
            .ltout(),
            .carryin(n13104),
            .carryout(n13105),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i19_LC_11_31_3.C_ON=1'b1;
    defparam blink_counter_660__i19_LC_11_31_3.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i19_LC_11_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i19_LC_11_31_3 (
            .in0(_gnd_net_),
            .in1(N__41019),
            .in2(_gnd_net_),
            .in3(N__41013),
            .lcout(n7_adj_678),
            .ltout(),
            .carryin(n13105),
            .carryout(n13106),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i20_LC_11_31_4.C_ON=1'b1;
    defparam blink_counter_660__i20_LC_11_31_4.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i20_LC_11_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i20_LC_11_31_4 (
            .in0(_gnd_net_),
            .in1(N__41214),
            .in2(_gnd_net_),
            .in3(N__41208),
            .lcout(n6_adj_677),
            .ltout(),
            .carryin(n13106),
            .carryout(n13107),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i21_LC_11_31_5.C_ON=1'b1;
    defparam blink_counter_660__i21_LC_11_31_5.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i21_LC_11_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i21_LC_11_31_5 (
            .in0(_gnd_net_),
            .in1(N__41197),
            .in2(_gnd_net_),
            .in3(N__41184),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n13107),
            .carryout(n13108),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i22_LC_11_31_6.C_ON=1'b1;
    defparam blink_counter_660__i22_LC_11_31_6.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i22_LC_11_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i22_LC_11_31_6 (
            .in0(_gnd_net_),
            .in1(N__41179),
            .in2(_gnd_net_),
            .in3(N__41166),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n13108),
            .carryout(n13109),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i23_LC_11_31_7.C_ON=1'b1;
    defparam blink_counter_660__i23_LC_11_31_7.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i23_LC_11_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i23_LC_11_31_7 (
            .in0(_gnd_net_),
            .in1(N__41161),
            .in2(_gnd_net_),
            .in3(N__41148),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n13109),
            .carryout(n13110),
            .clk(N__55814),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i24_LC_11_32_0.C_ON=1'b1;
    defparam blink_counter_660__i24_LC_11_32_0.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i24_LC_11_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i24_LC_11_32_0 (
            .in0(_gnd_net_),
            .in1(N__41143),
            .in2(_gnd_net_),
            .in3(N__41130),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_11_32_0_),
            .carryout(n13111),
            .clk(N__55818),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_660__i25_LC_11_32_1.C_ON=1'b0;
    defparam blink_counter_660__i25_LC_11_32_1.SEQ_MODE=4'b1000;
    defparam blink_counter_660__i25_LC_11_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_660__i25_LC_11_32_1 (
            .in0(_gnd_net_),
            .in1(N__41120),
            .in2(_gnd_net_),
            .in3(N__41127),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55818),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i19_LC_11_32_3.C_ON=1'b0;
    defparam pwm_setpoint_i19_LC_11_32_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i19_LC_11_32_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i19_LC_11_32_3 (
            .in0(N__43908),
            .in1(N__55334),
            .in2(_gnd_net_),
            .in3(N__41109),
            .lcout(pwm_setpoint_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55818),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i18_1_lut_LC_11_32_6.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i18_1_lut_LC_11_32_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i18_1_lut_LC_11_32_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i18_1_lut_LC_11_32_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43974),
            .lcout(n8_adj_588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i21_1_lut_LC_11_32_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i21_1_lut_LC_11_32_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i21_1_lut_LC_11_32_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i21_1_lut_LC_11_32_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44138),
            .lcout(n5_adj_585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_12_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_12_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_12_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_2_lut_LC_12_17_0 (
            .in0(_gnd_net_),
            .in1(N__42419),
            .in2(_gnd_net_),
            .in3(N__41439),
            .lcout(n1901),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(n12592),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_12_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_12_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_12_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_3_lut_LC_12_17_1 (
            .in0(_gnd_net_),
            .in1(N__53101),
            .in2(N__41436),
            .in3(N__41400),
            .lcout(n1900),
            .ltout(),
            .carryin(n12592),
            .carryout(n12593),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_12_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_12_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_12_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_4_lut_LC_12_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41397),
            .in3(N__41367),
            .lcout(n1899),
            .ltout(),
            .carryin(n12593),
            .carryout(n12594),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_12_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_12_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_12_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_5_lut_LC_12_17_3 (
            .in0(_gnd_net_),
            .in1(N__53102),
            .in2(N__41364),
            .in3(N__41325),
            .lcout(n1898),
            .ltout(),
            .carryin(n12594),
            .carryout(n12595),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_12_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_12_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_6_lut_LC_12_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41322),
            .in3(N__41295),
            .lcout(n1897),
            .ltout(),
            .carryin(n12595),
            .carryout(n12596),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_12_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_12_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_7_lut_LC_12_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41292),
            .in3(N__41265),
            .lcout(n1896),
            .ltout(),
            .carryin(n12596),
            .carryout(n12597),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_12_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_12_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_12_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_8_lut_LC_12_17_6 (
            .in0(_gnd_net_),
            .in1(N__53937),
            .in2(N__41262),
            .in3(N__41229),
            .lcout(n1895),
            .ltout(),
            .carryin(n12597),
            .carryout(n12598),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_12_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_12_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_12_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_9_lut_LC_12_17_7 (
            .in0(_gnd_net_),
            .in1(N__53103),
            .in2(N__41834),
            .in3(N__41217),
            .lcout(n1894),
            .ltout(),
            .carryin(n12598),
            .carryout(n12599),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_12_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_12_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_12_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_10_lut_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(N__53577),
            .in2(N__41693),
            .in3(N__41664),
            .lcout(n1893),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(n12600),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_12_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_12_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_12_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_11_lut_LC_12_18_1 (
            .in0(_gnd_net_),
            .in1(N__53584),
            .in2(N__41661),
            .in3(N__41631),
            .lcout(n1892),
            .ltout(),
            .carryin(n12600),
            .carryout(n12601),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_12_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_12_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_12_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_12_lut_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(N__53578),
            .in2(N__41628),
            .in3(N__41595),
            .lcout(n1891),
            .ltout(),
            .carryin(n12601),
            .carryout(n12602),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_12_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_12_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_12_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_13_lut_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(N__53585),
            .in2(N__41592),
            .in3(N__41556),
            .lcout(n1890),
            .ltout(),
            .carryin(n12602),
            .carryout(n12603),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_12_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_12_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_12_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_14_lut_LC_12_18_4 (
            .in0(_gnd_net_),
            .in1(N__53579),
            .in2(N__41552),
            .in3(N__41511),
            .lcout(n1889),
            .ltout(),
            .carryin(n12603),
            .carryout(n12604),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_12_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_12_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_12_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_15_lut_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(N__41855),
            .in2(N__53936),
            .in3(N__41502),
            .lcout(n1888),
            .ltout(),
            .carryin(n12604),
            .carryout(n12605),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_12_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_12_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_16_lut_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(N__53583),
            .in2(N__41499),
            .in3(N__41475),
            .lcout(n1887),
            .ltout(),
            .carryin(n12605),
            .carryout(n12606),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_12_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_12_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_12_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_17_lut_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(N__53586),
            .in2(N__41472),
            .in3(N__41451),
            .lcout(n1886),
            .ltout(),
            .carryin(n12606),
            .carryout(n12607),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_12_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_12_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_12_19_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 encoder0_position_31__I_0_add_1235_18_lut_LC_12_19_0 (
            .in0(N__52810),
            .in1(N__44518),
            .in2(_gnd_net_),
            .in3(N__41874),
            .lcout(n1885),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_12_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_12_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_12_19_2.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1104_3_lut_LC_12_19_2 (
            .in0(N__48027),
            .in1(N__48003),
            .in2(N__50195),
            .in3(_gnd_net_),
            .lcout(n1720),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3 (
            .in0(_gnd_net_),
            .in1(N__48112),
            .in2(N__48090),
            .in3(N__50187),
            .lcout(n1722),
            .ltout(n1722_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4 (
            .in0(N__41759),
            .in1(_gnd_net_),
            .in2(N__41859),
            .in3(N__44382),
            .lcout(n1821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_12_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_12_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_12_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1105_3_lut_LC_12_19_5 (
            .in0(_gnd_net_),
            .in1(N__48072),
            .in2(N__48045),
            .in3(N__50188),
            .lcout(n1721),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_12_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_12_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_12_19_7.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1179_3_lut_LC_12_19_7 (
            .in0(N__44478),
            .in1(_gnd_net_),
            .in2(N__50109),
            .in3(N__41758),
            .lcout(n1827),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12897_1_lut_LC_12_20_0.C_ON=1'b0;
    defparam i12897_1_lut_LC_12_20_0.SEQ_MODE=4'b0000;
    defparam i12897_1_lut_LC_12_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12897_1_lut_LC_12_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41785),
            .lcout(n15622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_12_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_12_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_12_20_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1039_3_lut_LC_12_20_1 (
            .in0(_gnd_net_),
            .in1(N__44640),
            .in2(N__48420),
            .in3(N__50672),
            .lcout(n1623_adj_610),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_12_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_12_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_12_20_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_12_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42290),
            .lcout(n16_adj_637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2177_2_lut_LC_12_20_5.C_ON=1'b0;
    defparam i2177_2_lut_LC_12_20_5.SEQ_MODE=4'b0000;
    defparam i2177_2_lut_LC_12_20_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2177_2_lut_LC_12_20_5 (
            .in0(_gnd_net_),
            .in1(N__46196),
            .in2(_gnd_net_),
            .in3(N__42330),
            .lcout(n402),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_12_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_12_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_12_20_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i18_3_lut_LC_12_20_6 (
            .in0(N__46197),
            .in1(N__42303),
            .in2(_gnd_net_),
            .in3(N__42291),
            .lcout(n302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_12_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_12_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_12_20_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i4_3_lut_LC_12_20_7 (
            .in0(N__42267),
            .in1(N__46198),
            .in2(_gnd_net_),
            .in3(N__42255),
            .lcout(n316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_12_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_12_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_12_21_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_12_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46183),
            .lcout(n2_adj_623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_12_21_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_12_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_12_21_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_12_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42009),
            .lcout(n18_adj_559),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_21_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41993),
            .lcout(n10_adj_631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_12_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_12_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_12_21_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_12_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42443),
            .lcout(n18_adj_639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_21_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_21_5 (
            .in0(N__46185),
            .in1(N__41931),
            .in2(_gnd_net_),
            .in3(N__41918),
            .lcout(n303),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_12_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_12_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_12_21_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i16_3_lut_LC_12_21_6 (
            .in0(N__41886),
            .in1(N__46186),
            .in2(_gnd_net_),
            .in3(N__42444),
            .lcout(n304),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_21_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_21_7 (
            .in0(N__46184),
            .in1(N__42390),
            .in2(_gnd_net_),
            .in3(N__42378),
            .lcout(n301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_12_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_12_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_12_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_2_lut_LC_12_22_0 (
            .in0(_gnd_net_),
            .in1(N__44744),
            .in2(_gnd_net_),
            .in3(N__42351),
            .lcout(n1001),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(n12493),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_12_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_12_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_12_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_3_lut_LC_12_22_1 (
            .in0(_gnd_net_),
            .in1(N__52901),
            .in2(N__44687),
            .in3(N__42348),
            .lcout(n1000),
            .ltout(),
            .carryin(n12493),
            .carryout(n12494),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_12_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_12_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_12_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_4_lut_LC_12_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42752),
            .in3(N__42345),
            .lcout(n999),
            .ltout(),
            .carryin(n12494),
            .carryout(n12495),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_12_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_12_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_12_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_5_lut_LC_12_22_3 (
            .in0(_gnd_net_),
            .in1(N__52902),
            .in2(N__42473),
            .in3(N__42342),
            .lcout(n998),
            .ltout(),
            .carryin(n12495),
            .carryout(n12496),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_12_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_12_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_12_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_6_lut_LC_12_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42546),
            .in3(N__42339),
            .lcout(n997),
            .ltout(),
            .carryin(n12496),
            .carryout(n12497),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_12_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_12_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_12_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_7_lut_LC_12_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42516),
            .in3(N__42336),
            .lcout(n996),
            .ltout(),
            .carryin(n12497),
            .carryout(n12498),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_12_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_12_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_12_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_8_lut_LC_12_22_6 (
            .in0(_gnd_net_),
            .in1(N__52903),
            .in2(N__44987),
            .in3(N__42333),
            .lcout(n995),
            .ltout(),
            .carryin(n12498),
            .carryout(n12499),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_12_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_12_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_12_22_7.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_632_9_lut_LC_12_22_7 (
            .in0(N__52904),
            .in1(N__42567),
            .in2(N__44964),
            .in3(N__42579),
            .lcout(n1026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i641_3_lut_LC_12_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i641_3_lut_LC_12_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i641_3_lut_LC_12_23_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i641_3_lut_LC_12_23_0 (
            .in0(_gnd_net_),
            .in1(N__44757),
            .in2(N__42576),
            .in3(N__44952),
            .lcout(n1033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_167_LC_12_23_1.C_ON=1'b0;
    defparam i1_2_lut_adj_167_LC_12_23_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_167_LC_12_23_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_167_LC_12_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42515),
            .in3(N__42538),
            .lcout(),
            .ltout(n14466_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_169_LC_12_23_2.C_ON=1'b0;
    defparam i1_4_lut_adj_169_LC_12_23_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_169_LC_12_23_2.LUT_INIT=16'b1111111011101110;
    LogicCell40 i1_4_lut_adj_169_LC_12_23_2 (
            .in0(N__44980),
            .in1(N__42566),
            .in2(N__42555),
            .in3(N__42552),
            .lcout(n960),
            .ltout(n960_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i637_3_lut_LC_12_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i637_3_lut_LC_12_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i637_3_lut_LC_12_23_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i637_3_lut_LC_12_23_3 (
            .in0(_gnd_net_),
            .in1(N__42539),
            .in2(N__42525),
            .in3(N__42522),
            .lcout(n1029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i636_3_lut_LC_12_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i636_3_lut_LC_12_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i636_3_lut_LC_12_23_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i636_3_lut_LC_12_23_4 (
            .in0(_gnd_net_),
            .in1(N__42511),
            .in2(N__42495),
            .in3(N__44954),
            .lcout(n1028),
            .ltout(n1028_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i703_3_lut_LC_12_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i703_3_lut_LC_12_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i703_3_lut_LC_12_23_5.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i703_3_lut_LC_12_23_5 (
            .in0(_gnd_net_),
            .in1(N__46408),
            .in2(N__42486),
            .in3(N__45096),
            .lcout(n1127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i638_3_lut_LC_12_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i638_3_lut_LC_12_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i638_3_lut_LC_12_23_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i638_3_lut_LC_12_23_6 (
            .in0(_gnd_net_),
            .in1(N__42483),
            .in2(N__42477),
            .in3(N__44953),
            .lcout(n1030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_12_24_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_12_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_12_24_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_12_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42456),
            .lcout(n17_adj_560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10984_3_lut_LC_12_24_1.C_ON=1'b0;
    defparam i10984_3_lut_LC_12_24_1.SEQ_MODE=4'b0000;
    defparam i10984_3_lut_LC_12_24_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 i10984_3_lut_LC_12_24_1 (
            .in0(_gnd_net_),
            .in1(N__42870),
            .in2(N__42609),
            .in3(N__42846),
            .lcout(),
            .ltout(n13648_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10985_3_lut_LC_12_24_2.C_ON=1'b0;
    defparam i10985_3_lut_LC_12_24_2.SEQ_MODE=4'b0000;
    defparam i10985_3_lut_LC_12_24_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 i10985_3_lut_LC_12_24_2 (
            .in0(_gnd_net_),
            .in1(N__46173),
            .in2(N__42822),
            .in3(N__42819),
            .lcout(n832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i639_3_lut_LC_12_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i639_3_lut_LC_12_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i639_3_lut_LC_12_24_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i639_3_lut_LC_12_24_4 (
            .in0(_gnd_net_),
            .in1(N__42762),
            .in2(N__42753),
            .in3(N__44955),
            .lcout(n1031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12441_3_lut_LC_12_24_5.C_ON=1'b0;
    defparam i12441_3_lut_LC_12_24_5.SEQ_MODE=4'b0000;
    defparam i12441_3_lut_LC_12_24_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 i12441_3_lut_LC_12_24_5 (
            .in0(_gnd_net_),
            .in1(N__42728),
            .in2(N__46199),
            .in3(N__42693),
            .lcout(n833),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_12_24_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_12_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_12_24_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_12_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42660),
            .lcout(n22_adj_555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_738_2_lut_LC_12_25_0.C_ON=1'b1;
    defparam add_738_2_lut_LC_12_25_0.SEQ_MODE=4'b0000;
    defparam add_738_2_lut_LC_12_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_738_2_lut_LC_12_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42645),
            .in3(N__42624),
            .lcout(n2542),
            .ltout(),
            .carryin(bfn_12_25_0_),
            .carryout(n12482),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_738_3_lut_LC_12_25_1.C_ON=1'b1;
    defparam add_738_3_lut_LC_12_25_1.SEQ_MODE=4'b0000;
    defparam add_738_3_lut_LC_12_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_738_3_lut_LC_12_25_1 (
            .in0(_gnd_net_),
            .in1(N__52427),
            .in2(N__42621),
            .in3(N__42600),
            .lcout(n2541),
            .ltout(),
            .carryin(n12482),
            .carryout(n12483),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_738_4_lut_LC_12_25_2.C_ON=1'b1;
    defparam add_738_4_lut_LC_12_25_2.SEQ_MODE=4'b0000;
    defparam add_738_4_lut_LC_12_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_738_4_lut_LC_12_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42597),
            .in3(N__42582),
            .lcout(n2540),
            .ltout(),
            .carryin(n12483),
            .carryout(n12484),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_738_5_lut_LC_12_25_3.C_ON=1'b1;
    defparam add_738_5_lut_LC_12_25_3.SEQ_MODE=4'b0000;
    defparam add_738_5_lut_LC_12_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_738_5_lut_LC_12_25_3 (
            .in0(_gnd_net_),
            .in1(N__52428),
            .in2(N__43308),
            .in3(N__43293),
            .lcout(n2539),
            .ltout(),
            .carryin(n12484),
            .carryout(n12485),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_738_6_lut_LC_12_25_4.C_ON=1'b1;
    defparam add_738_6_lut_LC_12_25_4.SEQ_MODE=4'b0000;
    defparam add_738_6_lut_LC_12_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_738_6_lut_LC_12_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43290),
            .in3(N__43272),
            .lcout(n2538),
            .ltout(),
            .carryin(n12485),
            .carryout(n12486),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_738_7_lut_LC_12_25_5.C_ON=1'b0;
    defparam add_738_7_lut_LC_12_25_5.SEQ_MODE=4'b0000;
    defparam add_738_7_lut_LC_12_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_738_7_lut_LC_12_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43269),
            .in3(N__43257),
            .lcout(n2537),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_12_25_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_12_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_12_25_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_12_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43248),
            .lcout(n19_adj_558),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_12_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_12_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_12_25_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2112_3_lut_LC_12_25_7 (
            .in0(_gnd_net_),
            .in1(N__43233),
            .in2(N__43197),
            .in3(N__43179),
            .lcout(n3208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i0_LC_12_26_0.C_ON=1'b1;
    defparam duty_i0_LC_12_26_0.SEQ_MODE=4'b1000;
    defparam duty_i0_LC_12_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i0_LC_12_26_0 (
            .in0(_gnd_net_),
            .in1(N__42978),
            .in2(N__48825),
            .in3(N__42948),
            .lcout(duty_0),
            .ltout(),
            .carryin(bfn_12_26_0_),
            .carryout(n12459),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i1_LC_12_26_1.C_ON=1'b1;
    defparam duty_i1_LC_12_26_1.SEQ_MODE=4'b1000;
    defparam duty_i1_LC_12_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i1_LC_12_26_1 (
            .in0(_gnd_net_),
            .in1(N__42945),
            .in2(N__48792),
            .in3(N__42912),
            .lcout(duty_1),
            .ltout(),
            .carryin(n12459),
            .carryout(n12460),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i2_LC_12_26_2.C_ON=1'b1;
    defparam duty_i2_LC_12_26_2.SEQ_MODE=4'b1000;
    defparam duty_i2_LC_12_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i2_LC_12_26_2 (
            .in0(_gnd_net_),
            .in1(N__48756),
            .in2(N__42909),
            .in3(N__42873),
            .lcout(duty_2),
            .ltout(),
            .carryin(n12460),
            .carryout(n12461),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i3_LC_12_26_3.C_ON=1'b1;
    defparam duty_i3_LC_12_26_3.SEQ_MODE=4'b1000;
    defparam duty_i3_LC_12_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i3_LC_12_26_3 (
            .in0(_gnd_net_),
            .in1(N__43527),
            .in2(N__49170),
            .in3(N__43500),
            .lcout(duty_3),
            .ltout(),
            .carryin(n12461),
            .carryout(n12462),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i4_LC_12_26_4.C_ON=1'b1;
    defparam duty_i4_LC_12_26_4.SEQ_MODE=4'b1000;
    defparam duty_i4_LC_12_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i4_LC_12_26_4 (
            .in0(_gnd_net_),
            .in1(N__49137),
            .in2(N__43497),
            .in3(N__43461),
            .lcout(duty_4),
            .ltout(),
            .carryin(n12462),
            .carryout(n12463),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i5_LC_12_26_5.C_ON=1'b1;
    defparam duty_i5_LC_12_26_5.SEQ_MODE=4'b1000;
    defparam duty_i5_LC_12_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i5_LC_12_26_5 (
            .in0(_gnd_net_),
            .in1(N__43458),
            .in2(N__49104),
            .in3(N__43434),
            .lcout(duty_5),
            .ltout(),
            .carryin(n12463),
            .carryout(n12464),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i6_LC_12_26_6.C_ON=1'b1;
    defparam duty_i6_LC_12_26_6.SEQ_MODE=4'b1000;
    defparam duty_i6_LC_12_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i6_LC_12_26_6 (
            .in0(_gnd_net_),
            .in1(N__43431),
            .in2(N__49067),
            .in3(N__43407),
            .lcout(duty_6),
            .ltout(),
            .carryin(n12464),
            .carryout(n12465),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i7_LC_12_26_7.C_ON=1'b1;
    defparam duty_i7_LC_12_26_7.SEQ_MODE=4'b1000;
    defparam duty_i7_LC_12_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i7_LC_12_26_7 (
            .in0(_gnd_net_),
            .in1(N__49020),
            .in2(N__43404),
            .in3(N__43374),
            .lcout(duty_7),
            .ltout(),
            .carryin(n12465),
            .carryout(n12466),
            .clk(N__55796),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i8_LC_12_27_0.C_ON=1'b1;
    defparam duty_i8_LC_12_27_0.SEQ_MODE=4'b1000;
    defparam duty_i8_LC_12_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i8_LC_12_27_0 (
            .in0(_gnd_net_),
            .in1(N__43371),
            .in2(N__48984),
            .in3(N__43362),
            .lcout(duty_8),
            .ltout(),
            .carryin(bfn_12_27_0_),
            .carryout(n12467),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i9_LC_12_27_1.C_ON=1'b1;
    defparam duty_i9_LC_12_27_1.SEQ_MODE=4'b1000;
    defparam duty_i9_LC_12_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i9_LC_12_27_1 (
            .in0(_gnd_net_),
            .in1(N__43359),
            .in2(N__48945),
            .in3(N__43335),
            .lcout(duty_9),
            .ltout(),
            .carryin(n12467),
            .carryout(n12468),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i10_LC_12_27_2.C_ON=1'b1;
    defparam duty_i10_LC_12_27_2.SEQ_MODE=4'b1000;
    defparam duty_i10_LC_12_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i10_LC_12_27_2 (
            .in0(_gnd_net_),
            .in1(N__43332),
            .in2(N__48900),
            .in3(N__43311),
            .lcout(duty_10),
            .ltout(),
            .carryin(n12468),
            .carryout(n12469),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i11_LC_12_27_3.C_ON=1'b1;
    defparam duty_i11_LC_12_27_3.SEQ_MODE=4'b1000;
    defparam duty_i11_LC_12_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i11_LC_12_27_3 (
            .in0(_gnd_net_),
            .in1(N__43734),
            .in2(N__49488),
            .in3(N__43728),
            .lcout(duty_11),
            .ltout(),
            .carryin(n12469),
            .carryout(n12470),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i12_LC_12_27_4.C_ON=1'b1;
    defparam duty_i12_LC_12_27_4.SEQ_MODE=4'b1000;
    defparam duty_i12_LC_12_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i12_LC_12_27_4 (
            .in0(_gnd_net_),
            .in1(N__43725),
            .in2(N__49443),
            .in3(N__43716),
            .lcout(duty_12),
            .ltout(),
            .carryin(n12470),
            .carryout(n12471),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i13_LC_12_27_5.C_ON=1'b1;
    defparam duty_i13_LC_12_27_5.SEQ_MODE=4'b1000;
    defparam duty_i13_LC_12_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i13_LC_12_27_5 (
            .in0(_gnd_net_),
            .in1(N__43713),
            .in2(N__49392),
            .in3(N__43683),
            .lcout(duty_13),
            .ltout(),
            .carryin(n12471),
            .carryout(n12472),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i14_LC_12_27_6.C_ON=1'b1;
    defparam duty_i14_LC_12_27_6.SEQ_MODE=4'b1000;
    defparam duty_i14_LC_12_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i14_LC_12_27_6 (
            .in0(_gnd_net_),
            .in1(N__43680),
            .in2(N__49344),
            .in3(N__43656),
            .lcout(duty_14),
            .ltout(),
            .carryin(n12472),
            .carryout(n12473),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i15_LC_12_27_7.C_ON=1'b1;
    defparam duty_i15_LC_12_27_7.SEQ_MODE=4'b1000;
    defparam duty_i15_LC_12_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i15_LC_12_27_7 (
            .in0(_gnd_net_),
            .in1(N__54881),
            .in2(N__43653),
            .in3(N__43611),
            .lcout(duty_15),
            .ltout(),
            .carryin(n12473),
            .carryout(n12474),
            .clk(N__55799),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i16_LC_12_28_0.C_ON=1'b1;
    defparam duty_i16_LC_12_28_0.SEQ_MODE=4'b1000;
    defparam duty_i16_LC_12_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i16_LC_12_28_0 (
            .in0(_gnd_net_),
            .in1(N__43608),
            .in2(N__49296),
            .in3(N__43578),
            .lcout(duty_16),
            .ltout(),
            .carryin(bfn_12_28_0_),
            .carryout(n12475),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i17_LC_12_28_1.C_ON=1'b1;
    defparam duty_i17_LC_12_28_1.SEQ_MODE=4'b1000;
    defparam duty_i17_LC_12_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i17_LC_12_28_1 (
            .in0(_gnd_net_),
            .in1(N__43575),
            .in2(N__49257),
            .in3(N__43563),
            .lcout(duty_17),
            .ltout(),
            .carryin(n12475),
            .carryout(n12476),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i18_LC_12_28_2.C_ON=1'b1;
    defparam duty_i18_LC_12_28_2.SEQ_MODE=4'b1000;
    defparam duty_i18_LC_12_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i18_LC_12_28_2 (
            .in0(_gnd_net_),
            .in1(N__43560),
            .in2(N__49215),
            .in3(N__43530),
            .lcout(duty_18),
            .ltout(),
            .carryin(n12476),
            .carryout(n12477),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i19_LC_12_28_3.C_ON=1'b1;
    defparam duty_i19_LC_12_28_3.SEQ_MODE=4'b1000;
    defparam duty_i19_LC_12_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i19_LC_12_28_3 (
            .in0(_gnd_net_),
            .in1(N__43917),
            .in2(N__54810),
            .in3(N__43887),
            .lcout(duty_19),
            .ltout(),
            .carryin(n12477),
            .carryout(n12478),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i20_LC_12_28_4.C_ON=1'b1;
    defparam duty_i20_LC_12_28_4.SEQ_MODE=4'b1000;
    defparam duty_i20_LC_12_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i20_LC_12_28_4 (
            .in0(_gnd_net_),
            .in1(N__49590),
            .in2(N__43884),
            .in3(N__43875),
            .lcout(duty_20),
            .ltout(),
            .carryin(n12478),
            .carryout(n12479),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i21_LC_12_28_5.C_ON=1'b1;
    defparam duty_i21_LC_12_28_5.SEQ_MODE=4'b1000;
    defparam duty_i21_LC_12_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i21_LC_12_28_5 (
            .in0(_gnd_net_),
            .in1(N__43872),
            .in2(N__54852),
            .in3(N__43863),
            .lcout(duty_21),
            .ltout(),
            .carryin(n12479),
            .carryout(n12480),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i22_LC_12_28_6.C_ON=1'b1;
    defparam duty_i22_LC_12_28_6.SEQ_MODE=4'b1000;
    defparam duty_i22_LC_12_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i22_LC_12_28_6 (
            .in0(_gnd_net_),
            .in1(N__43860),
            .in2(N__49548),
            .in3(N__43833),
            .lcout(duty_22),
            .ltout(),
            .carryin(n12480),
            .carryout(n12481),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i23_LC_12_28_7.C_ON=1'b0;
    defparam duty_i23_LC_12_28_7.SEQ_MODE=4'b1000;
    defparam duty_i23_LC_12_28_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 duty_i23_LC_12_28_7 (
            .in0(N__54763),
            .in1(N__43830),
            .in2(_gnd_net_),
            .in3(N__43824),
            .lcout(duty_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55803),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i35_2_lut_LC_12_29_2.C_ON=1'b0;
    defparam LessThan_299_i35_2_lut_LC_12_29_2.SEQ_MODE=4'b0000;
    defparam LessThan_299_i35_2_lut_LC_12_29_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i35_2_lut_LC_12_29_2 (
            .in0(_gnd_net_),
            .in1(N__46558),
            .in2(_gnd_net_),
            .in3(N__43934),
            .lcout(n35),
            .ltout(n35_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12540_4_lut_LC_12_29_3.C_ON=1'b0;
    defparam i12540_4_lut_LC_12_29_3.SEQ_MODE=4'b0000;
    defparam i12540_4_lut_LC_12_29_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12540_4_lut_LC_12_29_3 (
            .in0(N__43806),
            .in1(N__44064),
            .in2(N__43794),
            .in3(N__43791),
            .lcout(n15265),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i27_2_lut_LC_12_29_4.C_ON=1'b0;
    defparam LessThan_299_i27_2_lut_LC_12_29_4.SEQ_MODE=4'b0000;
    defparam LessThan_299_i27_2_lut_LC_12_29_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i27_2_lut_LC_12_29_4 (
            .in0(_gnd_net_),
            .in1(N__43782),
            .in2(_gnd_net_),
            .in3(N__46541),
            .lcout(n27_adj_671),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i12_LC_12_29_5.C_ON=1'b0;
    defparam pwm_setpoint_i12_LC_12_29_5.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i12_LC_12_29_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i12_LC_12_29_5 (
            .in0(N__44093),
            .in1(N__55260),
            .in2(_gnd_net_),
            .in3(N__44076),
            .lcout(pwm_setpoint_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55808),
            .ce(),
            .sr(_gnd_net_));
    defparam i12553_3_lut_LC_12_29_6.C_ON=1'b0;
    defparam i12553_3_lut_LC_12_29_6.SEQ_MODE=4'b0000;
    defparam i12553_3_lut_LC_12_29_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12553_3_lut_LC_12_29_6 (
            .in0(N__44063),
            .in1(N__44055),
            .in2(_gnd_net_),
            .in3(N__44031),
            .lcout(n15278),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12510_3_lut_LC_12_30_1.C_ON=1'b0;
    defparam i12510_3_lut_LC_12_30_1.SEQ_MODE=4'b0000;
    defparam i12510_3_lut_LC_12_30_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12510_3_lut_LC_12_30_1 (
            .in0(N__45270),
            .in1(N__47245),
            .in2(_gnd_net_),
            .in3(N__44022),
            .lcout(),
            .ltout(n15235_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12511_3_lut_LC_12_30_2.C_ON=1'b0;
    defparam i12511_3_lut_LC_12_30_2.SEQ_MODE=4'b0000;
    defparam i12511_3_lut_LC_12_30_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12511_3_lut_LC_12_30_2 (
            .in0(_gnd_net_),
            .in1(N__45471),
            .in2(N__44013),
            .in3(N__47744),
            .lcout(),
            .ltout(n15236_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12455_3_lut_LC_12_30_3.C_ON=1'b0;
    defparam i12455_3_lut_LC_12_30_3.SEQ_MODE=4'b0000;
    defparam i12455_3_lut_LC_12_30_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 i12455_3_lut_LC_12_30_3 (
            .in0(N__45458),
            .in1(_gnd_net_),
            .in2(N__44010),
            .in3(N__47723),
            .lcout(n15180),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i11_LC_12_30_4.C_ON=1'b0;
    defparam pwm_setpoint_i11_LC_12_30_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i11_LC_12_30_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i11_LC_12_30_4 (
            .in0(N__55271),
            .in1(N__44006),
            .in2(_gnd_net_),
            .in3(N__43986),
            .lcout(pwm_setpoint_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55815),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i17_LC_12_30_6.C_ON=1'b0;
    defparam pwm_setpoint_i17_LC_12_30_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i17_LC_12_30_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i17_LC_12_30_6 (
            .in0(N__55272),
            .in1(N__43973),
            .in2(_gnd_net_),
            .in3(N__43953),
            .lcout(pwm_setpoint_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55815),
            .ce(),
            .sr(_gnd_net_));
    defparam i12549_3_lut_LC_12_30_7.C_ON=1'b0;
    defparam i12549_3_lut_LC_12_30_7.SEQ_MODE=4'b0000;
    defparam i12549_3_lut_LC_12_30_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12549_3_lut_LC_12_30_7 (
            .in0(N__45366),
            .in1(N__45348),
            .in2(_gnd_net_),
            .in3(N__43923),
            .lcout(n15274),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i8_3_lut_3_lut_LC_12_31_0.C_ON=1'b0;
    defparam LessThan_299_i8_3_lut_3_lut_LC_12_31_0.SEQ_MODE=4'b0000;
    defparam LessThan_299_i8_3_lut_3_lut_LC_12_31_0.LUT_INIT=16'b1000100011101110;
    LogicCell40 LessThan_299_i8_3_lut_3_lut_LC_12_31_0 (
            .in0(N__47489),
            .in1(N__47364),
            .in2(_gnd_net_),
            .in3(N__47346),
            .lcout(),
            .ltout(n8_adj_657_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12494_4_lut_LC_12_31_1.C_ON=1'b0;
    defparam i12494_4_lut_LC_12_31_1.SEQ_MODE=4'b0000;
    defparam i12494_4_lut_LC_12_31_1.LUT_INIT=16'b1111111000010000;
    LogicCell40 i12494_4_lut_LC_12_31_1 (
            .in0(N__44166),
            .in1(N__45390),
            .in2(N__44208),
            .in3(N__44193),
            .lcout(),
            .ltout(n15219_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12530_4_lut_LC_12_31_2.C_ON=1'b0;
    defparam i12530_4_lut_LC_12_31_2.SEQ_MODE=4'b0000;
    defparam i12530_4_lut_LC_12_31_2.LUT_INIT=16'b1111000011100100;
    LogicCell40 i12530_4_lut_LC_12_31_2 (
            .in0(N__44164),
            .in1(N__44205),
            .in2(N__44196),
            .in3(N__47706),
            .lcout(n15255),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i24_3_lut_LC_12_31_3.C_ON=1'b0;
    defparam LessThan_299_i24_3_lut_LC_12_31_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i24_3_lut_LC_12_31_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 LessThan_299_i24_3_lut_LC_12_31_3 (
            .in0(N__44187),
            .in1(N__44163),
            .in2(_gnd_net_),
            .in3(N__44100),
            .lcout(n24_adj_669),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i45_2_lut_LC_12_31_4.C_ON=1'b0;
    defparam LessThan_299_i45_2_lut_LC_12_31_4.SEQ_MODE=4'b0000;
    defparam LessThan_299_i45_2_lut_LC_12_31_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i45_2_lut_LC_12_31_4 (
            .in0(_gnd_net_),
            .in1(N__44186),
            .in2(_gnd_net_),
            .in3(N__46497),
            .lcout(n45),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12545_3_lut_LC_12_31_5.C_ON=1'b0;
    defparam i12545_3_lut_LC_12_31_5.SEQ_MODE=4'b0000;
    defparam i12545_3_lut_LC_12_31_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12545_3_lut_LC_12_31_5 (
            .in0(N__45444),
            .in1(N__45432),
            .in2(_gnd_net_),
            .in3(N__44172),
            .lcout(),
            .ltout(n40_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12532_4_lut_LC_12_31_6.C_ON=1'b0;
    defparam i12532_4_lut_LC_12_31_6.SEQ_MODE=4'b0000;
    defparam i12532_4_lut_LC_12_31_6.LUT_INIT=16'b1100110011011000;
    LogicCell40 i12532_4_lut_LC_12_31_6 (
            .in0(N__44165),
            .in1(N__44148),
            .in2(N__44142),
            .in3(N__45414),
            .lcout(n15257),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i20_LC_12_32_0.C_ON=1'b0;
    defparam pwm_setpoint_i20_LC_12_32_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i20_LC_12_32_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i20_LC_12_32_0 (
            .in0(N__55309),
            .in1(N__44139),
            .in2(_gnd_net_),
            .in3(N__44121),
            .lcout(pwm_setpoint_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55823),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i22_1_lut_LC_12_32_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i22_1_lut_LC_12_32_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i22_1_lut_LC_12_32_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i22_1_lut_LC_12_32_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44312),
            .lcout(n4_adj_584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i16_3_lut_3_lut_LC_12_32_2.C_ON=1'b0;
    defparam LessThan_299_i16_3_lut_3_lut_LC_12_32_2.SEQ_MODE=4'b0000;
    defparam LessThan_299_i16_3_lut_3_lut_LC_12_32_2.LUT_INIT=16'b1101110101000100;
    LogicCell40 LessThan_299_i16_3_lut_3_lut_LC_12_32_2 (
            .in0(N__47188),
            .in1(N__45379),
            .in2(_gnd_net_),
            .in3(N__47306),
            .lcout(n16_adj_664),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2175_1_lut_LC_12_32_5.C_ON=1'b0;
    defparam i2175_1_lut_LC_12_32_5.SEQ_MODE=4'b0000;
    defparam i2175_1_lut_LC_12_32_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 i2175_1_lut_LC_12_32_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55308),
            .lcout(pwm_setpoint_23__N_195),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_3_lut_LC_12_32_6.C_ON=1'b0;
    defparam i14_3_lut_LC_12_32_6.SEQ_MODE=4'b0000;
    defparam i14_3_lut_LC_12_32_6.LUT_INIT=16'b0101111111111010;
    LogicCell40 i14_3_lut_LC_12_32_6 (
            .in0(N__47633),
            .in1(_gnd_net_),
            .in2(N__47598),
            .in3(N__47672),
            .lcout(n6_adj_717),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i21_LC_12_32_7.C_ON=1'b0;
    defparam pwm_setpoint_i21_LC_12_32_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i21_LC_12_32_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 pwm_setpoint_i21_LC_12_32_7 (
            .in0(N__44322),
            .in1(N__55310),
            .in2(_gnd_net_),
            .in3(N__44313),
            .lcout(pwm_setpoint_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55823),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_13_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_13_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_13_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_2_lut_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(N__45642),
            .in2(_gnd_net_),
            .in3(N__44286),
            .lcout(n1801),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(n12577),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_13_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_13_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_13_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_3_lut_LC_13_17_1 (
            .in0(_gnd_net_),
            .in1(N__52731),
            .in2(N__45665),
            .in3(N__44268),
            .lcout(n1800),
            .ltout(),
            .carryin(n12577),
            .carryout(n12578),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_13_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_13_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_13_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_4_lut_LC_13_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45593),
            .in3(N__44253),
            .lcout(n1799),
            .ltout(),
            .carryin(n12578),
            .carryout(n12579),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_13_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_13_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_13_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_5_lut_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(N__52732),
            .in2(N__45686),
            .in3(N__44241),
            .lcout(n1798),
            .ltout(),
            .carryin(n12579),
            .carryout(n12580),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_13_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_13_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_13_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_6_lut_LC_13_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45536),
            .in3(N__44229),
            .lcout(n1797),
            .ltout(),
            .carryin(n12580),
            .carryout(n12581),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_13_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_13_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_7_lut_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45494),
            .in3(N__44211),
            .lcout(n1796),
            .ltout(),
            .carryin(n12581),
            .carryout(n12582),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_13_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_13_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_8_lut_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(N__52734),
            .in2(N__50105),
            .in3(N__44469),
            .lcout(n1795),
            .ltout(),
            .carryin(n12582),
            .carryout(n12583),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_13_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_13_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_13_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_9_lut_LC_13_17_7 (
            .in0(_gnd_net_),
            .in1(N__52733),
            .in2(N__49791),
            .in3(N__44454),
            .lcout(n1794),
            .ltout(),
            .carryin(n12583),
            .carryout(n12584),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_13_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_13_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_13_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_10_lut_LC_13_18_0 (
            .in0(_gnd_net_),
            .in1(N__52724),
            .in2(N__50339),
            .in3(N__44442),
            .lcout(n1793),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(n12585),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_13_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_13_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_13_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_11_lut_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(N__53085),
            .in2(N__50285),
            .in3(N__44427),
            .lcout(n1792),
            .ltout(),
            .carryin(n12585),
            .carryout(n12586),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_13_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_13_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_13_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_12_lut_LC_13_18_2 (
            .in0(_gnd_net_),
            .in1(N__52725),
            .in2(N__50312),
            .in3(N__44415),
            .lcout(n1791),
            .ltout(),
            .carryin(n12586),
            .carryout(n12587),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_13_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_13_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_13_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_13_lut_LC_13_18_3 (
            .in0(_gnd_net_),
            .in1(N__53086),
            .in2(N__50249),
            .in3(N__44400),
            .lcout(n1790),
            .ltout(),
            .carryin(n12587),
            .carryout(n12588),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_13_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_13_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_13_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_14_lut_LC_13_18_4 (
            .in0(_gnd_net_),
            .in1(N__52726),
            .in2(N__44397),
            .in3(N__44376),
            .lcout(n1789),
            .ltout(),
            .carryin(n12588),
            .carryout(n12589),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_13_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_13_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_13_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_15_lut_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(N__44372),
            .in2(N__53002),
            .in3(N__44343),
            .lcout(n1788),
            .ltout(),
            .carryin(n12589),
            .carryout(n12590),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_13_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_13_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_13_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_16_lut_LC_13_18_6 (
            .in0(_gnd_net_),
            .in1(N__44579),
            .in2(N__53449),
            .in3(N__44553),
            .lcout(n1787),
            .ltout(),
            .carryin(n12590),
            .carryout(n12591),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_13_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_13_18_7.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1168_17_lut_LC_13_18_7 (
            .in0(N__52730),
            .in1(N__44543),
            .in2(N__47943),
            .in3(N__44526),
            .lcout(n1818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_13_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_13_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_13_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_2_lut_LC_13_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48223),
            .in3(N__44499),
            .lcout(n1601),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(n12550),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_13_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_13_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_13_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_3_lut_LC_13_19_1 (
            .in0(_gnd_net_),
            .in1(N__52721),
            .in2(N__45762),
            .in3(N__44496),
            .lcout(n1600),
            .ltout(),
            .carryin(n12550),
            .carryout(n12551),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_13_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_13_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_13_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_4_lut_LC_13_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48168),
            .in3(N__44493),
            .lcout(n1599),
            .ltout(),
            .carryin(n12551),
            .carryout(n12552),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_13_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_13_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_13_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_5_lut_LC_13_19_3 (
            .in0(_gnd_net_),
            .in1(N__52722),
            .in2(N__45557),
            .in3(N__44490),
            .lcout(n1598),
            .ltout(),
            .carryin(n12552),
            .carryout(n12553),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_13_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_13_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_13_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_6_lut_LC_13_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50580),
            .in3(N__44487),
            .lcout(n1597),
            .ltout(),
            .carryin(n12553),
            .carryout(n12554),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_13_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_13_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_13_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_7_lut_LC_13_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50751),
            .in3(N__44484),
            .lcout(n1596),
            .ltout(),
            .carryin(n12554),
            .carryout(n12555),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_13_19_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_13_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_13_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_8_lut_LC_13_19_6 (
            .in0(_gnd_net_),
            .in1(N__52786),
            .in2(N__49987),
            .in3(N__44481),
            .lcout(n1595),
            .ltout(),
            .carryin(n12555),
            .carryout(n12556),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_13_19_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_13_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_13_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_9_lut_LC_13_19_7 (
            .in0(_gnd_net_),
            .in1(N__52723),
            .in2(N__50798),
            .in3(N__44649),
            .lcout(n1594),
            .ltout(),
            .carryin(n12556),
            .carryout(n12557),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_13_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_13_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_13_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_10_lut_LC_13_20_0 (
            .in0(_gnd_net_),
            .in1(N__52711),
            .in2(N__50052),
            .in3(N__44646),
            .lcout(n1593),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(n12558),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_13_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_13_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_13_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_11_lut_LC_13_20_1 (
            .in0(_gnd_net_),
            .in1(N__52713),
            .in2(N__48444),
            .in3(N__44643),
            .lcout(n1592),
            .ltout(),
            .carryin(n12558),
            .carryout(n12559),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_13_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_13_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_13_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_12_lut_LC_13_20_2 (
            .in0(_gnd_net_),
            .in1(N__48416),
            .in2(N__53000),
            .in3(N__44634),
            .lcout(n1591),
            .ltout(),
            .carryin(n12559),
            .carryout(n12560),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_13_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_13_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_13_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_13_lut_LC_13_20_3 (
            .in0(_gnd_net_),
            .in1(N__52717),
            .in2(N__47916),
            .in3(N__44631),
            .lcout(n1590),
            .ltout(),
            .carryin(n12560),
            .carryout(n12561),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_13_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_13_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_13_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_14_lut_LC_13_20_4 (
            .in0(_gnd_net_),
            .in1(N__48263),
            .in2(N__53001),
            .in3(N__44628),
            .lcout(n1589),
            .ltout(),
            .carryin(n12561),
            .carryout(n12562),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_13_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_13_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_13_20_5.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1034_15_lut_LC_13_20_5 (
            .in0(N__52712),
            .in1(N__45725),
            .in2(N__50820),
            .in3(N__44625),
            .lcout(n1620_adj_607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i843_3_lut_LC_13_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i843_3_lut_LC_13_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i843_3_lut_LC_13_21_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i843_3_lut_LC_13_21_1 (
            .in0(_gnd_net_),
            .in1(N__48606),
            .in2(N__48627),
            .in3(N__51590),
            .lcout(n1331),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_13_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_13_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_13_21_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i21_3_lut_LC_13_21_2 (
            .in0(N__44622),
            .in1(N__46189),
            .in2(_gnd_net_),
            .in3(N__44610),
            .lcout(n299),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_13_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_13_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_13_21_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i7_3_lut_LC_13_21_3 (
            .in0(N__46190),
            .in1(N__44904),
            .in2(_gnd_net_),
            .in3(N__44895),
            .lcout(n313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_13_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_13_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_13_21_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i23_3_lut_LC_13_21_4 (
            .in0(N__44805),
            .in1(N__44817),
            .in2(_gnd_net_),
            .in3(N__46188),
            .lcout(n297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_21_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44804),
            .lcout(n11_adj_632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_13_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_13_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_13_21_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i25_3_lut_LC_13_21_6 (
            .in0(N__44730),
            .in1(N__44769),
            .in2(_gnd_net_),
            .in3(N__46187),
            .lcout(n295),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_13_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_13_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_13_21_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_13_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44729),
            .lcout(n9_adj_630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i640_3_lut_LC_13_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i640_3_lut_LC_13_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i640_3_lut_LC_13_22_0.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i640_3_lut_LC_13_22_0 (
            .in0(N__44691),
            .in1(_gnd_net_),
            .in2(N__44664),
            .in3(N__44956),
            .lcout(n1032),
            .ltout(n1032_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9947_3_lut_LC_13_22_1.C_ON=1'b0;
    defparam i9947_3_lut_LC_13_22_1.SEQ_MODE=4'b0000;
    defparam i9947_3_lut_LC_13_22_1.LUT_INIT=16'b1111000010100000;
    LogicCell40 i9947_3_lut_LC_13_22_1 (
            .in0(N__46266),
            .in1(_gnd_net_),
            .in2(N__44655),
            .in3(N__45934),
            .lcout(),
            .ltout(n11914_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_170_LC_13_22_2.C_ON=1'b0;
    defparam i1_4_lut_adj_170_LC_13_22_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_170_LC_13_22_2.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_170_LC_13_22_2 (
            .in0(N__45133),
            .in1(N__45025),
            .in2(N__44652),
            .in3(N__45874),
            .lcout(),
            .ltout(n13716_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12777_4_lut_LC_13_22_3.C_ON=1'b0;
    defparam i12777_4_lut_LC_13_22_3.SEQ_MODE=4'b0000;
    defparam i12777_4_lut_LC_13_22_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12777_4_lut_LC_13_22_3 (
            .in0(N__45107),
            .in1(N__45047),
            .in2(N__45000),
            .in3(N__45082),
            .lcout(n1059),
            .ltout(n1059_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i702_3_lut_LC_13_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i702_3_lut_LC_13_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i702_3_lut_LC_13_22_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i702_3_lut_LC_13_22_4 (
            .in0(N__45083),
            .in1(_gnd_net_),
            .in2(N__44997),
            .in3(N__45069),
            .lcout(n1126),
            .ltout(n1126_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_171_LC_13_22_5.C_ON=1'b0;
    defparam i1_3_lut_adj_171_LC_13_22_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_171_LC_13_22_5.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_171_LC_13_22_5 (
            .in0(_gnd_net_),
            .in1(N__51787),
            .in2(N__44994),
            .in3(N__51748),
            .lcout(n14428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i704_3_lut_LC_13_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i704_3_lut_LC_13_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i704_3_lut_LC_13_22_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i704_3_lut_LC_13_22_6 (
            .in0(_gnd_net_),
            .in1(N__45120),
            .in2(N__45140),
            .in3(N__46409),
            .lcout(n1128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i635_rep_55_3_lut_LC_13_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i635_rep_55_3_lut_LC_13_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i635_rep_55_3_lut_LC_13_22_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i635_rep_55_3_lut_LC_13_22_7 (
            .in0(N__44991),
            .in1(_gnd_net_),
            .in2(N__44963),
            .in3(N__44925),
            .lcout(n1027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_13_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_13_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_13_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_2_lut_LC_13_23_0 (
            .in0(_gnd_net_),
            .in1(N__46264),
            .in2(_gnd_net_),
            .in3(N__44919),
            .lcout(n1101),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(n12500),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_13_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_13_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_13_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_3_lut_LC_13_23_1 (
            .in0(_gnd_net_),
            .in1(N__52557),
            .in2(N__45941),
            .in3(N__44916),
            .lcout(n1100),
            .ltout(),
            .carryin(n12500),
            .carryout(n12501),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_13_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_13_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_13_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_4_lut_LC_13_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45915),
            .in3(N__44913),
            .lcout(n1099),
            .ltout(),
            .carryin(n12501),
            .carryout(n12502),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_13_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_13_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_13_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_5_lut_LC_13_23_3 (
            .in0(_gnd_net_),
            .in1(N__52558),
            .in2(N__45875),
            .in3(N__44910),
            .lcout(n1098),
            .ltout(),
            .carryin(n12502),
            .carryout(n12503),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_13_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_13_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_13_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_6_lut_LC_13_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45030),
            .in3(N__44907),
            .lcout(n1097),
            .ltout(),
            .carryin(n12503),
            .carryout(n12504),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_13_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_13_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_13_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_7_lut_LC_13_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45141),
            .in3(N__45114),
            .lcout(n1096),
            .ltout(),
            .carryin(n12504),
            .carryout(n12505),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_13_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_13_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_13_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_8_lut_LC_13_23_6 (
            .in0(_gnd_net_),
            .in1(N__52590),
            .in2(N__45111),
            .in3(N__45090),
            .lcout(n1095),
            .ltout(),
            .carryin(n12505),
            .carryout(n12506),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_13_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_13_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_13_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_9_lut_LC_13_23_7 (
            .in0(_gnd_net_),
            .in1(N__52559),
            .in2(N__45087),
            .in3(N__45063),
            .lcout(n1094),
            .ltout(),
            .carryin(n12506),
            .carryout(n12507),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_13_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_13_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_13_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_10_lut_LC_13_24_0 (
            .in0(_gnd_net_),
            .in1(N__52429),
            .in2(N__45057),
            .in3(N__45060),
            .lcout(n1093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i701_3_lut_LC_13_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i701_3_lut_LC_13_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i701_3_lut_LC_13_24_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i701_3_lut_LC_13_24_1 (
            .in0(_gnd_net_),
            .in1(N__45056),
            .in2(N__46424),
            .in3(N__45036),
            .lcout(n1125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i705_3_lut_LC_13_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i705_3_lut_LC_13_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i705_3_lut_LC_13_24_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i705_3_lut_LC_13_24_6 (
            .in0(_gnd_net_),
            .in1(N__45029),
            .in2(N__45009),
            .in3(N__46414),
            .lcout(n1129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_13_25_0.C_ON=1'b0;
    defparam i9_4_lut_LC_13_25_0.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_13_25_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i9_4_lut_LC_13_25_0 (
            .in0(N__49211),
            .in1(N__49388),
            .in2(N__49442),
            .in3(N__49340),
            .lcout(n23_adj_700),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_25_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_25_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_25_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.pwm_counter_661__i0_LC_13_26_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i0_LC_13_26_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i0_LC_13_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i0_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__45197),
            .in2(_gnd_net_),
            .in3(N__45183),
            .lcout(pwm_counter_0),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\PWM.n13056 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i1_LC_13_26_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i1_LC_13_26_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i1_LC_13_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i1_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__45179),
            .in2(_gnd_net_),
            .in3(N__45165),
            .lcout(pwm_counter_1),
            .ltout(),
            .carryin(\PWM.n13056 ),
            .carryout(\PWM.n13057 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i2_LC_13_26_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i2_LC_13_26_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i2_LC_13_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i2_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__46811),
            .in2(_gnd_net_),
            .in3(N__45162),
            .lcout(pwm_counter_2),
            .ltout(),
            .carryin(\PWM.n13057 ),
            .carryout(\PWM.n13058 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i3_LC_13_26_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i3_LC_13_26_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i3_LC_13_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i3_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__46793),
            .in2(_gnd_net_),
            .in3(N__45159),
            .lcout(pwm_counter_3),
            .ltout(),
            .carryin(\PWM.n13058 ),
            .carryout(\PWM.n13059 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i4_LC_13_26_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i4_LC_13_26_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i4_LC_13_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i4_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__47468),
            .in2(_gnd_net_),
            .in3(N__45156),
            .lcout(pwm_counter_4),
            .ltout(),
            .carryin(\PWM.n13059 ),
            .carryout(\PWM.n13060 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i5_LC_13_26_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i5_LC_13_26_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i5_LC_13_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i5_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(N__46772),
            .in2(_gnd_net_),
            .in3(N__45153),
            .lcout(pwm_counter_5),
            .ltout(),
            .carryin(\PWM.n13060 ),
            .carryout(\PWM.n13061 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i6_LC_13_26_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i6_LC_13_26_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i6_LC_13_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i6_LC_13_26_6  (
            .in0(_gnd_net_),
            .in1(N__46708),
            .in2(_gnd_net_),
            .in3(N__45150),
            .lcout(pwm_counter_6),
            .ltout(),
            .carryin(\PWM.n13061 ),
            .carryout(\PWM.n13062 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i7_LC_13_26_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i7_LC_13_26_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i7_LC_13_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i7_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(N__46741),
            .in2(_gnd_net_),
            .in3(N__45147),
            .lcout(pwm_counter_7),
            .ltout(),
            .carryin(\PWM.n13062 ),
            .carryout(\PWM.n13063 ),
            .clk(N__55800),
            .ce(),
            .sr(N__47118));
    defparam \PWM.pwm_counter_661__i8_LC_13_27_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i8_LC_13_27_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i8_LC_13_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i8_LC_13_27_0  (
            .in0(_gnd_net_),
            .in1(N__47338),
            .in2(_gnd_net_),
            .in3(N__45144),
            .lcout(pwm_counter_8),
            .ltout(),
            .carryin(bfn_13_27_0_),
            .carryout(\PWM.n13064 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i9_LC_13_27_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i9_LC_13_27_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i9_LC_13_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i9_LC_13_27_1  (
            .in0(_gnd_net_),
            .in1(N__47269),
            .in2(_gnd_net_),
            .in3(N__45228),
            .lcout(pwm_counter_9),
            .ltout(),
            .carryin(\PWM.n13064 ),
            .carryout(\PWM.n13065 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i10_LC_13_27_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i10_LC_13_27_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i10_LC_13_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i10_LC_13_27_2  (
            .in0(_gnd_net_),
            .in1(N__46658),
            .in2(_gnd_net_),
            .in3(N__45225),
            .lcout(pwm_counter_10),
            .ltout(),
            .carryin(\PWM.n13065 ),
            .carryout(\PWM.n13066 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i11_LC_13_27_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i11_LC_13_27_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i11_LC_13_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i11_LC_13_27_3  (
            .in0(_gnd_net_),
            .in1(N__46679),
            .in2(_gnd_net_),
            .in3(N__45222),
            .lcout(pwm_counter_11),
            .ltout(),
            .carryin(\PWM.n13066 ),
            .carryout(\PWM.n13067 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i12_LC_13_27_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i12_LC_13_27_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i12_LC_13_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i12_LC_13_27_4  (
            .in0(_gnd_net_),
            .in1(N__47155),
            .in2(_gnd_net_),
            .in3(N__45219),
            .lcout(pwm_counter_12),
            .ltout(),
            .carryin(\PWM.n13067 ),
            .carryout(\PWM.n13068 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i13_LC_13_27_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i13_LC_13_27_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i13_LC_13_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i13_LC_13_27_5  (
            .in0(_gnd_net_),
            .in1(N__46537),
            .in2(_gnd_net_),
            .in3(N__45216),
            .lcout(pwm_counter_13),
            .ltout(),
            .carryin(\PWM.n13068 ),
            .carryout(\PWM.n13069 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i14_LC_13_27_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i14_LC_13_27_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i14_LC_13_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i14_LC_13_27_6  (
            .in0(_gnd_net_),
            .in1(N__46633),
            .in2(_gnd_net_),
            .in3(N__45213),
            .lcout(pwm_counter_14),
            .ltout(),
            .carryin(\PWM.n13069 ),
            .carryout(\PWM.n13070 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i15_LC_13_27_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i15_LC_13_27_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i15_LC_13_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i15_LC_13_27_7  (
            .in0(_gnd_net_),
            .in1(N__46444),
            .in2(_gnd_net_),
            .in3(N__45210),
            .lcout(pwm_counter_15),
            .ltout(),
            .carryin(\PWM.n13070 ),
            .carryout(\PWM.n13071 ),
            .clk(N__55804),
            .ce(),
            .sr(N__47110));
    defparam \PWM.pwm_counter_661__i16_LC_13_28_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i16_LC_13_28_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i16_LC_13_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i16_LC_13_28_0  (
            .in0(_gnd_net_),
            .in1(N__46590),
            .in2(_gnd_net_),
            .in3(N__45207),
            .lcout(pwm_counter_16),
            .ltout(),
            .carryin(bfn_13_28_0_),
            .carryout(\PWM.n13072 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i17_LC_13_28_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i17_LC_13_28_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i17_LC_13_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i17_LC_13_28_1  (
            .in0(_gnd_net_),
            .in1(N__46560),
            .in2(_gnd_net_),
            .in3(N__45204),
            .lcout(pwm_counter_17),
            .ltout(),
            .carryin(\PWM.n13072 ),
            .carryout(\PWM.n13073 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i18_LC_13_28_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i18_LC_13_28_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i18_LC_13_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i18_LC_13_28_2  (
            .in0(_gnd_net_),
            .in1(N__46475),
            .in2(_gnd_net_),
            .in3(N__45255),
            .lcout(pwm_counter_18),
            .ltout(),
            .carryin(\PWM.n13073 ),
            .carryout(\PWM.n13074 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i19_LC_13_28_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i19_LC_13_28_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i19_LC_13_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i19_LC_13_28_3  (
            .in0(_gnd_net_),
            .in1(N__47087),
            .in2(_gnd_net_),
            .in3(N__45252),
            .lcout(pwm_counter_19),
            .ltout(),
            .carryin(\PWM.n13074 ),
            .carryout(\PWM.n13075 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i20_LC_13_28_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i20_LC_13_28_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i20_LC_13_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i20_LC_13_28_4  (
            .in0(_gnd_net_),
            .in1(N__46613),
            .in2(_gnd_net_),
            .in3(N__45249),
            .lcout(pwm_counter_20),
            .ltout(),
            .carryin(\PWM.n13075 ),
            .carryout(\PWM.n13076 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i21_LC_13_28_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i21_LC_13_28_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i21_LC_13_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i21_LC_13_28_5  (
            .in0(_gnd_net_),
            .in1(N__47179),
            .in2(_gnd_net_),
            .in3(N__45246),
            .lcout(pwm_counter_21),
            .ltout(),
            .carryin(\PWM.n13076 ),
            .carryout(\PWM.n13077 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i22_LC_13_28_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i22_LC_13_28_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i22_LC_13_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i22_LC_13_28_6  (
            .in0(_gnd_net_),
            .in1(N__46496),
            .in2(_gnd_net_),
            .in3(N__45243),
            .lcout(pwm_counter_22),
            .ltout(),
            .carryin(\PWM.n13077 ),
            .carryout(\PWM.n13078 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i23_LC_13_28_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i23_LC_13_28_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i23_LC_13_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i23_LC_13_28_7  (
            .in0(_gnd_net_),
            .in1(N__46514),
            .in2(_gnd_net_),
            .in3(N__45240),
            .lcout(pwm_counter_23),
            .ltout(),
            .carryin(\PWM.n13078 ),
            .carryout(\PWM.n13079 ),
            .clk(N__55809),
            .ce(),
            .sr(N__47109));
    defparam \PWM.pwm_counter_661__i24_LC_13_29_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i24_LC_13_29_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i24_LC_13_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i24_LC_13_29_0  (
            .in0(_gnd_net_),
            .in1(N__47052),
            .in2(_gnd_net_),
            .in3(N__45237),
            .lcout(pwm_counter_24),
            .ltout(),
            .carryin(bfn_13_29_0_),
            .carryout(\PWM.n13080 ),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam \PWM.pwm_counter_661__i25_LC_13_29_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i25_LC_13_29_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i25_LC_13_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i25_LC_13_29_1  (
            .in0(_gnd_net_),
            .in1(N__46989),
            .in2(_gnd_net_),
            .in3(N__45234),
            .lcout(pwm_counter_25),
            .ltout(),
            .carryin(\PWM.n13080 ),
            .carryout(\PWM.n13081 ),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam \PWM.pwm_counter_661__i26_LC_13_29_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i26_LC_13_29_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i26_LC_13_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i26_LC_13_29_2  (
            .in0(_gnd_net_),
            .in1(N__47013),
            .in2(_gnd_net_),
            .in3(N__45231),
            .lcout(pwm_counter_26),
            .ltout(),
            .carryin(\PWM.n13081 ),
            .carryout(\PWM.n13082 ),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam \PWM.pwm_counter_661__i27_LC_13_29_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i27_LC_13_29_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i27_LC_13_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i27_LC_13_29_3  (
            .in0(_gnd_net_),
            .in1(N__47027),
            .in2(_gnd_net_),
            .in3(N__45333),
            .lcout(pwm_counter_27),
            .ltout(),
            .carryin(\PWM.n13082 ),
            .carryout(\PWM.n13083 ),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam \PWM.pwm_counter_661__i28_LC_13_29_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i28_LC_13_29_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i28_LC_13_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i28_LC_13_29_4  (
            .in0(_gnd_net_),
            .in1(N__46974),
            .in2(_gnd_net_),
            .in3(N__45330),
            .lcout(pwm_counter_28),
            .ltout(),
            .carryin(\PWM.n13083 ),
            .carryout(\PWM.n13084 ),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam \PWM.pwm_counter_661__i29_LC_13_29_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i29_LC_13_29_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i29_LC_13_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i29_LC_13_29_5  (
            .in0(_gnd_net_),
            .in1(N__47040),
            .in2(_gnd_net_),
            .in3(N__45327),
            .lcout(pwm_counter_29),
            .ltout(),
            .carryin(\PWM.n13084 ),
            .carryout(\PWM.n13085 ),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam \PWM.pwm_counter_661__i30_LC_13_29_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_661__i30_LC_13_29_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i30_LC_13_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i30_LC_13_29_6  (
            .in0(_gnd_net_),
            .in1(N__47001),
            .in2(_gnd_net_),
            .in3(N__45324),
            .lcout(pwm_counter_30),
            .ltout(),
            .carryin(\PWM.n13085 ),
            .carryout(\PWM.n13086 ),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam \PWM.pwm_counter_661__i31_LC_13_29_7 .C_ON=1'b0;
    defparam \PWM.pwm_counter_661__i31_LC_13_29_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_661__i31_LC_13_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_661__i31_LC_13_29_7  (
            .in0(_gnd_net_),
            .in1(N__46953),
            .in2(_gnd_net_),
            .in3(N__45321),
            .lcout(pwm_counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55816),
            .ce(),
            .sr(N__47111));
    defparam commutation_state_i0_LC_13_30_0.C_ON=1'b0;
    defparam commutation_state_i0_LC_13_30_0.SEQ_MODE=4'b1001;
    defparam commutation_state_i0_LC_13_30_0.LUT_INIT=16'b0000000001100110;
    LogicCell40 commutation_state_i0_LC_13_30_0 (
            .in0(N__47637),
            .in1(N__47597),
            .in2(_gnd_net_),
            .in3(N__47690),
            .lcout(commutation_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55819),
            .ce(N__45318),
            .sr(N__47697));
    defparam LessThan_299_i11_2_lut_LC_13_30_2.C_ON=1'b0;
    defparam LessThan_299_i11_2_lut_LC_13_30_2.SEQ_MODE=4'b0000;
    defparam LessThan_299_i11_2_lut_LC_13_30_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i11_2_lut_LC_13_30_2 (
            .in0(_gnd_net_),
            .in1(N__45302),
            .in2(_gnd_net_),
            .in3(N__46773),
            .lcout(n11_adj_660),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i13_2_lut_LC_13_30_3.C_ON=1'b0;
    defparam LessThan_299_i13_2_lut_LC_13_30_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i13_2_lut_LC_13_30_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i13_2_lut_LC_13_30_3 (
            .in0(_gnd_net_),
            .in1(N__45285),
            .in2(_gnd_net_),
            .in3(N__46709),
            .lcout(n13_adj_662),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i21_2_lut_LC_13_30_4.C_ON=1'b0;
    defparam LessThan_299_i21_2_lut_LC_13_30_4.SEQ_MODE=4'b0000;
    defparam LessThan_299_i21_2_lut_LC_13_30_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i21_2_lut_LC_13_30_4 (
            .in0(_gnd_net_),
            .in1(N__45269),
            .in2(_gnd_net_),
            .in3(N__46659),
            .lcout(n21_adj_667),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i23_2_lut_LC_13_30_5.C_ON=1'b0;
    defparam LessThan_299_i23_2_lut_LC_13_30_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i23_2_lut_LC_13_30_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i23_2_lut_LC_13_30_5 (
            .in0(N__46680),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45470),
            .lcout(n23_adj_668),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i25_2_lut_LC_13_30_6.C_ON=1'b0;
    defparam LessThan_299_i25_2_lut_LC_13_30_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i25_2_lut_LC_13_30_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i25_2_lut_LC_13_30_6 (
            .in0(_gnd_net_),
            .in1(N__45459),
            .in2(_gnd_net_),
            .in3(N__47157),
            .lcout(n25_adj_670),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i41_2_lut_LC_13_31_1.C_ON=1'b0;
    defparam LessThan_299_i41_2_lut_LC_13_31_1.SEQ_MODE=4'b0000;
    defparam LessThan_299_i41_2_lut_LC_13_31_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i41_2_lut_LC_13_31_1 (
            .in0(_gnd_net_),
            .in1(N__45443),
            .in2(_gnd_net_),
            .in3(N__46614),
            .lcout(n41),
            .ltout(n41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12387_4_lut_LC_13_31_2.C_ON=1'b0;
    defparam i12387_4_lut_LC_13_31_2.SEQ_MODE=4'b0000;
    defparam i12387_4_lut_LC_13_31_2.LUT_INIT=16'b1010101010101011;
    LogicCell40 i12387_4_lut_LC_13_31_2 (
            .in0(N__47757),
            .in1(N__45347),
            .in2(N__45426),
            .in3(N__45423),
            .lcout(n15112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.pwm_out_12_LC_13_31_6 .C_ON=1'b0;
    defparam \PWM.pwm_out_12_LC_13_31_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_out_12_LC_13_31_6 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \PWM.pwm_out_12_LC_13_31_6  (
            .in0(N__46518),
            .in1(N__45408),
            .in2(_gnd_net_),
            .in3(N__45396),
            .lcout(pwm_out),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55824),
            .ce(),
            .sr(N__46935));
    defparam i12383_2_lut_4_lut_LC_13_32_1.C_ON=1'b0;
    defparam i12383_2_lut_4_lut_LC_13_32_1.SEQ_MODE=4'b0000;
    defparam i12383_2_lut_4_lut_LC_13_32_1.LUT_INIT=16'b0111101111011110;
    LogicCell40 i12383_2_lut_4_lut_LC_13_32_1 (
            .in0(N__47277),
            .in1(N__45381),
            .in2(N__47310),
            .in3(N__47190),
            .lcout(n15108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i43_2_lut_LC_13_32_3.C_ON=1'b0;
    defparam LessThan_299_i43_2_lut_LC_13_32_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i43_2_lut_LC_13_32_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i43_2_lut_LC_13_32_3 (
            .in0(_gnd_net_),
            .in1(N__47189),
            .in2(_gnd_net_),
            .in3(N__45380),
            .lcout(n43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i39_2_lut_LC_13_32_5.C_ON=1'b0;
    defparam LessThan_299_i39_2_lut_LC_13_32_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i39_2_lut_LC_13_32_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i39_2_lut_LC_13_32_5 (
            .in0(N__45365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47088),
            .lcout(n39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12878_1_lut_LC_14_17_0.C_ON=1'b0;
    defparam i12878_1_lut_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam i12878_1_lut_LC_14_17_0.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12878_1_lut_LC_14_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50170),
            .in3(_gnd_net_),
            .lcout(n15603),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1043_rep_35_3_lut_LC_14_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1043_rep_35_3_lut_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1043_rep_35_3_lut_LC_14_17_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1043_rep_35_3_lut_LC_14_17_1 (
            .in0(_gnd_net_),
            .in1(N__47802),
            .in2(N__49955),
            .in3(N__50144),
            .lcout(),
            .ltout(n14910_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12442_3_lut_4_lut_LC_14_17_2.C_ON=1'b0;
    defparam i12442_3_lut_4_lut_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam i12442_3_lut_4_lut_LC_14_17_2.LUT_INIT=16'b1101100011110000;
    LogicCell40 i12442_3_lut_4_lut_LC_14_17_2 (
            .in0(N__50145),
            .in1(N__49991),
            .in2(N__45540),
            .in3(N__50668),
            .lcout(n1726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_14_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_14_17_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1107_3_lut_LC_14_17_3 (
            .in0(N__47787),
            .in1(_gnd_net_),
            .in2(N__47769),
            .in3(N__50146),
            .lcout(n1723),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_14_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_14_17_4.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1114_3_lut_LC_14_17_4 (
            .in0(N__47841),
            .in1(_gnd_net_),
            .in2(N__50169),
            .in3(N__47861),
            .lcout(n1730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_76_LC_14_17_5.C_ON=1'b0;
    defparam i1_4_lut_adj_76_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_76_LC_14_17_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_76_LC_14_17_5 (
            .in0(N__47786),
            .in1(N__45702),
            .in2(N__48125),
            .in3(N__50079),
            .lcout(),
            .ltout(n14514_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12881_4_lut_LC_14_17_6.C_ON=1'b0;
    defparam i12881_4_lut_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam i12881_4_lut_LC_14_17_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12881_4_lut_LC_14_17_6 (
            .in0(N__48026),
            .in1(N__48070),
            .in2(N__45510),
            .in3(N__47963),
            .lcout(n1653),
            .ltout(n1653_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_14_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_14_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_14_17_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1117_3_lut_LC_14_17_7 (
            .in0(_gnd_net_),
            .in1(N__47511),
            .in2(N__45507),
            .in3(N__47544),
            .lcout(n1733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_14_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_14_18_0.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1046_3_lut_LC_14_18_0 (
            .in0(N__45504),
            .in1(_gnd_net_),
            .in2(N__45558),
            .in3(N__50653),
            .lcout(n1630_adj_617),
            .ltout(n1630_adj_617_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_14_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_14_18_1.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1113_3_lut_LC_14_18_1 (
            .in0(N__50167),
            .in1(N__47817),
            .in2(N__45498),
            .in3(_gnd_net_),
            .lcout(n1729),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9935_3_lut_LC_14_18_2.C_ON=1'b0;
    defparam i9935_3_lut_LC_14_18_2.SEQ_MODE=4'b0000;
    defparam i9935_3_lut_LC_14_18_2.LUT_INIT=16'b1110111000000000;
    LogicCell40 i9935_3_lut_LC_14_18_2 (
            .in0(N__47542),
            .in1(N__48181),
            .in2(_gnd_net_),
            .in3(N__47884),
            .lcout(),
            .ltout(n11902_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_75_LC_14_18_3.C_ON=1'b0;
    defparam i1_4_lut_adj_75_LC_14_18_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_75_LC_14_18_3.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_75_LC_14_18_3 (
            .in0(N__47857),
            .in1(N__47828),
            .in2(N__45705),
            .in3(N__50554),
            .lcout(n13736),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_14_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_14_18_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1047_3_lut_LC_14_18_4 (
            .in0(_gnd_net_),
            .in1(N__45696),
            .in2(N__48167),
            .in3(N__50652),
            .lcout(n1631_adj_618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_14_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_14_18_5.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1115_3_lut_LC_14_18_5 (
            .in0(N__50168),
            .in1(N__47871),
            .in2(N__47891),
            .in3(_gnd_net_),
            .lcout(n1731),
            .ltout(n1731_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10002_4_lut_LC_14_18_6.C_ON=1'b0;
    defparam i10002_4_lut_LC_14_18_6.SEQ_MODE=4'b0000;
    defparam i10002_4_lut_LC_14_18_6.LUT_INIT=16'b1111111011110000;
    LogicCell40 i10002_4_lut_LC_14_18_6 (
            .in0(N__45658),
            .in1(N__45641),
            .in2(N__45612),
            .in3(N__45586),
            .lcout(n11970),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_14_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_14_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_14_18_7.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1116_3_lut_LC_14_18_7 (
            .in0(N__50166),
            .in1(N__47499),
            .in2(N__48188),
            .in3(_gnd_net_),
            .lcout(n1732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_14_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_14_19_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1038_3_lut_LC_14_19_0 (
            .in0(_gnd_net_),
            .in1(N__47909),
            .in2(N__50662),
            .in3(N__45570),
            .lcout(n1622_adj_609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i976_3_lut_LC_14_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i976_3_lut_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i976_3_lut_LC_14_19_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i976_3_lut_LC_14_19_1 (
            .in0(_gnd_net_),
            .in1(N__51056),
            .in2(N__51400),
            .in3(N__51036),
            .lcout(n1528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_14_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_14_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_14_19_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1037_3_lut_LC_14_19_2 (
            .in0(_gnd_net_),
            .in1(N__45564),
            .in2(N__50661),
            .in3(N__48264),
            .lcout(n1621_adj_608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i979_3_lut_LC_14_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i979_3_lut_LC_14_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i979_3_lut_LC_14_19_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 encoder0_position_31__I_0_i979_3_lut_LC_14_19_3 (
            .in0(N__51387),
            .in1(N__50427),
            .in2(_gnd_net_),
            .in3(N__50453),
            .lcout(n1531),
            .ltout(n1531_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10006_4_lut_LC_14_19_4.C_ON=1'b0;
    defparam i10006_4_lut_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam i10006_4_lut_LC_14_19_4.LUT_INIT=16'b1111111011110000;
    LogicCell40 i10006_4_lut_LC_14_19_4 (
            .in0(N__48224),
            .in1(N__45761),
            .in2(N__45774),
            .in3(N__48160),
            .lcout(n11974),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_14_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_14_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_14_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1040_3_lut_LC_14_19_5 (
            .in0(_gnd_net_),
            .in1(N__48440),
            .in2(N__45771),
            .in3(N__50633),
            .lcout(n1624_adj_611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i981_3_lut_LC_14_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i981_3_lut_LC_14_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i981_3_lut_LC_14_19_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i981_3_lut_LC_14_19_6 (
            .in0(N__50529),
            .in1(N__50502),
            .in2(_gnd_net_),
            .in3(N__51386),
            .lcout(n1533),
            .ltout(n1533_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_14_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_14_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_14_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1048_3_lut_LC_14_19_7 (
            .in0(_gnd_net_),
            .in1(N__45747),
            .in2(N__45741),
            .in3(N__50632),
            .lcout(n1632_adj_619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i970_3_lut_LC_14_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i970_3_lut_LC_14_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i970_3_lut_LC_14_20_0.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i970_3_lut_LC_14_20_0 (
            .in0(N__51391),
            .in1(_gnd_net_),
            .in2(N__50859),
            .in3(N__50879),
            .lcout(n1522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12857_1_lut_LC_14_20_1.C_ON=1'b0;
    defparam i12857_1_lut_LC_14_20_1.SEQ_MODE=4'b0000;
    defparam i12857_1_lut_LC_14_20_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12857_1_lut_LC_14_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50654),
            .lcout(n15582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_72_LC_14_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_72_LC_14_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_72_LC_14_20_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_72_LC_14_20_2 (
            .in0(N__48436),
            .in1(N__48409),
            .in2(N__50051),
            .in3(N__45840),
            .lcout(),
            .ltout(n14294_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_73_LC_14_20_3.C_ON=1'b0;
    defparam i1_4_lut_adj_73_LC_14_20_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_73_LC_14_20_3.LUT_INIT=16'b1111100011110000;
    LogicCell40 i1_4_lut_adj_73_LC_14_20_3 (
            .in0(N__50575),
            .in1(N__50746),
            .in2(N__45714),
            .in3(N__45711),
            .lcout(n14296),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i975_3_lut_LC_14_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i975_3_lut_LC_14_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i975_3_lut_LC_14_20_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i975_3_lut_LC_14_20_4 (
            .in0(_gnd_net_),
            .in1(N__51016),
            .in2(N__51401),
            .in3(N__50994),
            .lcout(n1527),
            .ltout(n1527_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_71_LC_14_20_5.C_ON=1'b0;
    defparam i1_2_lut_adj_71_LC_14_20_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_71_LC_14_20_5.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_71_LC_14_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45843),
            .in3(N__49977),
            .lcout(n14288),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i909_3_lut_LC_14_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i909_3_lut_LC_14_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i909_3_lut_LC_14_20_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i909_3_lut_LC_14_20_6 (
            .in0(_gnd_net_),
            .in1(N__48305),
            .in2(N__48285),
            .in3(N__51281),
            .lcout(n1429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_14_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_14_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_14_21_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i20_3_lut_LC_14_21_0 (
            .in0(N__45816),
            .in1(N__45834),
            .in2(_gnd_net_),
            .in3(N__46191),
            .lcout(n300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i842_3_lut_LC_14_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i842_3_lut_LC_14_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i842_3_lut_LC_14_21_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i842_3_lut_LC_14_21_1 (
            .in0(_gnd_net_),
            .in1(N__48591),
            .in2(N__51601),
            .in3(N__51638),
            .lcout(n1330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i908_3_lut_LC_14_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i908_3_lut_LC_14_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i908_3_lut_LC_14_21_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i908_3_lut_LC_14_21_3 (
            .in0(N__48725),
            .in1(_gnd_net_),
            .in2(N__51287),
            .in3(N__48273),
            .lcout(n1428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i910_3_lut_LC_14_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i910_3_lut_LC_14_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i910_3_lut_LC_14_21_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i910_3_lut_LC_14_21_4 (
            .in0(_gnd_net_),
            .in1(N__48315),
            .in2(N__48341),
            .in3(N__51266),
            .lcout(n1430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i836_3_lut_LC_14_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i836_3_lut_LC_14_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i836_3_lut_LC_14_21_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i836_3_lut_LC_14_21_5 (
            .in0(N__48855),
            .in1(_gnd_net_),
            .in2(N__51602),
            .in3(N__52200),
            .lcout(n1324),
            .ltout(n1324_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i903_3_lut_LC_14_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i903_3_lut_LC_14_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i903_3_lut_LC_14_21_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i903_3_lut_LC_14_21_6 (
            .in0(_gnd_net_),
            .in1(N__48522),
            .in2(N__45819),
            .in3(N__51270),
            .lcout(n1423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_14_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_14_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_14_21_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_14_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45815),
            .lcout(n14_adj_635),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i707_3_lut_LC_14_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i707_3_lut_LC_14_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i707_3_lut_LC_14_22_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i707_3_lut_LC_14_22_0 (
            .in0(_gnd_net_),
            .in1(N__45914),
            .in2(N__45900),
            .in3(N__46410),
            .lcout(n1131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9941_3_lut_LC_14_22_1.C_ON=1'b0;
    defparam i9941_3_lut_LC_14_22_1.SEQ_MODE=4'b0000;
    defparam i9941_3_lut_LC_14_22_1.LUT_INIT=16'b1111000010100000;
    LogicCell40 i9941_3_lut_LC_14_22_1 (
            .in0(N__48391),
            .in1(_gnd_net_),
            .in2(N__48482),
            .in3(N__48703),
            .lcout(),
            .ltout(n11908_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_176_LC_14_22_2.C_ON=1'b0;
    defparam i1_4_lut_adj_176_LC_14_22_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_176_LC_14_22_2.LUT_INIT=16'b1010100000000000;
    LogicCell40 i1_4_lut_adj_176_LC_14_22_2 (
            .in0(N__48304),
            .in1(N__48334),
            .in2(N__45891),
            .in3(N__48721),
            .lcout(),
            .ltout(n13708_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12822_4_lut_LC_14_22_3.C_ON=1'b0;
    defparam i12822_4_lut_LC_14_22_3.SEQ_MODE=4'b0000;
    defparam i12822_4_lut_LC_14_22_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12822_4_lut_LC_14_22_3 (
            .in0(N__48533),
            .in1(N__48839),
            .in2(N__45888),
            .in3(N__51075),
            .lcout(n1356),
            .ltout(n1356_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i912_3_lut_LC_14_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i912_3_lut_LC_14_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i912_3_lut_LC_14_22_4.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i912_3_lut_LC_14_22_4 (
            .in0(N__48704),
            .in1(N__48363),
            .in2(N__45885),
            .in3(_gnd_net_),
            .lcout(n1432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12819_1_lut_LC_14_22_5.C_ON=1'b0;
    defparam i12819_1_lut_LC_14_22_5.SEQ_MODE=4'b0000;
    defparam i12819_1_lut_LC_14_22_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12819_1_lut_LC_14_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51277),
            .in3(_gnd_net_),
            .lcout(n15544),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i913_3_lut_LC_14_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i913_3_lut_LC_14_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i913_3_lut_LC_14_22_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i913_3_lut_LC_14_22_6 (
            .in0(_gnd_net_),
            .in1(N__48392),
            .in2(N__48375),
            .in3(N__51248),
            .lcout(n1433),
            .ltout(n1433_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9939_3_lut_LC_14_22_7.C_ON=1'b0;
    defparam i9939_3_lut_LC_14_22_7.SEQ_MODE=4'b0000;
    defparam i9939_3_lut_LC_14_22_7.LUT_INIT=16'b1111101000000000;
    LogicCell40 i9939_3_lut_LC_14_22_7 (
            .in0(N__50521),
            .in1(_gnd_net_),
            .in2(N__45882),
            .in3(N__50443),
            .lcout(n11906),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i706_3_lut_LC_14_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i706_3_lut_LC_14_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i706_3_lut_LC_14_23_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i706_3_lut_LC_14_23_0 (
            .in0(_gnd_net_),
            .in1(N__45879),
            .in2(N__46420),
            .in3(N__45849),
            .lcout(n1130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i709_3_lut_LC_14_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i709_3_lut_LC_14_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i709_3_lut_LC_14_23_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i709_3_lut_LC_14_23_1 (
            .in0(_gnd_net_),
            .in1(N__46265),
            .in2(N__46239),
            .in3(N__46404),
            .lcout(n1133),
            .ltout(n1133_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10032_4_lut_LC_14_23_2.C_ON=1'b0;
    defparam i10032_4_lut_LC_14_23_2.SEQ_MODE=4'b0000;
    defparam i10032_4_lut_LC_14_23_2.LUT_INIT=16'b1111111010101010;
    LogicCell40 i10032_4_lut_LC_14_23_2 (
            .in0(N__51913),
            .in1(N__51463),
            .in2(N__46227),
            .in3(N__51953),
            .lcout(),
            .ltout(n12000_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12791_4_lut_LC_14_23_3.C_ON=1'b0;
    defparam i12791_4_lut_LC_14_23_3.SEQ_MODE=4'b0000;
    defparam i12791_4_lut_LC_14_23_3.LUT_INIT=16'b0000000100010001;
    LogicCell40 i12791_4_lut_LC_14_23_3 (
            .in0(N__52337),
            .in1(N__46224),
            .in2(N__46218),
            .in3(N__46341),
            .lcout(n1158),
            .ltout(n1158_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i777_3_lut_LC_14_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i777_3_lut_LC_14_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i777_3_lut_LC_14_23_4.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i777_3_lut_LC_14_23_4 (
            .in0(N__51441),
            .in1(N__51464),
            .in2(N__46215),
            .in3(_gnd_net_),
            .lcout(n1233),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i776_3_lut_LC_14_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i776_3_lut_LC_14_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i776_3_lut_LC_14_23_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i776_3_lut_LC_14_23_5 (
            .in0(_gnd_net_),
            .in1(N__51969),
            .in2(N__51429),
            .in3(N__52239),
            .lcout(n1232),
            .ltout(n1232_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9943_3_lut_LC_14_23_6.C_ON=1'b0;
    defparam i9943_3_lut_LC_14_23_6.SEQ_MODE=4'b0000;
    defparam i9943_3_lut_LC_14_23_6.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9943_3_lut_LC_14_23_6 (
            .in0(_gnd_net_),
            .in1(N__48685),
            .in2(N__46212),
            .in3(N__48655),
            .lcout(n11910),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_14_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_14_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_14_23_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i22_3_lut_LC_14_23_7 (
            .in0(N__46209),
            .in1(N__46194),
            .in2(_gnd_net_),
            .in3(N__46335),
            .lcout(n298),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i708_3_lut_LC_14_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i708_3_lut_LC_14_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i708_3_lut_LC_14_24_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i708_3_lut_LC_14_24_0 (
            .in0(_gnd_net_),
            .in1(N__45954),
            .in2(N__45948),
            .in3(N__46418),
            .lcout(n1132),
            .ltout(n1132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i775_3_lut_LC_14_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i775_3_lut_LC_14_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i775_3_lut_LC_14_24_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i775_3_lut_LC_14_24_1 (
            .in0(_gnd_net_),
            .in1(N__52240),
            .in2(N__45918),
            .in3(N__51939),
            .lcout(n1231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12774_1_lut_LC_14_24_3.C_ON=1'b0;
    defparam i12774_1_lut_LC_14_24_3.SEQ_MODE=4'b0000;
    defparam i12774_1_lut_LC_14_24_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 i12774_1_lut_LC_14_24_3 (
            .in0(N__46419),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n15499),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_53_LC_14_24_4.C_ON=1'b0;
    defparam i10_4_lut_adj_53_LC_14_24_4.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_53_LC_14_24_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_53_LC_14_24_4 (
            .in0(N__49249),
            .in1(N__54764),
            .in2(N__49589),
            .in3(N__49484),
            .lcout(n24_adj_561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_172_LC_14_24_6.C_ON=1'b0;
    defparam i1_2_lut_adj_172_LC_14_24_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_172_LC_14_24_6.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_172_LC_14_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51874),
            .in3(N__51824),
            .lcout(n14470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_14_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_14_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_14_24_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_14_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46327),
            .lcout(n12_adj_633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_14_25_0.C_ON=1'b0;
    defparam i2_2_lut_LC_14_25_0.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_14_25_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i2_2_lut_LC_14_25_0 (
            .in0(N__49537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49470),
            .lcout(),
            .ltout(n16_adj_701_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_LC_14_25_1.C_ON=1'b0;
    defparam i11_4_lut_LC_14_25_1.SEQ_MODE=4'b0000;
    defparam i11_4_lut_LC_14_25_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i11_4_lut_LC_14_25_1 (
            .in0(N__49585),
            .in1(N__49289),
            .in2(N__46290),
            .in3(N__46872),
            .lcout(n25_adj_698),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_14_26_0.C_ON=1'b0;
    defparam i4_4_lut_LC_14_26_0.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_14_26_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i4_4_lut_LC_14_26_0 (
            .in0(N__48888),
            .in1(N__49008),
            .in2(N__49056),
            .in3(N__48972),
            .lcout(n10_adj_567),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i828_4_lut_LC_14_26_2.C_ON=1'b0;
    defparam i828_4_lut_LC_14_26_2.SEQ_MODE=4'b0000;
    defparam i828_4_lut_LC_14_26_2.LUT_INIT=16'b1111000011110001;
    LogicCell40 i828_4_lut_LC_14_26_2 (
            .in0(N__46857),
            .in1(N__46287),
            .in2(N__54765),
            .in3(N__46278),
            .lcout(direction_N_340),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_14_26_4.C_ON=1'b0;
    defparam i3_4_lut_LC_14_26_4.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_14_26_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i3_4_lut_LC_14_26_4 (
            .in0(N__49156),
            .in1(N__48811),
            .in2(N__48784),
            .in3(N__48745),
            .lcout(),
            .ltout(n13932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_14_26_5.C_ON=1'b0;
    defparam i2_3_lut_LC_14_26_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_14_26_5.LUT_INIT=16'b1100000000000000;
    LogicCell40 i2_3_lut_LC_14_26_5 (
            .in0(_gnd_net_),
            .in1(N__49090),
            .in2(N__46269),
            .in3(N__49126),
            .lcout(),
            .ltout(n14110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_49_LC_14_26_6.C_ON=1'b0;
    defparam i1_4_lut_adj_49_LC_14_26_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_49_LC_14_26_6.LUT_INIT=16'b1010101010101000;
    LogicCell40 i1_4_lut_adj_49_LC_14_26_6 (
            .in0(N__49242),
            .in1(N__48927),
            .in2(N__46881),
            .in3(N__46878),
            .lcout(n15_adj_702),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9888_2_lut_LC_14_26_7.C_ON=1'b0;
    defparam i9888_2_lut_LC_14_26_7.SEQ_MODE=4'b0000;
    defparam i9888_2_lut_LC_14_26_7.LUT_INIT=16'b1111111111001100;
    LogicCell40 i9888_2_lut_LC_14_26_7 (
            .in0(_gnd_net_),
            .in1(N__49089),
            .in2(_gnd_net_),
            .in3(N__49125),
            .lcout(n11853),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_adj_54_LC_14_27_0.C_ON=1'b0;
    defparam i9_4_lut_adj_54_LC_14_27_0.SEQ_MODE=4'b0000;
    defparam i9_4_lut_adj_54_LC_14_27_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_adj_54_LC_14_27_0 (
            .in0(N__49194),
            .in1(N__49281),
            .in2(N__49333),
            .in3(N__54873),
            .lcout(n23_adj_562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12425_3_lut_4_lut_LC_14_27_4.C_ON=1'b0;
    defparam i12425_3_lut_4_lut_LC_14_27_4.SEQ_MODE=4'b0000;
    defparam i12425_3_lut_4_lut_LC_14_27_4.LUT_INIT=16'b0111101111011110;
    LogicCell40 i12425_3_lut_4_lut_LC_14_27_4 (
            .in0(N__46848),
            .in1(N__46827),
            .in2(N__46812),
            .in3(N__46789),
            .lcout(n15150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i2_3_lut_LC_14_27_5 .C_ON=1'b0;
    defparam \PWM.i2_3_lut_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \PWM.i2_3_lut_LC_14_27_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \PWM.i2_3_lut_LC_14_27_5  (
            .in0(N__46771),
            .in1(N__46740),
            .in2(_gnd_net_),
            .in3(N__46707),
            .lcout(\PWM.n13995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i11_4_lut_LC_14_27_6 .C_ON=1'b0;
    defparam \PWM.i11_4_lut_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \PWM.i11_4_lut_LC_14_27_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i11_4_lut_LC_14_27_6  (
            .in0(N__46678),
            .in1(N__46657),
            .in2(N__46638),
            .in3(N__46612),
            .lcout(\PWM.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i12_4_lut_LC_14_28_1 .C_ON=1'b0;
    defparam \PWM.i12_4_lut_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \PWM.i12_4_lut_LC_14_28_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i12_4_lut_LC_14_28_1  (
            .in0(N__46589),
            .in1(N__46559),
            .in2(N__46542),
            .in3(N__46513),
            .lcout(\PWM.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i10_4_lut_LC_14_28_2 .C_ON=1'b0;
    defparam \PWM.i10_4_lut_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \PWM.i10_4_lut_LC_14_28_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i10_4_lut_LC_14_28_2  (
            .in0(N__46495),
            .in1(N__46474),
            .in2(N__46455),
            .in3(N__47178),
            .lcout(),
            .ltout(\PWM.n26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i13_4_lut_LC_14_28_3 .C_ON=1'b0;
    defparam \PWM.i13_4_lut_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \PWM.i13_4_lut_LC_14_28_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i13_4_lut_LC_14_28_3  (
            .in0(N__47156),
            .in1(N__47058),
            .in2(N__47136),
            .in3(N__46962),
            .lcout(),
            .ltout(\PWM.n29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i9624_4_lut_LC_14_28_4 .C_ON=1'b0;
    defparam \PWM.i9624_4_lut_LC_14_28_4 .SEQ_MODE=4'b0000;
    defparam \PWM.i9624_4_lut_LC_14_28_4 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \PWM.i9624_4_lut_LC_14_28_4  (
            .in0(N__46952),
            .in1(N__47133),
            .in2(N__47127),
            .in3(N__47124),
            .lcout(\PWM.pwm_counter_31__N_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i1_4_lut_LC_14_28_6 .C_ON=1'b0;
    defparam \PWM.i1_4_lut_LC_14_28_6 .SEQ_MODE=4'b0000;
    defparam \PWM.i1_4_lut_LC_14_28_6 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \PWM.i1_4_lut_LC_14_28_6  (
            .in0(N__47086),
            .in1(N__47337),
            .in2(N__47067),
            .in3(N__47268),
            .lcout(\PWM.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_14_29_1.C_ON=1'b0;
    defparam i5_4_lut_LC_14_29_1.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_14_29_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_LC_14_29_1 (
            .in0(N__47051),
            .in1(N__47039),
            .in2(N__47028),
            .in3(N__47012),
            .lcout(),
            .ltout(n12_adj_566_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_14_29_2.C_ON=1'b0;
    defparam i6_4_lut_LC_14_29_2.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_14_29_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_14_29_2 (
            .in0(N__47000),
            .in1(N__46988),
            .in2(N__46977),
            .in3(N__46973),
            .lcout(n5162),
            .ltout(n5162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_14_29_3.C_ON=1'b0;
    defparam i1_2_lut_LC_14_29_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_14_29_3.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_LC_14_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46956),
            .in3(N__46951),
            .lcout(n5164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i8_LC_14_29_4.C_ON=1'b0;
    defparam pwm_setpoint_i8_LC_14_29_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i8_LC_14_29_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i8_LC_14_29_4 (
            .in0(N__55322),
            .in1(N__46923),
            .in2(_gnd_net_),
            .in3(N__46907),
            .lcout(pwm_setpoint_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55820),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i9_2_lut_LC_14_29_5.C_ON=1'b0;
    defparam LessThan_299_i9_2_lut_LC_14_29_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i9_2_lut_LC_14_29_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i9_2_lut_LC_14_29_5 (
            .in0(_gnd_net_),
            .in1(N__47490),
            .in2(_gnd_net_),
            .in3(N__47469),
            .lcout(n9_adj_658),
            .ltout(n9_adj_658_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12480_4_lut_LC_14_29_6.C_ON=1'b0;
    defparam i12480_4_lut_LC_14_29_6.SEQ_MODE=4'b0000;
    defparam i12480_4_lut_LC_14_29_6.LUT_INIT=16'b1111111111001101;
    LogicCell40 i12480_4_lut_LC_14_29_6 (
            .in0(N__47454),
            .in1(N__47435),
            .in2(N__47424),
            .in3(N__47417),
            .lcout(n15205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12476_4_lut_LC_14_30_0.C_ON=1'b0;
    defparam i12476_4_lut_LC_14_30_0.SEQ_MODE=4'b0000;
    defparam i12476_4_lut_LC_14_30_0.LUT_INIT=16'b1110111011101111;
    LogicCell40 i12476_4_lut_LC_14_30_0 (
            .in0(N__47210),
            .in1(N__47228),
            .in2(N__47403),
            .in3(N__47388),
            .lcout(),
            .ltout(n15201_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12536_4_lut_LC_14_30_1.C_ON=1'b0;
    defparam i12536_4_lut_LC_14_30_1.SEQ_MODE=4'b0000;
    defparam i12536_4_lut_LC_14_30_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12536_4_lut_LC_14_30_1 (
            .in0(N__47743),
            .in1(N__47722),
            .in2(N__47382),
            .in3(N__47246),
            .lcout(n15261),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i17_2_lut_LC_14_30_4.C_ON=1'b0;
    defparam LessThan_299_i17_2_lut_LC_14_30_4.SEQ_MODE=4'b0000;
    defparam LessThan_299_i17_2_lut_LC_14_30_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i17_2_lut_LC_14_30_4 (
            .in0(_gnd_net_),
            .in1(N__47357),
            .in2(_gnd_net_),
            .in3(N__47345),
            .lcout(n17_adj_665),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i19_2_lut_LC_14_30_5.C_ON=1'b0;
    defparam LessThan_299_i19_2_lut_LC_14_30_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i19_2_lut_LC_14_30_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i19_2_lut_LC_14_30_5 (
            .in0(_gnd_net_),
            .in1(N__47305),
            .in2(_gnd_net_),
            .in3(N__47276),
            .lcout(n19_adj_666),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12380_2_lut_4_lut_LC_14_30_6.C_ON=1'b0;
    defparam i12380_2_lut_4_lut_LC_14_30_6.SEQ_MODE=4'b0000;
    defparam i12380_2_lut_4_lut_LC_14_30_6.LUT_INIT=16'b0000100000000010;
    LogicCell40 i12380_2_lut_4_lut_LC_14_30_6 (
            .in0(N__49764),
            .in1(N__54693),
            .in2(N__54637),
            .in3(N__56100),
            .lcout(n15088),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12416_2_lut_4_lut_LC_14_30_7.C_ON=1'b0;
    defparam i12416_2_lut_4_lut_LC_14_30_7.SEQ_MODE=4'b0000;
    defparam i12416_2_lut_4_lut_LC_14_30_7.LUT_INIT=16'b0010000100000000;
    LogicCell40 i12416_2_lut_4_lut_LC_14_30_7 (
            .in0(N__56099),
            .in1(N__54624),
            .in2(N__54699),
            .in3(N__49610),
            .lcout(n15091),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12407_4_lut_LC_14_31_0.C_ON=1'b0;
    defparam i12407_4_lut_LC_14_31_0.SEQ_MODE=4'b0000;
    defparam i12407_4_lut_LC_14_31_0.LUT_INIT=16'b1010101010101011;
    LogicCell40 i12407_4_lut_LC_14_31_0 (
            .in0(N__47247),
            .in1(N__47229),
            .in2(N__47217),
            .in3(N__47199),
            .lcout(),
            .ltout(n15132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12385_4_lut_LC_14_31_1.C_ON=1'b0;
    defparam i12385_4_lut_LC_14_31_1.SEQ_MODE=4'b0000;
    defparam i12385_4_lut_LC_14_31_1.LUT_INIT=16'b1010101010101011;
    LogicCell40 i12385_4_lut_LC_14_31_1 (
            .in0(N__47756),
            .in1(N__47745),
            .in2(N__47727),
            .in3(N__47724),
            .lcout(n15110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12420_2_lut_4_lut_LC_14_31_2.C_ON=1'b0;
    defparam i12420_2_lut_4_lut_LC_14_31_2.SEQ_MODE=4'b0000;
    defparam i12420_2_lut_4_lut_LC_14_31_2.LUT_INIT=16'b0000100100000000;
    LogicCell40 i12420_2_lut_4_lut_LC_14_31_2 (
            .in0(N__54684),
            .in1(N__56101),
            .in2(N__54636),
            .in3(N__49735),
            .lcout(n15095),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i1_LC_14_31_4.C_ON=1'b0;
    defparam commutation_state_i1_LC_14_31_4.SEQ_MODE=4'b1000;
    defparam commutation_state_i1_LC_14_31_4.LUT_INIT=16'b1011001100010000;
    LogicCell40 commutation_state_i1_LC_14_31_4 (
            .in0(N__47635),
            .in1(N__47689),
            .in2(N__56029),
            .in3(N__47586),
            .lcout(commutation_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55826),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_14_31_5.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_14_31_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_14_31_5.LUT_INIT=16'b0000000001000100;
    LogicCell40 i2_2_lut_3_lut_LC_14_31_5 (
            .in0(N__47585),
            .in1(N__47685),
            .in2(_gnd_net_),
            .in3(N__47634),
            .lcout(commutation_state_7__N_261),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12419_2_lut_4_lut_LC_14_32_1.C_ON=1'b0;
    defparam i12419_2_lut_4_lut_LC_14_32_1.SEQ_MODE=4'b0000;
    defparam i12419_2_lut_4_lut_LC_14_32_1.LUT_INIT=16'b0010000000010000;
    LogicCell40 i12419_2_lut_4_lut_LC_14_32_1 (
            .in0(N__56118),
            .in1(N__54623),
            .in2(N__49703),
            .in3(N__54671),
            .lcout(n15094),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i2_LC_14_32_6.C_ON=1'b0;
    defparam commutation_state_i2_LC_14_32_6.SEQ_MODE=4'b1000;
    defparam commutation_state_i2_LC_14_32_6.LUT_INIT=16'b1010001000110010;
    LogicCell40 commutation_state_i2_LC_14_32_6 (
            .in0(N__47691),
            .in1(N__47636),
            .in2(N__55950),
            .in3(N__47596),
            .lcout(commutation_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55829),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_15_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_15_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_15_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_2_lut_LC_15_17_0 (
            .in0(_gnd_net_),
            .in1(N__47543),
            .in2(_gnd_net_),
            .in3(N__47502),
            .lcout(n1701),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(n12563),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_15_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_15_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_15_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_3_lut_LC_15_17_1 (
            .in0(_gnd_net_),
            .in1(N__54188),
            .in2(N__48192),
            .in3(N__47493),
            .lcout(n1700),
            .ltout(),
            .carryin(n12563),
            .carryout(n12564),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_15_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_15_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_15_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_4_lut_LC_15_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47895),
            .in3(N__47865),
            .lcout(n1699),
            .ltout(),
            .carryin(n12564),
            .carryout(n12565),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_15_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_15_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_15_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_5_lut_LC_15_17_3 (
            .in0(_gnd_net_),
            .in1(N__54189),
            .in2(N__47862),
            .in3(N__47835),
            .lcout(n1698),
            .ltout(),
            .carryin(n12565),
            .carryout(n12566),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_15_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_15_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_15_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_6_lut_LC_15_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47832),
            .in3(N__47811),
            .lcout(n1697),
            .ltout(),
            .carryin(n12566),
            .carryout(n12567),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_15_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_15_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_15_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_7_lut_LC_15_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50555),
            .in3(N__47808),
            .lcout(n1696),
            .ltout(),
            .carryin(n12567),
            .carryout(n12568),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_15_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_15_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_15_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_8_lut_LC_15_17_6 (
            .in0(_gnd_net_),
            .in1(N__54190),
            .in2(N__50711),
            .in3(N__47805),
            .lcout(n1695),
            .ltout(),
            .carryin(n12568),
            .carryout(n12569),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_15_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_15_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_15_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_9_lut_LC_15_17_7 (
            .in0(_gnd_net_),
            .in1(N__49928),
            .in2(N__54359),
            .in3(N__47796),
            .lcout(n1694),
            .ltout(),
            .carryin(n12569),
            .carryout(n12570),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_15_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_15_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_15_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_10_lut_LC_15_18_0 (
            .in0(_gnd_net_),
            .in1(N__53090),
            .in2(N__50769),
            .in3(N__47793),
            .lcout(n1693_adj_621),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(n12571),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_15_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_15_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_11_lut_LC_15_18_1 (
            .in0(_gnd_net_),
            .in1(N__53095),
            .in2(N__50012),
            .in3(N__47790),
            .lcout(n1692),
            .ltout(),
            .carryin(n12571),
            .carryout(n12572),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_15_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_15_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_15_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_12_lut_LC_15_18_2 (
            .in0(_gnd_net_),
            .in1(N__47785),
            .in2(N__53451),
            .in3(N__47760),
            .lcout(n1691),
            .ltout(),
            .carryin(n12572),
            .carryout(n12573),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_15_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_15_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_15_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_13_lut_LC_15_18_3 (
            .in0(_gnd_net_),
            .in1(N__53099),
            .in2(N__48126),
            .in3(N__48075),
            .lcout(n1690),
            .ltout(),
            .carryin(n12573),
            .carryout(n12574),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_15_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_15_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_15_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_14_lut_LC_15_18_4 (
            .in0(_gnd_net_),
            .in1(N__53091),
            .in2(N__48071),
            .in3(N__48030),
            .lcout(n1689),
            .ltout(),
            .carryin(n12574),
            .carryout(n12575),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_15_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_15_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_15_lut_LC_15_18_5 (
            .in0(_gnd_net_),
            .in1(N__48022),
            .in2(N__53450),
            .in3(N__47991),
            .lcout(n1688),
            .ltout(),
            .carryin(n12575),
            .carryout(n12576),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_15_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_15_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_15_18_6.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1101_16_lut_LC_15_18_6 (
            .in0(N__53100),
            .in1(N__47981),
            .in2(N__47970),
            .in3(N__47946),
            .lcout(n1719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_15_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_15_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_15_18_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1108_3_lut_LC_15_18_7 (
            .in0(_gnd_net_),
            .in1(N__47922),
            .in2(N__50013),
            .in3(N__50165),
            .lcout(n1724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i978_3_lut_LC_15_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i978_3_lut_LC_15_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i978_3_lut_LC_15_19_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i978_3_lut_LC_15_19_0 (
            .in0(_gnd_net_),
            .in1(N__50414),
            .in2(N__51398),
            .in3(N__50394),
            .lcout(n1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i911_3_lut_LC_15_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i911_3_lut_LC_15_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i911_3_lut_LC_15_19_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i911_3_lut_LC_15_19_1 (
            .in0(_gnd_net_),
            .in1(N__48354),
            .in2(N__48486),
            .in3(N__51282),
            .lcout(n1431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i971_3_lut_LC_15_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i971_3_lut_LC_15_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i971_3_lut_LC_15_19_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i971_3_lut_LC_15_19_2 (
            .in0(_gnd_net_),
            .in1(N__51212),
            .in2(N__51399),
            .in3(N__50895),
            .lcout(n1523),
            .ltout(n1523_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12860_4_lut_LC_15_19_3.C_ON=1'b0;
    defparam i12860_4_lut_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam i12860_4_lut_LC_15_19_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12860_4_lut_LC_15_19_3 (
            .in0(N__50813),
            .in1(N__48262),
            .in2(N__48246),
            .in3(N__48243),
            .lcout(n1554),
            .ltout(n1554_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_15_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_15_19_4.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1049_3_lut_LC_15_19_4 (
            .in0(N__48237),
            .in1(_gnd_net_),
            .in2(N__48228),
            .in3(N__48225),
            .lcout(n1633_adj_620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i977_3_lut_LC_15_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i977_3_lut_LC_15_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i977_3_lut_LC_15_19_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i977_3_lut_LC_15_19_5 (
            .in0(_gnd_net_),
            .in1(N__50355),
            .in2(N__50385),
            .in3(N__51379),
            .lcout(n1529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i980_3_lut_LC_15_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i980_3_lut_LC_15_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i980_3_lut_LC_15_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i980_3_lut_LC_15_19_7 (
            .in0(_gnd_net_),
            .in1(N__50466),
            .in2(N__50490),
            .in3(N__51375),
            .lcout(n1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_178_LC_15_20_0.C_ON=1'b0;
    defparam i1_4_lut_adj_178_LC_15_20_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_178_LC_15_20_0.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_178_LC_15_20_0 (
            .in0(N__50410),
            .in1(N__51055),
            .in2(N__48141),
            .in3(N__50371),
            .lcout(n13727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i906_3_lut_LC_15_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i906_3_lut_LC_15_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i906_3_lut_LC_15_20_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i906_3_lut_LC_15_20_1 (
            .in0(_gnd_net_),
            .in1(N__51120),
            .in2(N__51295),
            .in3(N__48561),
            .lcout(n1426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i905_3_lut_LC_15_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i905_3_lut_LC_15_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i905_3_lut_LC_15_20_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i905_3_lut_LC_15_20_2 (
            .in0(N__48552),
            .in1(_gnd_net_),
            .in2(N__51099),
            .in3(N__51283),
            .lcout(n1425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_177_LC_15_20_3.C_ON=1'b0;
    defparam i1_2_lut_adj_177_LC_15_20_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_177_LC_15_20_3.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_177_LC_15_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51020),
            .in3(N__50978),
            .lcout(),
            .ltout(n14490_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_179_LC_15_20_4.C_ON=1'b0;
    defparam i1_4_lut_adj_179_LC_15_20_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_179_LC_15_20_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_179_LC_15_20_4 (
            .in0(N__50920),
            .in1(N__50947),
            .in2(N__48129),
            .in3(N__51211),
            .lcout(),
            .ltout(n14496_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12841_4_lut_LC_15_20_5.C_ON=1'b0;
    defparam i12841_4_lut_LC_15_20_5.SEQ_MODE=4'b0000;
    defparam i12841_4_lut_LC_15_20_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12841_4_lut_LC_15_20_5 (
            .in0(N__50875),
            .in1(N__48456),
            .in2(N__48450),
            .in3(N__50840),
            .lcout(n1455),
            .ltout(n1455_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i973_3_lut_LC_15_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i973_3_lut_LC_15_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i973_3_lut_LC_15_20_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i973_3_lut_LC_15_20_6 (
            .in0(_gnd_net_),
            .in1(N__50948),
            .in2(N__48447),
            .in3(N__50934),
            .lcout(n1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i972_3_lut_LC_15_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i972_3_lut_LC_15_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i972_3_lut_LC_15_20_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i972_3_lut_LC_15_20_7 (
            .in0(_gnd_net_),
            .in1(N__50921),
            .in2(N__50907),
            .in3(N__51392),
            .lcout(n1524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_15_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_15_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_15_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_2_lut_LC_15_21_0 (
            .in0(_gnd_net_),
            .in1(N__48393),
            .in2(_gnd_net_),
            .in3(N__48366),
            .lcout(n1401),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(n12527),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_15_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_15_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_15_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_3_lut_LC_15_21_1 (
            .in0(_gnd_net_),
            .in1(N__53196),
            .in2(N__48705),
            .in3(N__48357),
            .lcout(n1400),
            .ltout(),
            .carryin(n12527),
            .carryout(n12528),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_15_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_15_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_15_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_4_lut_LC_15_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48481),
            .in3(N__48345),
            .lcout(n1399),
            .ltout(),
            .carryin(n12528),
            .carryout(n12529),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_15_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_15_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_15_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_5_lut_LC_15_21_3 (
            .in0(_gnd_net_),
            .in1(N__53197),
            .in2(N__48342),
            .in3(N__48309),
            .lcout(n1398),
            .ltout(),
            .carryin(n12529),
            .carryout(n12530),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_15_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_15_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_6_lut_LC_15_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48306),
            .in3(N__48276),
            .lcout(n1397),
            .ltout(),
            .carryin(n12530),
            .carryout(n12531),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_15_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_15_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_15_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_7_lut_LC_15_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48726),
            .in3(N__48267),
            .lcout(n1396),
            .ltout(),
            .carryin(n12531),
            .carryout(n12532),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_15_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_15_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_15_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_8_lut_LC_15_21_6 (
            .in0(_gnd_net_),
            .in1(N__53198),
            .in2(N__51137),
            .in3(N__48564),
            .lcout(n1395),
            .ltout(),
            .carryin(n12532),
            .carryout(n12533),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_15_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_15_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_15_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_9_lut_LC_15_21_7 (
            .in0(_gnd_net_),
            .in1(N__51119),
            .in2(N__53576),
            .in3(N__48555),
            .lcout(n1394),
            .ltout(),
            .carryin(n12533),
            .carryout(n12534),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_15_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_15_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_15_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_10_lut_LC_15_22_0 (
            .in0(_gnd_net_),
            .in1(N__52898),
            .in2(N__51098),
            .in3(N__48543),
            .lcout(n1393),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(n12535),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_15_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_15_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_15_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_11_lut_LC_15_22_1 (
            .in0(_gnd_net_),
            .in1(N__52979),
            .in2(N__51687),
            .in3(N__48540),
            .lcout(n1392),
            .ltout(),
            .carryin(n12535),
            .carryout(n12536),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_15_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_15_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_15_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_12_lut_LC_15_22_2 (
            .in0(_gnd_net_),
            .in1(N__52899),
            .in2(N__48537),
            .in3(N__48516),
            .lcout(n1391),
            .ltout(),
            .carryin(n12536),
            .carryout(n12537),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_15_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_15_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_15_22_3.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_900_13_lut_LC_15_22_3 (
            .in0(N__52900),
            .in1(N__48840),
            .in2(N__48506),
            .in3(N__48489),
            .lcout(n1422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i771_3_lut_LC_15_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i771_3_lut_LC_15_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i771_3_lut_LC_15_22_4.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i771_3_lut_LC_15_22_4 (
            .in0(_gnd_net_),
            .in1(N__52245),
            .in2(N__51803),
            .in3(N__51771),
            .lcout(n1227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i844_3_lut_LC_15_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i844_3_lut_LC_15_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i844_3_lut_LC_15_22_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i844_3_lut_LC_15_22_5 (
            .in0(N__48659),
            .in1(_gnd_net_),
            .in2(N__48639),
            .in3(N__51582),
            .lcout(n1332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i841_3_lut_LC_15_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i841_3_lut_LC_15_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i841_3_lut_LC_15_22_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i841_3_lut_LC_15_22_6 (
            .in0(_gnd_net_),
            .in1(N__48579),
            .in2(N__51597),
            .in3(N__51488),
            .lcout(n1329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i845_3_lut_LC_15_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i845_3_lut_LC_15_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i845_3_lut_LC_15_22_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i845_3_lut_LC_15_22_7 (
            .in0(N__48669),
            .in1(N__48687),
            .in2(_gnd_net_),
            .in3(N__51581),
            .lcout(n1333),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_15_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_15_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_15_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_2_lut_LC_15_23_0 (
            .in0(_gnd_net_),
            .in1(N__48686),
            .in2(_gnd_net_),
            .in3(N__48663),
            .lcout(n1301),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(n12517),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_15_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_15_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_15_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_3_lut_LC_15_23_1 (
            .in0(_gnd_net_),
            .in1(N__52973),
            .in2(N__48660),
            .in3(N__48630),
            .lcout(n1300),
            .ltout(),
            .carryin(n12517),
            .carryout(n12518),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_15_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_15_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_15_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_4_lut_LC_15_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48623),
            .in3(N__48594),
            .lcout(n1299),
            .ltout(),
            .carryin(n12518),
            .carryout(n12519),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_15_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_15_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_15_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_5_lut_LC_15_23_3 (
            .in0(_gnd_net_),
            .in1(N__52974),
            .in2(N__51637),
            .in3(N__48582),
            .lcout(n1298),
            .ltout(),
            .carryin(n12519),
            .carryout(n12520),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_15_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_15_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_15_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_6_lut_LC_15_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51489),
            .in3(N__48573),
            .lcout(n1297),
            .ltout(),
            .carryin(n12520),
            .carryout(n12521),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_15_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_15_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_15_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_7_lut_LC_15_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51669),
            .in3(N__48570),
            .lcout(n1296),
            .ltout(),
            .carryin(n12521),
            .carryout(n12522),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_15_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_15_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_15_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_8_lut_LC_15_23_6 (
            .in0(_gnd_net_),
            .in1(N__52975),
            .in2(N__51507),
            .in3(N__48567),
            .lcout(n1295),
            .ltout(),
            .carryin(n12522),
            .carryout(n12523),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_15_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_15_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_15_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_9_lut_LC_15_23_7 (
            .in0(_gnd_net_),
            .in1(N__51166),
            .in2(N__53339),
            .in3(N__48861),
            .lcout(n1294),
            .ltout(),
            .carryin(n12523),
            .carryout(n12524),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_15_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_15_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_15_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_10_lut_LC_15_24_0 (
            .in0(_gnd_net_),
            .in1(N__52891),
            .in2(N__51720),
            .in3(N__48858),
            .lcout(n1293),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(n12525),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_15_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_15_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_15_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_11_lut_LC_15_24_1 (
            .in0(_gnd_net_),
            .in1(N__52971),
            .in2(N__52196),
            .in3(N__48846),
            .lcout(n1292),
            .ltout(),
            .carryin(n12525),
            .carryout(n12526),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_15_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_15_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_15_24_2.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_833_12_lut_LC_15_24_2 (
            .in0(N__52972),
            .in1(N__51521),
            .in2(N__52323),
            .in3(N__48843),
            .lcout(n1323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12788_1_lut_LC_15_24_4.C_ON=1'b0;
    defparam i12788_1_lut_LC_15_24_4.SEQ_MODE=4'b0000;
    defparam i12788_1_lut_LC_15_24_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12788_1_lut_LC_15_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52241),
            .lcout(n15513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_305_1_LC_15_25_0.C_ON=1'b1;
    defparam add_305_1_LC_15_25_0.SEQ_MODE=4'b0000;
    defparam add_305_1_LC_15_25_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_305_1_LC_15_25_0 (
            .in0(_gnd_net_),
            .in1(N__52035),
            .in2(N__52082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(n12435),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i0_LC_15_25_1.C_ON=1'b1;
    defparam encoder0_position_target_i0_i0_LC_15_25_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i0_LC_15_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i0_LC_15_25_1 (
            .in0(_gnd_net_),
            .in1(N__48815),
            .in2(N__52146),
            .in3(N__48795),
            .lcout(encoder0_position_target_0),
            .ltout(),
            .carryin(n12435),
            .carryout(n12436),
            .clk(N__55805),
            .ce(N__55399),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i1_LC_15_25_2.C_ON=1'b1;
    defparam encoder0_position_target_i0_i1_LC_15_25_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i1_LC_15_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i1_LC_15_25_2 (
            .in0(_gnd_net_),
            .in1(N__52036),
            .in2(N__48788),
            .in3(N__48759),
            .lcout(encoder0_position_target_1),
            .ltout(),
            .carryin(n12436),
            .carryout(n12437),
            .clk(N__55805),
            .ce(N__55399),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i2_LC_15_25_3.C_ON=1'b1;
    defparam encoder0_position_target_i0_i2_LC_15_25_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i2_LC_15_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i2_LC_15_25_3 (
            .in0(_gnd_net_),
            .in1(N__52042),
            .in2(N__48755),
            .in3(N__48729),
            .lcout(encoder0_position_target_2),
            .ltout(),
            .carryin(n12437),
            .carryout(n12438),
            .clk(N__55805),
            .ce(N__55399),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i3_LC_15_25_4.C_ON=1'b1;
    defparam encoder0_position_target_i0_i3_LC_15_25_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i3_LC_15_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i3_LC_15_25_4 (
            .in0(_gnd_net_),
            .in1(N__52037),
            .in2(N__49166),
            .in3(N__49140),
            .lcout(encoder0_position_target_3),
            .ltout(),
            .carryin(n12438),
            .carryout(n12439),
            .clk(N__55805),
            .ce(N__55399),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i4_LC_15_25_5.C_ON=1'b1;
    defparam encoder0_position_target_i0_i4_LC_15_25_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i4_LC_15_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i4_LC_15_25_5 (
            .in0(_gnd_net_),
            .in1(N__52043),
            .in2(N__49136),
            .in3(N__49107),
            .lcout(encoder0_position_target_4),
            .ltout(),
            .carryin(n12439),
            .carryout(n12440),
            .clk(N__55805),
            .ce(N__55399),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i5_LC_15_25_6.C_ON=1'b1;
    defparam encoder0_position_target_i0_i5_LC_15_25_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i5_LC_15_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i5_LC_15_25_6 (
            .in0(_gnd_net_),
            .in1(N__52038),
            .in2(N__49100),
            .in3(N__49071),
            .lcout(encoder0_position_target_5),
            .ltout(),
            .carryin(n12440),
            .carryout(n12441),
            .clk(N__55805),
            .ce(N__55399),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i6_LC_15_25_7.C_ON=1'b1;
    defparam encoder0_position_target_i0_i6_LC_15_25_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i6_LC_15_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i6_LC_15_25_7 (
            .in0(_gnd_net_),
            .in1(N__52044),
            .in2(N__49057),
            .in3(N__49023),
            .lcout(encoder0_position_target_6),
            .ltout(),
            .carryin(n12441),
            .carryout(n12442),
            .clk(N__55805),
            .ce(N__55399),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i7_LC_15_26_0.C_ON=1'b1;
    defparam encoder0_position_target_i0_i7_LC_15_26_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i7_LC_15_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i7_LC_15_26_0 (
            .in0(_gnd_net_),
            .in1(N__52045),
            .in2(N__49018),
            .in3(N__48987),
            .lcout(encoder0_position_target_7),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(n12443),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i8_LC_15_26_1.C_ON=1'b1;
    defparam encoder0_position_target_i0_i8_LC_15_26_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i8_LC_15_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i8_LC_15_26_1 (
            .in0(_gnd_net_),
            .in1(N__48976),
            .in2(N__52083),
            .in3(N__48948),
            .lcout(encoder0_position_target_8),
            .ltout(),
            .carryin(n12443),
            .carryout(n12444),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i9_LC_15_26_2.C_ON=1'b1;
    defparam encoder0_position_target_i0_i9_LC_15_26_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i9_LC_15_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i9_LC_15_26_2 (
            .in0(_gnd_net_),
            .in1(N__52049),
            .in2(N__48941),
            .in3(N__48903),
            .lcout(encoder0_position_target_9),
            .ltout(),
            .carryin(n12444),
            .carryout(n12445),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i10_LC_15_26_3.C_ON=1'b1;
    defparam encoder0_position_target_i0_i10_LC_15_26_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i10_LC_15_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i10_LC_15_26_3 (
            .in0(_gnd_net_),
            .in1(N__48889),
            .in2(N__52084),
            .in3(N__48864),
            .lcout(encoder0_position_target_10),
            .ltout(),
            .carryin(n12445),
            .carryout(n12446),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i11_LC_15_26_4.C_ON=1'b1;
    defparam encoder0_position_target_i0_i11_LC_15_26_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i11_LC_15_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i11_LC_15_26_4 (
            .in0(_gnd_net_),
            .in1(N__52053),
            .in2(N__49483),
            .in3(N__49446),
            .lcout(encoder0_position_target_11),
            .ltout(),
            .carryin(n12446),
            .carryout(n12447),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i12_LC_15_26_5.C_ON=1'b1;
    defparam encoder0_position_target_i0_i12_LC_15_26_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i12_LC_15_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i12_LC_15_26_5 (
            .in0(_gnd_net_),
            .in1(N__49425),
            .in2(N__52085),
            .in3(N__49395),
            .lcout(encoder0_position_target_12),
            .ltout(),
            .carryin(n12447),
            .carryout(n12448),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i13_LC_15_26_6.C_ON=1'b1;
    defparam encoder0_position_target_i0_i13_LC_15_26_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i13_LC_15_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i13_LC_15_26_6 (
            .in0(_gnd_net_),
            .in1(N__52057),
            .in2(N__49387),
            .in3(N__49347),
            .lcout(encoder0_position_target_13),
            .ltout(),
            .carryin(n12448),
            .carryout(n12449),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i14_LC_15_26_7.C_ON=1'b1;
    defparam encoder0_position_target_i0_i14_LC_15_26_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i14_LC_15_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i14_LC_15_26_7 (
            .in0(_gnd_net_),
            .in1(N__49332),
            .in2(N__52086),
            .in3(N__49302),
            .lcout(encoder0_position_target_14),
            .ltout(),
            .carryin(n12449),
            .carryout(n12450),
            .clk(N__55810),
            .ce(N__55389),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i15_LC_15_27_0.C_ON=1'b1;
    defparam encoder0_position_target_i0_i15_LC_15_27_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i15_LC_15_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i15_LC_15_27_0 (
            .in0(_gnd_net_),
            .in1(N__52087),
            .in2(N__54882),
            .in3(N__49299),
            .lcout(encoder0_position_target_15),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(n12451),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i16_LC_15_27_1.C_ON=1'b1;
    defparam encoder0_position_target_i0_i16_LC_15_27_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i16_LC_15_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i16_LC_15_27_1 (
            .in0(_gnd_net_),
            .in1(N__49288),
            .in2(N__52106),
            .in3(N__49260),
            .lcout(encoder0_position_target_16),
            .ltout(),
            .carryin(n12451),
            .carryout(n12452),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i17_LC_15_27_2.C_ON=1'b1;
    defparam encoder0_position_target_i0_i17_LC_15_27_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i17_LC_15_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i17_LC_15_27_2 (
            .in0(_gnd_net_),
            .in1(N__52091),
            .in2(N__49253),
            .in3(N__49218),
            .lcout(encoder0_position_target_17),
            .ltout(),
            .carryin(n12452),
            .carryout(n12453),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i18_LC_15_27_3.C_ON=1'b1;
    defparam encoder0_position_target_i0_i18_LC_15_27_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i18_LC_15_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i18_LC_15_27_3 (
            .in0(_gnd_net_),
            .in1(N__49207),
            .in2(N__52107),
            .in3(N__49176),
            .lcout(encoder0_position_target_18),
            .ltout(),
            .carryin(n12453),
            .carryout(n12454),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i19_LC_15_27_4.C_ON=1'b1;
    defparam encoder0_position_target_i0_i19_LC_15_27_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i19_LC_15_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i19_LC_15_27_4 (
            .in0(_gnd_net_),
            .in1(N__52095),
            .in2(N__54805),
            .in3(N__49173),
            .lcout(encoder0_position_target_19),
            .ltout(),
            .carryin(n12454),
            .carryout(n12455),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i20_LC_15_27_5.C_ON=1'b1;
    defparam encoder0_position_target_i0_i20_LC_15_27_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i20_LC_15_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i20_LC_15_27_5 (
            .in0(_gnd_net_),
            .in1(N__49581),
            .in2(N__52108),
            .in3(N__49554),
            .lcout(encoder0_position_target_20),
            .ltout(),
            .carryin(n12455),
            .carryout(n12456),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i21_LC_15_27_6.C_ON=1'b1;
    defparam encoder0_position_target_i0_i21_LC_15_27_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i21_LC_15_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i21_LC_15_27_6 (
            .in0(_gnd_net_),
            .in1(N__52099),
            .in2(N__54847),
            .in3(N__49551),
            .lcout(encoder0_position_target_21),
            .ltout(),
            .carryin(n12456),
            .carryout(n12457),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i22_LC_15_27_7.C_ON=1'b1;
    defparam encoder0_position_target_i0_i22_LC_15_27_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i22_LC_15_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i22_LC_15_27_7 (
            .in0(_gnd_net_),
            .in1(N__49533),
            .in2(N__52109),
            .in3(N__49506),
            .lcout(encoder0_position_target_22),
            .ltout(),
            .carryin(n12457),
            .carryout(n12458),
            .clk(N__55817),
            .ce(N__55402),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i23_LC_15_28_0.C_ON=1'b0;
    defparam encoder0_position_target_i0_i23_LC_15_28_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i23_LC_15_28_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 encoder0_position_target_i0_i23_LC_15_28_0 (
            .in0(N__52110),
            .in1(N__54755),
            .in2(_gnd_net_),
            .in3(N__49503),
            .lcout(encoder0_position_target_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55821),
            .ce(N__55404),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_60_LC_15_29_6.C_ON=1'b0;
    defparam i2_2_lut_adj_60_LC_15_29_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_60_LC_15_29_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_adj_60_LC_15_29_6 (
            .in0(_gnd_net_),
            .in1(N__49699),
            .in2(_gnd_net_),
            .in3(N__49736),
            .lcout(n10_adj_719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12417_2_lut_4_lut_LC_15_30_1.C_ON=1'b0;
    defparam i12417_2_lut_4_lut_LC_15_30_1.SEQ_MODE=4'b0000;
    defparam i12417_2_lut_4_lut_LC_15_30_1.LUT_INIT=16'b0000100000000100;
    LogicCell40 i12417_2_lut_4_lut_LC_15_30_1 (
            .in0(N__56110),
            .in1(N__49639),
            .in2(N__54638),
            .in3(N__54688),
            .lcout(n15092),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_61_LC_15_30_3.C_ON=1'b0;
    defparam i6_4_lut_adj_61_LC_15_30_3.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_61_LC_15_30_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_61_LC_15_30_3 (
            .in0(N__49609),
            .in1(N__49861),
            .in2(N__49643),
            .in3(N__49840),
            .lcout(),
            .ltout(n14_adj_718_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_15_30_4.C_ON=1'b0;
    defparam i7_4_lut_LC_15_30_4.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_15_30_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i7_4_lut_LC_15_30_4 (
            .in0(N__49666),
            .in1(N__49762),
            .in2(N__49500),
            .in3(N__49497),
            .lcout(n5119),
            .ltout(n5119_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9549_2_lut_LC_15_30_5.C_ON=1'b0;
    defparam i9549_2_lut_LC_15_30_5.SEQ_MODE=4'b0000;
    defparam i9549_2_lut_LC_15_30_5.LUT_INIT=16'b1010000010100000;
    LogicCell40 i9549_2_lut_LC_15_30_5 (
            .in0(N__55029),
            .in1(_gnd_net_),
            .in2(N__49491),
            .in3(_gnd_net_),
            .lcout(n11514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12422_2_lut_4_lut_LC_15_30_6.C_ON=1'b0;
    defparam i12422_2_lut_4_lut_LC_15_30_6.SEQ_MODE=4'b0000;
    defparam i12422_2_lut_4_lut_LC_15_30_6.LUT_INIT=16'b0000000010000010;
    LogicCell40 i12422_2_lut_4_lut_LC_15_30_6 (
            .in0(N__49862),
            .in1(N__56112),
            .in2(N__54698),
            .in3(N__54634),
            .lcout(n15089),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12418_2_lut_4_lut_LC_15_30_7.C_ON=1'b0;
    defparam i12418_2_lut_4_lut_LC_15_30_7.SEQ_MODE=4'b0000;
    defparam i12418_2_lut_4_lut_LC_15_30_7.LUT_INIT=16'b0000100000000100;
    LogicCell40 i12418_2_lut_4_lut_LC_15_30_7 (
            .in0(N__56111),
            .in1(N__49667),
            .in2(N__54639),
            .in3(N__54689),
            .lcout(n15093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i0_LC_15_31_0.C_ON=1'b1;
    defparam dti_counter_659__i0_LC_15_31_0.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i0_LC_15_31_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 dti_counter_659__i0_LC_15_31_0 (
            .in0(N__49773),
            .in1(N__49763),
            .in2(N__54576),
            .in3(N__49746),
            .lcout(dti_counter_0),
            .ltout(),
            .carryin(bfn_15_31_0_),
            .carryout(n12961),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i1_LC_15_31_1.C_ON=1'b1;
    defparam dti_counter_659__i1_LC_15_31_1.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i1_LC_15_31_1.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_659__i1_LC_15_31_1 (
            .in0(N__49743),
            .in1(N__49737),
            .in2(N__49909),
            .in3(N__49713),
            .lcout(dti_counter_1),
            .ltout(),
            .carryin(n12961),
            .carryout(n12962),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i2_LC_15_31_2.C_ON=1'b1;
    defparam dti_counter_659__i2_LC_15_31_2.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i2_LC_15_31_2.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_659__i2_LC_15_31_2 (
            .in0(N__49710),
            .in1(N__49899),
            .in2(N__49704),
            .in3(N__49677),
            .lcout(dti_counter_2),
            .ltout(),
            .carryin(n12962),
            .carryout(n12963),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i3_LC_15_31_3.C_ON=1'b1;
    defparam dti_counter_659__i3_LC_15_31_3.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i3_LC_15_31_3.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_659__i3_LC_15_31_3 (
            .in0(N__49674),
            .in1(N__49668),
            .in2(N__49910),
            .in3(N__49653),
            .lcout(dti_counter_3),
            .ltout(),
            .carryin(n12963),
            .carryout(n12964),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i4_LC_15_31_4.C_ON=1'b1;
    defparam dti_counter_659__i4_LC_15_31_4.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i4_LC_15_31_4.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_659__i4_LC_15_31_4 (
            .in0(N__49650),
            .in1(N__49903),
            .in2(N__49644),
            .in3(N__49620),
            .lcout(dti_counter_4),
            .ltout(),
            .carryin(n12964),
            .carryout(n12965),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i5_LC_15_31_5.C_ON=1'b1;
    defparam dti_counter_659__i5_LC_15_31_5.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i5_LC_15_31_5.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_659__i5_LC_15_31_5 (
            .in0(N__49617),
            .in1(N__49611),
            .in2(N__49911),
            .in3(N__49593),
            .lcout(dti_counter_5),
            .ltout(),
            .carryin(n12965),
            .carryout(n12966),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i6_LC_15_31_6.C_ON=1'b1;
    defparam dti_counter_659__i6_LC_15_31_6.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i6_LC_15_31_6.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_659__i6_LC_15_31_6 (
            .in0(N__49824),
            .in1(N__49907),
            .in2(N__49845),
            .in3(N__49914),
            .lcout(dti_counter_6),
            .ltout(),
            .carryin(n12966),
            .carryout(n12967),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_659__i7_LC_15_31_7.C_ON=1'b0;
    defparam dti_counter_659__i7_LC_15_31_7.SEQ_MODE=4'b1000;
    defparam dti_counter_659__i7_LC_15_31_7.LUT_INIT=16'b1110010001001110;
    LogicCell40 dti_counter_659__i7_LC_15_31_7 (
            .in0(N__49908),
            .in1(N__49878),
            .in2(N__49869),
            .in3(N__49872),
            .lcout(dti_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55830),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_62_LC_15_32_1.C_ON=1'b0;
    defparam i1_4_lut_adj_62_LC_15_32_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_62_LC_15_32_1.LUT_INIT=16'b0110111111110110;
    LogicCell40 i1_4_lut_adj_62_LC_15_32_1 (
            .in0(N__49812),
            .in1(N__55920),
            .in2(N__56017),
            .in3(N__49818),
            .lcout(n4_adj_716),
            .ltout(n4_adj_716_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12404_2_lut_4_lut_LC_15_32_2.C_ON=1'b0;
    defparam i12404_2_lut_4_lut_LC_15_32_2.SEQ_MODE=4'b0000;
    defparam i12404_2_lut_4_lut_LC_15_32_2.LUT_INIT=16'b0000100100000000;
    LogicCell40 i12404_2_lut_4_lut_LC_15_32_2 (
            .in0(N__54670),
            .in1(N__56124),
            .in2(N__49848),
            .in3(N__49841),
            .lcout(n15090),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i0_LC_15_32_3.C_ON=1'b0;
    defparam commutation_state_prev_i0_LC_15_32_3.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i0_LC_15_32_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 commutation_state_prev_i0_LC_15_32_3 (
            .in0(N__56125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(commutation_state_prev_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55831),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i1_LC_15_32_5.C_ON=1'b0;
    defparam commutation_state_prev_i1_LC_15_32_5.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i1_LC_15_32_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 commutation_state_prev_i1_LC_15_32_5 (
            .in0(N__56002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(commutation_state_prev_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55831),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i2_LC_15_32_6.C_ON=1'b0;
    defparam commutation_state_prev_i2_LC_15_32_6.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i2_LC_15_32_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 commutation_state_prev_i2_LC_15_32_6 (
            .in0(N__55921),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(commutation_state_prev_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55831),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_16_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_16_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_16_17_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1109_3_lut_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(N__50765),
            .in2(N__50186),
            .in3(N__49806),
            .lcout(n1725),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1111_3_lut_LC_16_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1111_3_lut_LC_16_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1111_3_lut_LC_16_17_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1111_3_lut_LC_16_17_1 (
            .in0(_gnd_net_),
            .in1(N__49800),
            .in2(N__50712),
            .in3(N__50175),
            .lcout(n1727),
            .ltout(n1727_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_77_LC_16_17_2.C_ON=1'b0;
    defparam i1_3_lut_adj_77_LC_16_17_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_77_LC_16_17_2.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_77_LC_16_17_2 (
            .in0(_gnd_net_),
            .in1(N__50092),
            .in2(N__50346),
            .in3(N__50338),
            .lcout(),
            .ltout(n14166_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_78_LC_16_17_3.C_ON=1'b0;
    defparam i1_4_lut_adj_78_LC_16_17_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_78_LC_16_17_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_78_LC_16_17_3 (
            .in0(N__50299),
            .in1(N__50267),
            .in2(N__50256),
            .in3(N__50248),
            .lcout(n14172),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_16_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_16_17_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1112_3_lut_LC_16_17_5 (
            .in0(_gnd_net_),
            .in1(N__50208),
            .in2(N__50556),
            .in3(N__50171),
            .lcout(n1728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_74_LC_16_17_7.C_ON=1'b0;
    defparam i1_4_lut_adj_74_LC_16_17_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_74_LC_16_17_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_74_LC_16_17_7 (
            .in0(N__50764),
            .in1(N__50704),
            .in2(N__49929),
            .in3(N__50005),
            .lcout(n14508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i907_3_lut_LC_16_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i907_3_lut_LC_16_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i907_3_lut_LC_16_18_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i907_3_lut_LC_16_18_0 (
            .in0(N__51138),
            .in1(_gnd_net_),
            .in2(N__50070),
            .in3(N__51294),
            .lcout(n1427),
            .ltout(n1427_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i974_3_lut_LC_16_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i974_3_lut_LC_16_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i974_3_lut_LC_16_18_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i974_3_lut_LC_16_18_1 (
            .in0(_gnd_net_),
            .in1(N__50961),
            .in2(N__50055),
            .in3(N__51397),
            .lcout(n1526),
            .ltout(n1526_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_16_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_16_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_16_18_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1041_3_lut_LC_16_18_2 (
            .in0(_gnd_net_),
            .in1(N__50648),
            .in2(N__50028),
            .in3(N__50025),
            .lcout(n1625_adj_612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1043_3_lut_LC_16_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1043_3_lut_LC_16_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1043_3_lut_LC_16_18_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1043_3_lut_LC_16_18_4 (
            .in0(_gnd_net_),
            .in1(N__49992),
            .in2(N__49956),
            .in3(N__50647),
            .lcout(n1627_adj_614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_16_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_16_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_16_18_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1042_3_lut_LC_16_18_5 (
            .in0(_gnd_net_),
            .in1(N__50802),
            .in2(N__50667),
            .in3(N__50781),
            .lcout(n1626_adj_613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_16_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_16_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_16_18_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_16_18_6 (
            .in0(_gnd_net_),
            .in1(N__50747),
            .in2(N__50727),
            .in3(N__50646),
            .lcout(n1628_adj_615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_16_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_16_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_16_18_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1045_3_lut_LC_16_18_7 (
            .in0(_gnd_net_),
            .in1(N__50688),
            .in2(N__50666),
            .in3(N__50576),
            .lcout(n1629_adj_616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_16_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_16_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_16_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_2_lut_LC_16_19_0 (
            .in0(_gnd_net_),
            .in1(N__50528),
            .in2(_gnd_net_),
            .in3(N__50493),
            .lcout(n1501),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(n12538),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_16_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_16_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_16_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_3_lut_LC_16_19_1 (
            .in0(_gnd_net_),
            .in1(N__53609),
            .in2(N__50489),
            .in3(N__50460),
            .lcout(n1500),
            .ltout(),
            .carryin(n12538),
            .carryout(n12539),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_16_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_16_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_16_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_4_lut_LC_16_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50457),
            .in3(N__50418),
            .lcout(n1499),
            .ltout(),
            .carryin(n12539),
            .carryout(n12540),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_16_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_16_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_16_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_5_lut_LC_16_19_3 (
            .in0(_gnd_net_),
            .in1(N__53610),
            .in2(N__50415),
            .in3(N__50388),
            .lcout(n1498),
            .ltout(),
            .carryin(n12540),
            .carryout(n12541),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_16_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_16_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_16_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_6_lut_LC_16_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50384),
            .in3(N__50349),
            .lcout(n1497),
            .ltout(),
            .carryin(n12541),
            .carryout(n12542),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_16_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_16_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_16_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_7_lut_LC_16_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51063),
            .in3(N__51027),
            .lcout(n1496),
            .ltout(),
            .carryin(n12542),
            .carryout(n12543),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_16_19_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_16_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_16_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_8_lut_LC_16_19_6 (
            .in0(_gnd_net_),
            .in1(N__53615),
            .in2(N__51024),
            .in3(N__50982),
            .lcout(n1495),
            .ltout(),
            .carryin(n12543),
            .carryout(n12544),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_16_19_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_16_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_16_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_9_lut_LC_16_19_7 (
            .in0(_gnd_net_),
            .in1(N__53611),
            .in2(N__50979),
            .in3(N__50955),
            .lcout(n1494),
            .ltout(),
            .carryin(n12544),
            .carryout(n12545),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_16_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_16_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_16_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_10_lut_LC_16_20_0 (
            .in0(_gnd_net_),
            .in1(N__53607),
            .in2(N__50952),
            .in3(N__50928),
            .lcout(n1493),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(n12546),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_16_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_16_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_16_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_11_lut_LC_16_20_1 (
            .in0(_gnd_net_),
            .in1(N__53612),
            .in2(N__50925),
            .in3(N__50898),
            .lcout(n1492),
            .ltout(),
            .carryin(n12546),
            .carryout(n12547),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_16_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_16_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_16_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_12_lut_LC_16_20_2 (
            .in0(_gnd_net_),
            .in1(N__53608),
            .in2(N__51213),
            .in3(N__50889),
            .lcout(n1491),
            .ltout(),
            .carryin(n12547),
            .carryout(n12548),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_16_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_16_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_16_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_13_lut_LC_16_20_3 (
            .in0(_gnd_net_),
            .in1(N__53613),
            .in2(N__50886),
            .in3(N__50847),
            .lcout(n1490),
            .ltout(),
            .carryin(n12548),
            .carryout(n12549),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_16_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_16_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_16_20_4.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_967_14_lut_LC_16_20_4 (
            .in0(N__53614),
            .in1(N__51317),
            .in2(N__50844),
            .in3(N__50823),
            .lcout(n1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12837_1_lut_LC_16_20_5.C_ON=1'b0;
    defparam i12837_1_lut_LC_16_20_5.SEQ_MODE=4'b0000;
    defparam i12837_1_lut_LC_16_20_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12837_1_lut_LC_16_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51393),
            .lcout(n15562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i904_3_lut_LC_16_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i904_3_lut_LC_16_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i904_3_lut_LC_16_21_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i904_3_lut_LC_16_21_0 (
            .in0(N__51306),
            .in1(N__51683),
            .in2(_gnd_net_),
            .in3(N__51296),
            .lcout(n1424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i838_3_lut_LC_16_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i838_3_lut_LC_16_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i838_3_lut_LC_16_21_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i838_3_lut_LC_16_21_1 (
            .in0(_gnd_net_),
            .in1(N__51168),
            .in2(N__51589),
            .in3(N__51189),
            .lcout(n1326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i839_3_lut_LC_16_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i839_3_lut_LC_16_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i839_3_lut_LC_16_21_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i839_3_lut_LC_16_21_2 (
            .in0(N__51506),
            .in1(_gnd_net_),
            .in2(N__51180),
            .in3(N__51569),
            .lcout(n1327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_173_LC_16_21_3.C_ON=1'b0;
    defparam i1_3_lut_adj_173_LC_16_21_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_173_LC_16_21_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_173_LC_16_21_3 (
            .in0(_gnd_net_),
            .in1(N__51167),
            .in2(N__51719),
            .in3(N__51505),
            .lcout(),
            .ltout(n14482_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12806_4_lut_LC_16_21_4.C_ON=1'b0;
    defparam i12806_4_lut_LC_16_21_4.SEQ_MODE=4'b0000;
    defparam i12806_4_lut_LC_16_21_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12806_4_lut_LC_16_21_4 (
            .in0(N__52322),
            .in1(N__52195),
            .in2(N__51153),
            .in3(N__51609),
            .lcout(n1257),
            .ltout(n1257_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i840_3_lut_LC_16_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i840_3_lut_LC_16_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i840_3_lut_LC_16_21_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i840_3_lut_LC_16_21_5 (
            .in0(_gnd_net_),
            .in1(N__51150),
            .in2(N__51141),
            .in3(N__51668),
            .lcout(n1328),
            .ltout(n1328_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_175_LC_16_21_6.C_ON=1'b0;
    defparam i1_4_lut_adj_175_LC_16_21_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_175_LC_16_21_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_175_LC_16_21_6 (
            .in0(N__51118),
            .in1(N__51682),
            .in2(N__51102),
            .in3(N__51091),
            .lcout(n14282),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i770_3_lut_LC_16_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i770_3_lut_LC_16_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i770_3_lut_LC_16_22_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i770_3_lut_LC_16_22_0 (
            .in0(_gnd_net_),
            .in1(N__51762),
            .in2(N__52278),
            .in3(N__51732),
            .lcout(n1226),
            .ltout(n1226_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i837_3_lut_LC_16_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i837_3_lut_LC_16_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i837_3_lut_LC_16_22_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i837_3_lut_LC_16_22_1 (
            .in0(N__51568),
            .in1(_gnd_net_),
            .in2(N__51699),
            .in3(N__51696),
            .lcout(n1325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i773_3_lut_LC_16_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i773_3_lut_LC_16_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i773_3_lut_LC_16_22_2.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i773_3_lut_LC_16_22_2 (
            .in0(N__51852),
            .in1(N__51882),
            .in2(N__52276),
            .in3(_gnd_net_),
            .lcout(n1229),
            .ltout(n1229_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_174_LC_16_22_3.C_ON=1'b0;
    defparam i1_4_lut_adj_174_LC_16_22_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_174_LC_16_22_3.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_174_LC_16_22_3 (
            .in0(N__51654),
            .in1(N__51487),
            .in2(N__51642),
            .in3(N__51639),
            .lcout(n13711),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12803_1_lut_LC_16_22_4.C_ON=1'b0;
    defparam i12803_1_lut_LC_16_22_4.SEQ_MODE=4'b0000;
    defparam i12803_1_lut_LC_16_22_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12803_1_lut_LC_16_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51567),
            .lcout(n15528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i772_3_lut_LC_16_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i772_3_lut_LC_16_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i772_3_lut_LC_16_22_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i772_3_lut_LC_16_22_6 (
            .in0(_gnd_net_),
            .in1(N__51843),
            .in2(N__52277),
            .in3(N__51813),
            .lcout(n1228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i774_3_lut_LC_16_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i774_3_lut_LC_16_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i774_3_lut_LC_16_22_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i774_3_lut_LC_16_22_7 (
            .in0(_gnd_net_),
            .in1(N__51920),
            .in2(N__51894),
            .in3(N__52264),
            .lcout(n1230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_16_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_16_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_16_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_2_lut_LC_16_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51468),
            .in3(N__51432),
            .lcout(n1201),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(n12508),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_16_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_16_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_16_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_3_lut_LC_16_23_1 (
            .in0(_gnd_net_),
            .in1(N__52894),
            .in2(N__51428),
            .in3(N__51960),
            .lcout(n1200),
            .ltout(),
            .carryin(n12508),
            .carryout(n12509),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_16_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_16_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_16_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_4_lut_LC_16_23_2 (
            .in0(_gnd_net_),
            .in1(N__51957),
            .in2(_gnd_net_),
            .in3(N__51927),
            .lcout(n1199),
            .ltout(),
            .carryin(n12509),
            .carryout(n12510),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_16_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_16_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_16_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_5_lut_LC_16_23_3 (
            .in0(_gnd_net_),
            .in1(N__52895),
            .in2(N__51924),
            .in3(N__51885),
            .lcout(n1198),
            .ltout(),
            .carryin(n12510),
            .carryout(n12511),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_16_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_16_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_16_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_6_lut_LC_16_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51881),
            .in3(N__51846),
            .lcout(n1197),
            .ltout(),
            .carryin(n12511),
            .carryout(n12512),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_16_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_16_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_16_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_7_lut_LC_16_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51842),
            .in3(N__51807),
            .lcout(n1196),
            .ltout(),
            .carryin(n12512),
            .carryout(n12513),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_16_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_16_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_16_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_8_lut_LC_16_23_6 (
            .in0(_gnd_net_),
            .in1(N__52897),
            .in2(N__51804),
            .in3(N__51765),
            .lcout(n1195),
            .ltout(),
            .carryin(n12513),
            .carryout(n12514),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_16_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_16_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_16_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_9_lut_LC_16_23_7 (
            .in0(_gnd_net_),
            .in1(N__52896),
            .in2(N__51761),
            .in3(N__51726),
            .lcout(n1194),
            .ltout(),
            .carryin(n12514),
            .carryout(n12515),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_16_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_16_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_16_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_10_lut_LC_16_24_0 (
            .in0(_gnd_net_),
            .in1(N__52892),
            .in2(N__52305),
            .in3(N__51723),
            .lcout(n1193),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(n12516),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_16_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_16_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_16_24_1.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_766_11_lut_LC_16_24_1 (
            .in0(N__52893),
            .in1(N__52355),
            .in2(N__52344),
            .in3(N__52326),
            .lcout(n1224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i769_3_lut_LC_16_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i769_3_lut_LC_16_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i769_3_lut_LC_16_24_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i769_3_lut_LC_16_24_6 (
            .in0(N__52304),
            .in1(_gnd_net_),
            .in2(N__52287),
            .in3(N__52274),
            .lcout(n1225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9618_4_lut_LC_16_25_0.C_ON=1'b0;
    defparam i9618_4_lut_LC_16_25_0.SEQ_MODE=4'b0000;
    defparam i9618_4_lut_LC_16_25_0.LUT_INIT=16'b1000000011111111;
    LogicCell40 i9618_4_lut_LC_16_25_0 (
            .in0(N__52170),
            .in1(N__54714),
            .in2(N__52161),
            .in3(N__54762),
            .lcout(direction_N_342),
            .ltout(direction_N_342_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_303_i1_3_lut_LC_16_25_1.C_ON=1'b0;
    defparam mux_303_i1_3_lut_LC_16_25_1.SEQ_MODE=4'b0000;
    defparam mux_303_i1_3_lut_LC_16_25_1.LUT_INIT=16'b0011111100001100;
    LogicCell40 mux_303_i1_3_lut_LC_16_25_1 (
            .in0(_gnd_net_),
            .in1(N__52033),
            .in2(N__52149),
            .in3(N__52136),
            .lcout(n1693),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20_3_lut_LC_16_25_5.C_ON=1'b0;
    defparam i20_3_lut_LC_16_25_5.SEQ_MODE=4'b0000;
    defparam i20_3_lut_LC_16_25_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 i20_3_lut_LC_16_25_5 (
            .in0(N__52137),
            .in1(N__52119),
            .in2(_gnd_net_),
            .in3(N__52034),
            .lcout(),
            .ltout(n13661_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam direction_167_LC_16_25_6.C_ON=1'b0;
    defparam direction_167_LC_16_25_6.SEQ_MODE=4'b1000;
    defparam direction_167_LC_16_25_6.LUT_INIT=16'b1111110100000010;
    LogicCell40 direction_167_LC_16_25_6 (
            .in0(N__54894),
            .in1(N__54990),
            .in2(N__52113),
            .in3(N__52081),
            .lcout(direction_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55811),
            .ce(),
            .sr(_gnd_net_));
    defparam i12764_2_lut_LC_16_25_7.C_ON=1'b0;
    defparam i12764_2_lut_LC_16_25_7.SEQ_MODE=4'b0000;
    defparam i12764_2_lut_LC_16_25_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i12764_2_lut_LC_16_25_7 (
            .in0(_gnd_net_),
            .in1(N__54893),
            .in2(_gnd_net_),
            .in3(N__54986),
            .lcout(n5197),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_adj_58_LC_16_26_2.C_ON=1'b0;
    defparam i9_4_lut_adj_58_LC_16_26_2.SEQ_MODE=4'b0000;
    defparam i9_4_lut_adj_58_LC_16_26_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_adj_58_LC_16_26_2 (
            .in0(N__54944),
            .in1(N__55437),
            .in2(N__54930),
            .in3(N__55115),
            .lcout(),
            .ltout(n22_adj_705_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_59_LC_16_26_3.C_ON=1'b0;
    defparam i11_4_lut_adj_59_LC_16_26_3.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_59_LC_16_26_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_59_LC_16_26_3 (
            .in0(N__55145),
            .in1(N__54911),
            .in2(N__51972),
            .in3(N__54705),
            .lcout(n24_adj_704),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_56_LC_16_27_1.C_ON=1'b0;
    defparam i1_2_lut_adj_56_LC_16_27_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_56_LC_16_27_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_56_LC_16_27_1 (
            .in0(_gnd_net_),
            .in1(N__55466),
            .in2(_gnd_net_),
            .in3(N__55130),
            .lcout(),
            .ltout(n6_adj_582_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_57_LC_16_27_2.C_ON=1'b0;
    defparam i4_4_lut_adj_57_LC_16_27_2.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_57_LC_16_27_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 i4_4_lut_adj_57_LC_16_27_2 (
            .in0(N__55052),
            .in1(N__55415),
            .in2(N__54897),
            .in3(N__55067),
            .lcout(n14108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_16_27_6.C_ON=1'b0;
    defparam i10_4_lut_LC_16_27_6.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_16_27_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 i10_4_lut_LC_16_27_6 (
            .in0(N__54874),
            .in1(N__54834),
            .in2(N__54801),
            .in3(N__54748),
            .lcout(n24_adj_699),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_LC_16_27_7.C_ON=1'b0;
    defparam i3_2_lut_LC_16_27_7.SEQ_MODE=4'b0000;
    defparam i3_2_lut_LC_16_27_7.LUT_INIT=16'b1111111111001100;
    LogicCell40 i3_2_lut_LC_16_27_7 (
            .in0(_gnd_net_),
            .in1(N__55100),
            .in2(_gnd_net_),
            .in3(N__55451),
            .lcout(n16_adj_707),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_163_LC_16_29_7.C_ON=1'b0;
    defparam dti_163_LC_16_29_7.SEQ_MODE=4'b1000;
    defparam dti_163_LC_16_29_7.LUT_INIT=16'b1111111100110011;
    LogicCell40 dti_163_LC_16_29_7 (
            .in0(_gnd_net_),
            .in1(N__55030),
            .in2(_gnd_net_),
            .in3(N__54567),
            .lcout(dti),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55827),
            .ce(N__54582),
            .sr(_gnd_net_));
    defparam i12594_2_lut_LC_16_30_1.C_ON=1'b0;
    defparam i12594_2_lut_LC_16_30_1.SEQ_MODE=4'b0000;
    defparam i12594_2_lut_LC_16_30_1.LUT_INIT=16'b1111111100110011;
    LogicCell40 i12594_2_lut_LC_16_30_1 (
            .in0(_gnd_net_),
            .in1(N__55028),
            .in2(_gnd_net_),
            .in3(N__54565),
            .lcout(),
            .ltout(dti_N_333_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_16_30_2.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_16_30_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_16_30_2.LUT_INIT=16'b1111111101101111;
    LogicCell40 i1_2_lut_4_lut_LC_16_30_2 (
            .in0(N__54697),
            .in1(N__56126),
            .in2(N__54642),
            .in3(N__54635),
            .lcout(n5169),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9550_1_lut_2_lut_LC_16_30_3.C_ON=1'b0;
    defparam i9550_1_lut_2_lut_LC_16_30_3.SEQ_MODE=4'b0000;
    defparam i9550_1_lut_2_lut_LC_16_30_3.LUT_INIT=16'b0011001111111111;
    LogicCell40 i9550_1_lut_2_lut_LC_16_30_3 (
            .in0(_gnd_net_),
            .in1(N__55027),
            .in2(_gnd_net_),
            .in3(N__54564),
            .lcout(n1377),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12554_4_lut_LC_16_31_6.C_ON=1'b0;
    defparam i12554_4_lut_LC_16_31_6.SEQ_MODE=4'b0000;
    defparam i12554_4_lut_LC_16_31_6.LUT_INIT=16'b1111011100000111;
    LogicCell40 i12554_4_lut_LC_16_31_6 (
            .in0(N__55951),
            .in1(N__56013),
            .in2(N__55035),
            .in3(N__54566),
            .lcout(n5183),
            .ltout(n5183_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3262_2_lut_LC_16_31_7.C_ON=1'b0;
    defparam i3262_2_lut_LC_16_31_7.SEQ_MODE=4'b0000;
    defparam i3262_2_lut_LC_16_31_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i3262_2_lut_LC_16_31_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__55038),
            .in3(N__55034),
            .lcout(n5235),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_3_lut_LC_17_25_4.C_ON=1'b0;
    defparam i7_3_lut_LC_17_25_4.SEQ_MODE=4'b0000;
    defparam i7_3_lut_LC_17_25_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i7_3_lut_LC_17_25_4 (
            .in0(N__54974),
            .in1(N__54959),
            .in2(_gnd_net_),
            .in3(N__55160),
            .lcout(),
            .ltout(n20_adj_706_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_LC_17_25_5.C_ON=1'b0;
    defparam i12_4_lut_LC_17_25_5.SEQ_MODE=4'b0000;
    defparam i12_4_lut_LC_17_25_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_LC_17_25_5 (
            .in0(N__55175),
            .in1(N__55086),
            .in2(N__54999),
            .in3(N__54996),
            .lcout(n13187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sweep_counter_657_658__i1_LC_17_26_0.C_ON=1'b1;
    defparam sweep_counter_657_658__i1_LC_17_26_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i1_LC_17_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i1_LC_17_26_0 (
            .in0(_gnd_net_),
            .in1(N__54975),
            .in2(_gnd_net_),
            .in3(N__54963),
            .lcout(sweep_counter_0),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(n12999),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i2_LC_17_26_1.C_ON=1'b1;
    defparam sweep_counter_657_658__i2_LC_17_26_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i2_LC_17_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i2_LC_17_26_1 (
            .in0(_gnd_net_),
            .in1(N__54960),
            .in2(_gnd_net_),
            .in3(N__54948),
            .lcout(sweep_counter_1),
            .ltout(),
            .carryin(n12999),
            .carryout(n13000),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i3_LC_17_26_2.C_ON=1'b1;
    defparam sweep_counter_657_658__i3_LC_17_26_2.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i3_LC_17_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i3_LC_17_26_2 (
            .in0(_gnd_net_),
            .in1(N__54945),
            .in2(_gnd_net_),
            .in3(N__54933),
            .lcout(sweep_counter_2),
            .ltout(),
            .carryin(n13000),
            .carryout(n13001),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i4_LC_17_26_3.C_ON=1'b1;
    defparam sweep_counter_657_658__i4_LC_17_26_3.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i4_LC_17_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i4_LC_17_26_3 (
            .in0(_gnd_net_),
            .in1(N__54929),
            .in2(_gnd_net_),
            .in3(N__54915),
            .lcout(sweep_counter_3),
            .ltout(),
            .carryin(n13001),
            .carryout(n13002),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i5_LC_17_26_4.C_ON=1'b1;
    defparam sweep_counter_657_658__i5_LC_17_26_4.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i5_LC_17_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i5_LC_17_26_4 (
            .in0(_gnd_net_),
            .in1(N__54912),
            .in2(_gnd_net_),
            .in3(N__54900),
            .lcout(sweep_counter_4),
            .ltout(),
            .carryin(n13002),
            .carryout(n13003),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i6_LC_17_26_5.C_ON=1'b1;
    defparam sweep_counter_657_658__i6_LC_17_26_5.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i6_LC_17_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i6_LC_17_26_5 (
            .in0(_gnd_net_),
            .in1(N__55176),
            .in2(_gnd_net_),
            .in3(N__55164),
            .lcout(sweep_counter_5),
            .ltout(),
            .carryin(n13003),
            .carryout(n13004),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i7_LC_17_26_6.C_ON=1'b1;
    defparam sweep_counter_657_658__i7_LC_17_26_6.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i7_LC_17_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i7_LC_17_26_6 (
            .in0(_gnd_net_),
            .in1(N__55161),
            .in2(_gnd_net_),
            .in3(N__55149),
            .lcout(sweep_counter_6),
            .ltout(),
            .carryin(n13004),
            .carryout(n13005),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i8_LC_17_26_7.C_ON=1'b1;
    defparam sweep_counter_657_658__i8_LC_17_26_7.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i8_LC_17_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i8_LC_17_26_7 (
            .in0(_gnd_net_),
            .in1(N__55146),
            .in2(_gnd_net_),
            .in3(N__55134),
            .lcout(sweep_counter_7),
            .ltout(),
            .carryin(n13005),
            .carryout(n13006),
            .clk(N__55822),
            .ce(),
            .sr(N__55400));
    defparam sweep_counter_657_658__i9_LC_17_27_0.C_ON=1'b1;
    defparam sweep_counter_657_658__i9_LC_17_27_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i9_LC_17_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i9_LC_17_27_0 (
            .in0(_gnd_net_),
            .in1(N__55131),
            .in2(_gnd_net_),
            .in3(N__55119),
            .lcout(sweep_counter_8),
            .ltout(),
            .carryin(bfn_17_27_0_),
            .carryout(n13007),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i10_LC_17_27_1.C_ON=1'b1;
    defparam sweep_counter_657_658__i10_LC_17_27_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i10_LC_17_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i10_LC_17_27_1 (
            .in0(_gnd_net_),
            .in1(N__55116),
            .in2(_gnd_net_),
            .in3(N__55104),
            .lcout(sweep_counter_9),
            .ltout(),
            .carryin(n13007),
            .carryout(n13008),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i11_LC_17_27_2.C_ON=1'b1;
    defparam sweep_counter_657_658__i11_LC_17_27_2.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i11_LC_17_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i11_LC_17_27_2 (
            .in0(_gnd_net_),
            .in1(N__55101),
            .in2(_gnd_net_),
            .in3(N__55089),
            .lcout(sweep_counter_10),
            .ltout(),
            .carryin(n13008),
            .carryout(n13009),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i12_LC_17_27_3.C_ON=1'b1;
    defparam sweep_counter_657_658__i12_LC_17_27_3.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i12_LC_17_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i12_LC_17_27_3 (
            .in0(_gnd_net_),
            .in1(N__55085),
            .in2(_gnd_net_),
            .in3(N__55071),
            .lcout(sweep_counter_11),
            .ltout(),
            .carryin(n13009),
            .carryout(n13010),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i13_LC_17_27_4.C_ON=1'b1;
    defparam sweep_counter_657_658__i13_LC_17_27_4.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i13_LC_17_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i13_LC_17_27_4 (
            .in0(_gnd_net_),
            .in1(N__55068),
            .in2(_gnd_net_),
            .in3(N__55056),
            .lcout(sweep_counter_12),
            .ltout(),
            .carryin(n13010),
            .carryout(n13011),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i14_LC_17_27_5.C_ON=1'b1;
    defparam sweep_counter_657_658__i14_LC_17_27_5.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i14_LC_17_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i14_LC_17_27_5 (
            .in0(_gnd_net_),
            .in1(N__55053),
            .in2(_gnd_net_),
            .in3(N__55041),
            .lcout(sweep_counter_13),
            .ltout(),
            .carryin(n13011),
            .carryout(n13012),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i15_LC_17_27_6.C_ON=1'b1;
    defparam sweep_counter_657_658__i15_LC_17_27_6.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i15_LC_17_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i15_LC_17_27_6 (
            .in0(_gnd_net_),
            .in1(N__55467),
            .in2(_gnd_net_),
            .in3(N__55455),
            .lcout(sweep_counter_14),
            .ltout(),
            .carryin(n13012),
            .carryout(n13013),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i16_LC_17_27_7.C_ON=1'b1;
    defparam sweep_counter_657_658__i16_LC_17_27_7.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i16_LC_17_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i16_LC_17_27_7 (
            .in0(_gnd_net_),
            .in1(N__55452),
            .in2(_gnd_net_),
            .in3(N__55440),
            .lcout(sweep_counter_15),
            .ltout(),
            .carryin(n13013),
            .carryout(n13014),
            .clk(N__55825),
            .ce(),
            .sr(N__55401));
    defparam sweep_counter_657_658__i17_LC_17_28_0.C_ON=1'b1;
    defparam sweep_counter_657_658__i17_LC_17_28_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i17_LC_17_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i17_LC_17_28_0 (
            .in0(_gnd_net_),
            .in1(N__55436),
            .in2(_gnd_net_),
            .in3(N__55422),
            .lcout(sweep_counter_16),
            .ltout(),
            .carryin(bfn_17_28_0_),
            .carryout(n13015),
            .clk(N__55828),
            .ce(),
            .sr(N__55403));
    defparam sweep_counter_657_658__i18_LC_17_28_1.C_ON=1'b0;
    defparam sweep_counter_657_658__i18_LC_17_28_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_657_658__i18_LC_17_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_657_658__i18_LC_17_28_1 (
            .in0(_gnd_net_),
            .in1(N__55416),
            .in2(_gnd_net_),
            .in3(N__55419),
            .lcout(sweep_counter_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55828),
            .ce(),
            .sr(N__55403));
    defparam dir_160_LC_17_32_2.C_ON=1'b0;
    defparam dir_160_LC_17_32_2.SEQ_MODE=4'b1000;
    defparam dir_160_LC_17_32_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 dir_160_LC_17_32_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55335),
            .lcout(dir),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55832),
            .ce(),
            .sr(_gnd_net_));
    defparam GHB_172_LC_18_31_5.C_ON=1'b0;
    defparam GHB_172_LC_18_31_5.SEQ_MODE=4'b1000;
    defparam GHB_172_LC_18_31_5.LUT_INIT=16'b1100110000100001;
    LogicCell40 GHB_172_LC_18_31_5 (
            .in0(N__56147),
            .in1(N__56036),
            .in2(N__55968),
            .in3(N__55881),
            .lcout(GHB),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55833),
            .ce(N__55633),
            .sr(N__55592));
    defparam GHA_170_LC_18_32_4.C_ON=1'b0;
    defparam GHA_170_LC_18_32_4.SEQ_MODE=4'b1000;
    defparam GHA_170_LC_18_32_4.LUT_INIT=16'b0000001110011000;
    LogicCell40 GHA_170_LC_18_32_4 (
            .in0(N__56148),
            .in1(N__56030),
            .in2(N__55962),
            .in3(N__55872),
            .lcout(GHA),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55834),
            .ce(N__55638),
            .sr(N__55590));
    defparam GLB_173_LC_19_31_1.C_ON=1'b0;
    defparam GLB_173_LC_19_31_1.SEQ_MODE=4'b1000;
    defparam GLB_173_LC_19_31_1.LUT_INIT=16'b0000100111110000;
    LogicCell40 GLB_173_LC_19_31_1 (
            .in0(N__56144),
            .in1(N__55964),
            .in2(N__56046),
            .in3(N__55890),
            .lcout(INLB_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55835),
            .ce(N__55629),
            .sr(N__55596));
    defparam GHC_174_LC_19_31_3.C_ON=1'b0;
    defparam GHC_174_LC_19_31_3.SEQ_MODE=4'b1000;
    defparam GHC_174_LC_19_31_3.LUT_INIT=16'b1100110001010010;
    LogicCell40 GHC_174_LC_19_31_3 (
            .in0(N__56143),
            .in1(N__55963),
            .in2(N__56045),
            .in3(N__55889),
            .lcout(GHC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55835),
            .ce(N__55629),
            .sr(N__55596));
    defparam GLA_171_LC_19_32_0.C_ON=1'b0;
    defparam GLA_171_LC_19_32_0.SEQ_MODE=4'b1000;
    defparam GLA_171_LC_19_32_0.LUT_INIT=16'b1001100000000011;
    LogicCell40 GLA_171_LC_19_32_0 (
            .in0(N__56146),
            .in1(N__56043),
            .in2(N__55961),
            .in3(N__55882),
            .lcout(INLA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55836),
            .ce(N__55637),
            .sr(N__55591));
    defparam GLC_175_LC_19_32_2.C_ON=1'b0;
    defparam GLC_175_LC_19_32_2.SEQ_MODE=4'b1000;
    defparam GLC_175_LC_19_32_2.LUT_INIT=16'b0100011011110000;
    LogicCell40 GLC_175_LC_19_32_2 (
            .in0(N__56145),
            .in1(N__56044),
            .in2(N__55960),
            .in3(N__55883),
            .lcout(INLC_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55836),
            .ce(N__55637),
            .sr(N__55591));
    defparam i9540_2_lut_LC_20_31_3.C_ON=1'b0;
    defparam i9540_2_lut_LC_20_31_3.SEQ_MODE=4'b0000;
    defparam i9540_2_lut_LC_20_31_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9540_2_lut_LC_20_31_3 (
            .in0(N__55504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55557),
            .lcout(INHB_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9541_2_lut_LC_20_31_4.C_ON=1'b0;
    defparam i9541_2_lut_LC_20_31_4.SEQ_MODE=4'b0000;
    defparam i9541_2_lut_LC_20_31_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9541_2_lut_LC_20_31_4 (
            .in0(N__55533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55505),
            .lcout(INHC_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9539_2_lut_LC_20_32_3.C_ON=1'b0;
    defparam i9539_2_lut_LC_20_32_3.SEQ_MODE=4'b0000;
    defparam i9539_2_lut_LC_20_32_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9539_2_lut_LC_20_32_3 (
            .in0(N__55512),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55488),
            .lcout(INHA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
