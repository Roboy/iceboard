// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Jan  6 14:15:37 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    output SCL;   // verilog/TinyFPGA_B.v(21[10:13])
    input SDA /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c_0;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(42[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(88[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(89[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(125[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(126[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(127[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(128[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(129[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(131[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(132[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(133[22:35])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(163[22:33])
    wire [22:0]pwm_setpoint_22__N_3;
    
    wire RX_N_2;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n1138;
    wire [23:0]displacement_23__N_26;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    wire [3:0]state_3__N_372;
    
    wire n4727, n4725, n15784, n15783, n15782, n15781, n15780, 
        n15779, n15778, n27243, n15777, n15776;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n5, n15775, n15774, n15773, n15772, n15771, n3, n4, 
        n5_adj_4758, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
        n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
        n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n15770, n15769, n122, n123, n7_adj_4759, n6_adj_4760, n771, 
        n10_adj_4761, n15768, n15767, n15766, n23506, n23505, n23504, 
        n14328, n23503, n23502, n23501, n23500, n23499, n4_adj_4762, 
        n23498, n23497, n23496, n23495, n23494, n23493, n23492, 
        n23491, n23490, n23489, n23488, n23487, n23486, n23485, 
        n19238, n15765, n15764, n3303;
    wire [31:0]\FRAME_MATCHER.state_31__N_2668 ;
    
    wire n15761, n15760, n15759, n15758, n15757, n15756, n15755, 
        n15754, n15753, n15752, n15751, n15750, n15749, n15748, 
        n15747, n15746, n15745, n15744, n15743, n15742, n15741, 
        n15740, n15739, n4452, n14282, n16247, n16246, n16245, 
        n16244, n16243, n16242, n16241, n16239, n16237, n16232, 
        n16231, n16230, n16229, n16228, n16227, n16226, n16225, 
        n16224, n16223, n16222, n16221, n16220, n16219, n16218, 
        n16217, n16216, n16215, n16214, n16213, n16212, n16211, 
        n16210, n16209, n16208, n16207, n16206, n16205, n16204, 
        n16203, n16199, n63, n4_adj_4763, n16023, n16022, n16021, 
        n16020, n16019, n16018, n16017, n16016, n16015, n16014, 
        n16013, n16012, n16011, n16010, n16009, n16008, n16007, 
        n6_adj_4764, n7_adj_4765, n8_adj_4766, n9_adj_4767, n10_adj_4768, 
        n11_adj_4769, n12_adj_4770, n13_adj_4771, n14_adj_4772, n15_adj_4773, 
        n16_adj_4774, n17_adj_4775, n18_adj_4776, n19_adj_4777, n20_adj_4778, 
        n21_adj_4779, n22_adj_4780, n23_adj_4781, n24_adj_4782, n25_adj_4783, 
        n16006, n16005, n23722, n16004, n16003, n16002, n16001, 
        n16000, n15548, n15999, n23721, n15998, n15997, n15996, 
        n15995, n15994, n23720, n15993, n15992, n15991, n15990, 
        n15989, n15988, n15987, n15986, n15985, n15984, n15983, 
        n15982, n15981, n15980, n15979, n15978, n15977, n15976, 
        n15975, n15974, n15973, n15972, n15971, n15970, n15969, 
        n15968, n15643, n15967, n15966, n15965, n15964, n15963, 
        n15962, n15961, n15960, n15959, n15958, n15957, n15956, 
        n15955, n15488, n4_adj_4784, n15954, n15953, n15952, n15951, 
        n15950, n15949, n15948, n15947, n15946, n15945, n15944, 
        n15943, n15942, n15941, n15940, n15939, n15938, n15937, 
        n15936, n15935, n15934, n15933, n15932, n15931, n15930, 
        quadA_debounced, quadB_debounced, n15451, n15929, n15928, 
        n15927, n15926, n15925, n15924, n15923, n15922, quadA_debounced_adj_4785, 
        quadB_debounced_adj_4786, n15921, n15920, n15919, n15918, 
        n15917, n15916, n15915, n15914, n15913, n15912, n15911, 
        n15910, n15909, n15908, n15907, n15906, n15905, n15904, 
        n15903, n15902, n15901, n15900, n15899, n15898, n15897, 
        n15896, n15895, n15894, n15893, n15892, n15891, n15890, 
        n15889, n15888, n15887, n15886, n4_adj_4787, n15885, n15884, 
        n15883, n15882, n63_adj_4788, n15881, n23719, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n4_adj_4789, n15880, n3_adj_4790, n15879;
    wire [2:0]r_SM_Main_2__N_3422;
    
    wire n15878, n15877, n15876, n15738, n15875, n15874, n15873, 
        n15872, n15871, n15870, n15869, n15868, n15867, n15866, 
        n15865, n15864;
    wire [2:0]r_SM_Main_adj_4867;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_4869;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3493;
    
    wire n2, n15863, n15862, n15861, n15860, n15859, n15858, n15857, 
        n15856, n15855, n15854, n15853, n15852, n15851, n15850, 
        n15849, n15848, n15847, n15846;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n5_adj_4795, n15845;
    wire [1:0]reg_B_adj_4879;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15844, n15843, n31935, n31149, n31148, n31147, n31146, 
        n31145, n1, n31144, n31143, n31142, n31141, n31140, n23718, 
        n31139, n31138, n31137, n31136, n23717, n31135, n31134, 
        n31133, n31132, n31131, n31130, n5_adj_4798, n31129, n31128, 
        n31127, n23716, n32553, n15737, n15736, n15735, n15734, 
        n15733, n15732, n15731, n15730, n15842, n15841, n15840, 
        n15839, n15838, n15837, n15836, n15835, n15834, n15833, 
        n15832, n15831, n15830, n15829, n15828, n15827, n15826, 
        n15825, n15824, n15823, n15822, n15821, n15820, n15819, 
        n15818, n15817, n15815, n15814, n15813, n15812, n15811, 
        n15810, n15809, n15726, n15724, n15723, n15722, n15721, 
        n15719, n15807, n15806, n15805, n15804, n15803, n15802, 
        n15801, n15800, n15718, n15716, n15715, n15714, n15713, 
        n15712, n15711, n15710, n15799, n15798, n15797, n15796, 
        n15795, n15794, n15793, n15792, n15791, n15790, n15789, 
        n15788, n15787, n15786, n15785, n30266, n27831, n28731, 
        n29426, n26593, n14318, n14295, n14309, n31082, n29773, 
        n31069, n28775, n8515, n27820, n27405, n23715, n15709, 
        n15708, n28749, n32898, n1_adj_4799, n1_adj_4800, n1_adj_4801, 
        n1_adj_4802, n1_adj_4803, n1_adj_4804, n1_adj_4805, n1_adj_4806, 
        n1_adj_4807, n1_adj_4808, n1_adj_4809, n1_adj_4810, n1_adj_4811, 
        n1_adj_4812, n1_adj_4813, n1_adj_4814, n1_adj_4815, n1_adj_4816, 
        n1_adj_4817, n1_adj_4818, n1_adj_4819, n1_adj_4820, n1_adj_4821, 
        n28639, n15707, n15706, n15705, n15704, n30290, n23714, 
        n23_adj_4822, n23713, n28597, n30174, n29458, n14287, n27755, 
        n11643, n29573, n6_adj_4823, n32532, n8_adj_4824, n32531, 
        n26505, n8353, n23712, n23711, n23710, n23709, n23708, 
        n23707, n23706, n23705, n23704, n23703, n23702, n23701, 
        n23700;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced, 
            quadB_debounced}), .reg_B({reg_B}), .n30174(n30174), .ENCODER0_B_c_0(ENCODER0_B_c_0), 
            .n16237(n16237), .ENCODER0_A_c_1(ENCODER0_A_c_1), .n15721(n15721)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(187[15] 192[4])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_40 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF h2_39 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i25551_2_lut (.I0(displacement[13]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31137));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25551_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_13_i1_3_lut (.I0(encoder0_position[13]), .I1(encoder1_position[13]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4809));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_13_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11195_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n26593), .I3(GND_net), .O(n15734));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11195_3_lut.LUT_INIT = 16'hacac;
    neopixel nx (.GND_net(GND_net), .timer({timer}), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .\state[1] (state[1]), .start(start), 
            .n28731(n28731), .n26593(n26593), .VCC_net(VCC_net), .n28597(n28597), 
            .n15451(n15451), .\state_3__N_372[1] (state_3__N_372[1]), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .neopxl_color({neopxl_color}), .LED_c(LED_c), .NEOPXL_c(NEOPXL_c), 
            .n15761(n15761), .n15760(n15760), .n15759(n15759), .n15758(n15758), 
            .n15757(n15757), .n15756(n15756), .n15755(n15755), .n15754(n15754), 
            .n15753(n15753), .n15752(n15752), .n15751(n15751), .n15750(n15750), 
            .n15749(n15749), .n15748(n15748), .n15747(n15747), .n15746(n15746), 
            .n15745(n15745), .n15744(n15744), .n15743(n15743), .n15742(n15742), 
            .n15741(n15741), .n15740(n15740), .n15739(n15739), .n15738(n15738), 
            .n15737(n15737), .n15736(n15736), .n15735(n15735), .n15734(n15734), 
            .n15733(n15733), .n15732(n15732), .n15731(n15731), .n26505(n26505), 
            .n29426(n29426), .n15726(n15726), .n15704(n15704)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(44[10] 50[2])
    SB_LUT4 i11278_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15817));   // verilog/coms.v(127[12] 300[6])
    defparam i11278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14742_4_lut (.I0(n1_adj_4809), .I1(n29773), .I2(n31137), 
            .I3(control_mode[1]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14742_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11196_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n26593), .I3(GND_net), .O(n15735));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11197_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n26593), .I3(GND_net), .O(n15736));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11279_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15818));   // verilog/coms.v(127[12] 300[6])
    defparam i11279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11198_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n26593), .I3(GND_net), .O(n15737));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11280_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n29573), 
            .I3(GND_net), .O(n15819));   // verilog/coms.v(127[12] 300[6])
    defparam i11280_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11281_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n29573), 
            .I3(GND_net), .O(n15820));   // verilog/coms.v(127[12] 300[6])
    defparam i11281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11199_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n26593), .I3(GND_net), .O(n15738));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11282_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n29573), 
            .I3(GND_net), .O(n15821));   // verilog/coms.v(127[12] 300[6])
    defparam i11282_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11200_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n26593), .I3(GND_net), .O(n15739));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11200_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dir_44 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_LUT4 i11201_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n26593), .I3(GND_net), .O(n15740));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11201_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11283_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n29573), 
            .I3(GND_net), .O(n15822));   // verilog/coms.v(127[12] 300[6])
    defparam i11283_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11202_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n26593), .I3(GND_net), .O(n15741));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11202_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11203_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n26593), .I3(GND_net), .O(n15742));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11284_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n29573), 
            .I3(GND_net), .O(n15823));   // verilog/coms.v(127[12] 300[6])
    defparam i11284_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11204_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n26593), .I3(GND_net), .O(n15743));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i25550_2_lut (.I0(displacement[14]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31136));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25550_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_14_i1_3_lut (.I0(encoder0_position[14]), .I1(encoder1_position[14]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4808));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14741_4_lut (.I0(n1_adj_4808), .I1(n29773), .I2(n31136), 
            .I3(control_mode[1]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14741_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11285_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n29573), 
            .I3(GND_net), .O(n15824));   // verilog/coms.v(127[12] 300[6])
    defparam i11285_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11205_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n26593), .I3(GND_net), .O(n15744));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11206_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n26593), .I3(GND_net), .O(n15745));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11286_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n29573), 
            .I3(GND_net), .O(n15825));   // verilog/coms.v(127[12] 300[6])
    defparam i11286_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11207_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n26593), .I3(GND_net), .O(n15746));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11208_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n26593), .I3(GND_net), .O(n15747));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11287_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n29573), 
            .I3(GND_net), .O(n15826));   // verilog/coms.v(127[12] 300[6])
    defparam i11287_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11209_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n26593), .I3(GND_net), .O(n15748));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11210_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n26593), .I3(GND_net), .O(n15749));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11211_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n26593), .I3(GND_net), .O(n15750));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11212_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n26593), .I3(GND_net), .O(n15751));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4781));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11213_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n26593), .I3(GND_net), .O(n15752));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4780));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11214_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n26593), .I3(GND_net), .O(n15753));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4779));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11288_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n29573), 
            .I3(GND_net), .O(n15827));   // verilog/coms.v(127[12] 300[6])
    defparam i11288_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11215_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n26593), .I3(GND_net), .O(n15754));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11216_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n26593), .I3(GND_net), .O(n15755));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11289_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n29573), 
            .I3(GND_net), .O(n15828));   // verilog/coms.v(127[12] 300[6])
    defparam i11289_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11217_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n26593), .I3(GND_net), .O(n15756));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11290_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n29573), 
            .I3(GND_net), .O(n15829));   // verilog/coms.v(127[12] 300[6])
    defparam i11290_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11218_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n26593), .I3(GND_net), .O(n15757));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11219_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n26593), .I3(GND_net), .O(n15758));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11291_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n29573), 
            .I3(GND_net), .O(n15830));   // verilog/coms.v(127[12] 300[6])
    defparam i11291_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11220_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n26593), .I3(GND_net), .O(n15759));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11221_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n26593), .I3(GND_net), .O(n15760));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11292_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n29573), 
            .I3(GND_net), .O(n15831));   // verilog/coms.v(127[12] 300[6])
    defparam i11292_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11293_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n29573), 
            .I3(GND_net), .O(n15832));   // verilog/coms.v(127[12] 300[6])
    defparam i11293_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11294_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n29573), 
            .I3(GND_net), .O(n15833));   // verilog/coms.v(127[12] 300[6])
    defparam i11294_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11295_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n29573), 
            .I3(GND_net), .O(n15834));   // verilog/coms.v(127[12] 300[6])
    defparam i11295_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11296_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n29573), 
            .I3(GND_net), .O(n15835));   // verilog/coms.v(127[12] 300[6])
    defparam i11296_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11297_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n29573), 
            .I3(GND_net), .O(n15836));   // verilog/coms.v(127[12] 300[6])
    defparam i11297_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11298_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n29573), 
            .I3(GND_net), .O(n15837));   // verilog/coms.v(127[12] 300[6])
    defparam i11298_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11299_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n29573), 
            .I3(GND_net), .O(n15838));   // verilog/coms.v(127[12] 300[6])
    defparam i11299_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4778));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11300_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n29573), 
            .I3(GND_net), .O(n15839));   // verilog/coms.v(127[12] 300[6])
    defparam i11300_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4777));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14751_4_lut (.I0(n1_adj_4818), .I1(n29773), .I2(n31146), 
            .I3(control_mode[1]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14751_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11222_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n26593), .I3(GND_net), .O(n15761));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4766));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4776));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25559_2_lut (.I0(displacement[5]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31145));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25559_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_5_i1_3_lut (.I0(encoder0_position[5]), .I1(encoder1_position[5]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4817));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_5_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4765));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4775));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11301_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n29573), 
            .I3(GND_net), .O(n15840));   // verilog/coms.v(127[12] 300[6])
    defparam i11301_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11302_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n29573), 
            .I3(GND_net), .O(n15841));   // verilog/coms.v(127[12] 300[6])
    defparam i11302_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4764));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11226_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n4725), .I3(GND_net), .O(n15765));   // verilog/coms.v(127[12] 300[6])
    defparam i11226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11227_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n4725), .I3(GND_net), .O(n15766));   // verilog/coms.v(127[12] 300[6])
    defparam i11227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11303_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n29573), 
            .I3(GND_net), .O(n15842));   // verilog/coms.v(127[12] 300[6])
    defparam i11303_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11304_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n29573), 
            .I3(GND_net), .O(n15843));   // verilog/coms.v(127[12] 300[6])
    defparam i11304_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11305_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n29573), 
            .I3(GND_net), .O(n15844));   // verilog/coms.v(127[12] 300[6])
    defparam i11305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11306_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n29573), 
            .I3(GND_net), .O(n15845));   // verilog/coms.v(127[12] 300[6])
    defparam i11306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11307_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n29573), 
            .I3(GND_net), .O(n15846));   // verilog/coms.v(127[12] 300[6])
    defparam i11307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11308_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n29573), 
            .I3(GND_net), .O(n15847));   // verilog/coms.v(127[12] 300[6])
    defparam i11308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11309_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n29573), 
            .I3(GND_net), .O(n15848));   // verilog/coms.v(127[12] 300[6])
    defparam i11309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11310_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n11643), .I3(GND_net), .O(n15849));   // verilog/coms.v(127[12] 300[6])
    defparam i11310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11311_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n11643), .I3(GND_net), .O(n15850));   // verilog/coms.v(127[12] 300[6])
    defparam i11311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11312_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n11643), .I3(GND_net), .O(n15851));   // verilog/coms.v(127[12] 300[6])
    defparam i11312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11313_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n11643), .I3(GND_net), .O(n15852));   // verilog/coms.v(127[12] 300[6])
    defparam i11313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11314_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n11643), .I3(GND_net), .O(n15853));   // verilog/coms.v(127[12] 300[6])
    defparam i11314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11315_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n11643), .I3(GND_net), .O(n15854));   // verilog/coms.v(127[12] 300[6])
    defparam i11315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11165_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n26593), .I3(GND_net), .O(n15704));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11165_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11166_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n4725), .I3(GND_net), .O(n15705));   // verilog/coms.v(127[12] 300[6])
    defparam i11166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11167_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n19238), 
            .I3(n14287), .O(n15706));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11167_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i11168_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n19238), 
            .I3(n14282), .O(n15707));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11168_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4789));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11169_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4784), 
            .I3(n14287), .O(n15708));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11169_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11170_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4784), 
            .I3(n14282), .O(n15709));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11170_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11171_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4787), 
            .I3(n14287), .O(n15710));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11171_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11172_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4787), 
            .I3(n14282), .O(n15711));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11172_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11316_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n11643), .I3(GND_net), .O(n15855));   // verilog/coms.v(127[12] 300[6])
    defparam i11316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11317_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n11643), .I3(GND_net), .O(n15856));   // verilog/coms.v(127[12] 300[6])
    defparam i11317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14750_4_lut (.I0(n1_adj_4817), .I1(n29773), .I2(n31145), 
            .I3(control_mode[1]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14750_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11318_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n11643), .I3(GND_net), .O(n15857));   // verilog/coms.v(127[12] 300[6])
    defparam i11318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11319_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n11643), .I3(GND_net), .O(n15858));   // verilog/coms.v(127[12] 300[6])
    defparam i11319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11320_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n11643), .I3(GND_net), .O(n15859));   // verilog/coms.v(127[12] 300[6])
    defparam i11320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11321_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n11643), .I3(GND_net), .O(n15860));   // verilog/coms.v(127[12] 300[6])
    defparam i11321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11322_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n11643), .I3(GND_net), .O(n15861));   // verilog/coms.v(127[12] 300[6])
    defparam i11322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11173_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4763), 
            .I3(n14287), .O(n15712));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11173_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11174_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15713));   // verilog/coms.v(127[12] 300[6])
    defparam i11174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11175_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n29573), 
            .I3(GND_net), .O(n15714));   // verilog/coms.v(127[12] 300[6])
    defparam i11175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11176_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n29573), 
            .I3(GND_net), .O(n15715));   // verilog/coms.v(127[12] 300[6])
    defparam i11176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11177_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n4727), .I3(GND_net), .O(n15716));   // verilog/coms.v(127[12] 300[6])
    defparam i11177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11179_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4725), .I3(GND_net), .O(n15718));   // verilog/coms.v(127[12] 300[6])
    defparam i11179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11323_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n11643), .I3(GND_net), .O(n15862));   // verilog/coms.v(127[12] 300[6])
    defparam i11323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11324_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n11643), .I3(GND_net), .O(n15863));   // verilog/coms.v(127[12] 300[6])
    defparam i11324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11325_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n11643), .I3(GND_net), .O(n15864));   // verilog/coms.v(127[12] 300[6])
    defparam i11325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11326_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n11643), .I3(GND_net), .O(n15865));   // verilog/coms.v(127[12] 300[6])
    defparam i11326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11327_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n11643), .I3(GND_net), .O(n15866));   // verilog/coms.v(127[12] 300[6])
    defparam i11327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11328_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n11643), .I3(GND_net), .O(n15867));   // verilog/coms.v(127[12] 300[6])
    defparam i11328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11329_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n11643), .I3(GND_net), .O(n15868));   // verilog/coms.v(127[12] 300[6])
    defparam i11329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11330_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n11643), .I3(GND_net), .O(n15869));   // verilog/coms.v(127[12] 300[6])
    defparam i11330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11331_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n11643), .I3(GND_net), .O(n15870));   // verilog/coms.v(127[12] 300[6])
    defparam i11331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11332_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n11643), .I3(GND_net), .O(n15871));   // verilog/coms.v(127[12] 300[6])
    defparam i11332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11333_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n11643), .I3(GND_net), .O(n15872));   // verilog/coms.v(127[12] 300[6])
    defparam i11333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11334_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n11643), .I3(GND_net), .O(n15873));   // verilog/coms.v(127[12] 300[6])
    defparam i11334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25558_2_lut (.I0(displacement[6]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31144));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25558_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11335_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n11643), .I3(GND_net), .O(n15874));   // verilog/coms.v(127[12] 300[6])
    defparam i11335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11336_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n11643), .I3(GND_net), .O(n15875));   // verilog/coms.v(127[12] 300[6])
    defparam i11336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11337_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n11643), .I3(GND_net), .O(n15876));   // verilog/coms.v(127[12] 300[6])
    defparam i11337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11338_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n11643), .I3(GND_net), .O(n15877));   // verilog/coms.v(127[12] 300[6])
    defparam i11338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11339_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n11643), .I3(GND_net), .O(n15878));   // verilog/coms.v(127[12] 300[6])
    defparam i11339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11340_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n11643), .I3(GND_net), .O(n15879));   // verilog/coms.v(127[12] 300[6])
    defparam i11340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11341_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n11643), .I3(GND_net), .O(n15880));   // verilog/coms.v(127[12] 300[6])
    defparam i11341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11228_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n4725), .I3(GND_net), .O(n15767));   // verilog/coms.v(127[12] 300[6])
    defparam i11228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11342_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n11643), .I3(GND_net), .O(n15881));   // verilog/coms.v(127[12] 300[6])
    defparam i11342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11343_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n11643), .I3(GND_net), .O(n15882));   // verilog/coms.v(127[12] 300[6])
    defparam i11343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11344_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n11643), .I3(GND_net), .O(n15883));   // verilog/coms.v(127[12] 300[6])
    defparam i11344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11345_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n11643), .I3(GND_net), .O(n15884));   // verilog/coms.v(127[12] 300[6])
    defparam i11345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_Mux_6_i1_3_lut (.I0(encoder0_position[6]), .I1(encoder1_position[6]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4816));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11346_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n11643), .I3(GND_net), .O(n15885));   // verilog/coms.v(127[12] 300[6])
    defparam i11346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11347_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n11643), .I3(GND_net), .O(n15886));   // verilog/coms.v(127[12] 300[6])
    defparam i11347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11348_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n11643), .I3(GND_net), .O(n15887));   // verilog/coms.v(127[12] 300[6])
    defparam i11348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11229_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n4725), .I3(GND_net), .O(n15768));   // verilog/coms.v(127[12] 300[6])
    defparam i11229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14749_4_lut (.I0(n1_adj_4816), .I1(n29773), .I2(n31144), 
            .I3(control_mode[1]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14749_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11349_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n11643), .I3(GND_net), .O(n15888));   // verilog/coms.v(127[12] 300[6])
    defparam i11349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11350_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n11643), .I3(GND_net), .O(n15889));   // verilog/coms.v(127[12] 300[6])
    defparam i11350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11351_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n11643), .I3(GND_net), .O(n15890));   // verilog/coms.v(127[12] 300[6])
    defparam i11351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11352_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n11643), .I3(GND_net), .O(n15891));   // verilog/coms.v(127[12] 300[6])
    defparam i11352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11353_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n11643), .I3(GND_net), .O(n15892));   // verilog/coms.v(127[12] 300[6])
    defparam i11353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11354_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n11643), .I3(GND_net), .O(n15893));   // verilog/coms.v(127[12] 300[6])
    defparam i11354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11355_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n11643), .I3(GND_net), .O(n15894));   // verilog/coms.v(127[12] 300[6])
    defparam i11355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11180_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n4725), .I3(GND_net), .O(n15719));   // verilog/coms.v(127[12] 300[6])
    defparam i11180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(n14318), .I1(n27755), .I2(n3303), .I3(n28639), 
            .O(n30266));
    defparam i2_4_lut.LUT_INIT = 16'hcdff;
    SB_LUT4 i1_4_lut (.I0(n63_adj_4788), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n30266), .I3(n30290), .O(n27243));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut.LUT_INIT = 16'hd5f5;
    SB_LUT4 i11182_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n30174), 
            .I3(GND_net), .O(n15721));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11183_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_4867[1]), .I2(n8353), 
            .I3(n4_adj_4762), .O(n15722));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11183_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i11184_3_lut (.I0(quadB_debounced_adj_4786), .I1(reg_B_adj_4879[0]), 
            .I2(n29458), .I3(GND_net), .O(n15723));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11185_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1138), .I3(GND_net), .O(n15724));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11187_4_lut (.I0(n28597), .I1(state[1]), .I2(state_3__N_372[1]), 
            .I3(n15451), .O(n15726));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11187_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4774));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4773));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4772));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11356_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n11643), .I3(GND_net), .O(n15895));   // verilog/coms.v(127[12] 300[6])
    defparam i11356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11357_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n11643), .I3(GND_net), .O(n15896));   // verilog/coms.v(127[12] 300[6])
    defparam i11357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11358_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n11643), .I3(GND_net), .O(n15897));   // verilog/coms.v(127[12] 300[6])
    defparam i11358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11359_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n11643), .I3(GND_net), .O(n15898));   // verilog/coms.v(127[12] 300[6])
    defparam i11359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11360_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n11643), .I3(GND_net), .O(n15899));   // verilog/coms.v(127[12] 300[6])
    defparam i11360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11361_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n11643), .I3(GND_net), .O(n15900));   // verilog/coms.v(127[12] 300[6])
    defparam i11361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11362_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n11643), .I3(GND_net), .O(n15901));   // verilog/coms.v(127[12] 300[6])
    defparam i11362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11363_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n11643), .I3(GND_net), .O(n15902));   // verilog/coms.v(127[12] 300[6])
    defparam i11363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11364_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n11643), .I3(GND_net), .O(n15903));   // verilog/coms.v(127[12] 300[6])
    defparam i11364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11365_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n11643), .I3(GND_net), .O(n15904));   // verilog/coms.v(127[12] 300[6])
    defparam i11365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11366_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n11643), .I3(GND_net), .O(n15905));   // verilog/coms.v(127[12] 300[6])
    defparam i11366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11367_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n11643), .I3(GND_net), .O(n15906));   // verilog/coms.v(127[12] 300[6])
    defparam i11367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11368_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n11643), .I3(GND_net), .O(n15907));   // verilog/coms.v(127[12] 300[6])
    defparam i11368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11369_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n11643), .I3(GND_net), .O(n15908));   // verilog/coms.v(127[12] 300[6])
    defparam i11369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11370_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n11643), .I3(GND_net), .O(n15909));   // verilog/coms.v(127[12] 300[6])
    defparam i11370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11371_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n11643), .I3(GND_net), .O(n15910));   // verilog/coms.v(127[12] 300[6])
    defparam i11371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11372_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n11643), .I3(GND_net), .O(n15911));   // verilog/coms.v(127[12] 300[6])
    defparam i11372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11373_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n11643), .I3(GND_net), .O(n15912));   // verilog/coms.v(127[12] 300[6])
    defparam i11373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11374_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n11643), .I3(GND_net), .O(n15913));   // verilog/coms.v(127[12] 300[6])
    defparam i11374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11375_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n11643), .I3(GND_net), .O(n15914));   // verilog/coms.v(127[12] 300[6])
    defparam i11375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11376_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n11643), .I3(GND_net), .O(n15915));   // verilog/coms.v(127[12] 300[6])
    defparam i11376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11377_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n11643), .I3(GND_net), .O(n15916));   // verilog/coms.v(127[12] 300[6])
    defparam i11377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11378_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n11643), .I3(GND_net), .O(n15917));   // verilog/coms.v(127[12] 300[6])
    defparam i11378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11379_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n11643), .I3(GND_net), .O(n15918));   // verilog/coms.v(127[12] 300[6])
    defparam i11379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11380_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n11643), .I3(GND_net), .O(n15919));   // verilog/coms.v(127[12] 300[6])
    defparam i11380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11381_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n11643), .I3(GND_net), .O(n15920));   // verilog/coms.v(127[12] 300[6])
    defparam i11381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11382_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n11643), .I3(GND_net), .O(n15921));   // verilog/coms.v(127[12] 300[6])
    defparam i11382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11383_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n11643), .I3(GND_net), .O(n15922));   // verilog/coms.v(127[12] 300[6])
    defparam i11383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11384_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n11643), .I3(GND_net), .O(n15923));   // verilog/coms.v(127[12] 300[6])
    defparam i11384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11385_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n11643), .I3(GND_net), .O(n15924));   // verilog/coms.v(127[12] 300[6])
    defparam i11385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11386_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n11643), .I3(GND_net), .O(n15925));   // verilog/coms.v(127[12] 300[6])
    defparam i11386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11387_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n11643), .I3(GND_net), .O(n15926));   // verilog/coms.v(127[12] 300[6])
    defparam i11387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11388_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n11643), .I3(GND_net), .O(n15927));   // verilog/coms.v(127[12] 300[6])
    defparam i11388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11389_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n11643), .I3(GND_net), .O(n15928));   // verilog/coms.v(127[12] 300[6])
    defparam i11389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11390_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n11643), 
            .I3(GND_net), .O(n15929));   // verilog/coms.v(127[12] 300[6])
    defparam i11390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4771));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11391_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n11643), 
            .I3(GND_net), .O(n15930));   // verilog/coms.v(127[12] 300[6])
    defparam i11391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11392_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n11643), 
            .I3(GND_net), .O(n15931));   // verilog/coms.v(127[12] 300[6])
    defparam i11392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11393_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n11643), 
            .I3(GND_net), .O(n15932));   // verilog/coms.v(127[12] 300[6])
    defparam i11393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11394_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n11643), 
            .I3(GND_net), .O(n15933));   // verilog/coms.v(127[12] 300[6])
    defparam i11394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11395_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n11643), 
            .I3(GND_net), .O(n15934));   // verilog/coms.v(127[12] 300[6])
    defparam i11395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11396_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n11643), 
            .I3(GND_net), .O(n15935));   // verilog/coms.v(127[12] 300[6])
    defparam i11396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11397_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n11643), 
            .I3(GND_net), .O(n15936));   // verilog/coms.v(127[12] 300[6])
    defparam i11397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11398_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n11643), 
            .I3(GND_net), .O(n15937));   // verilog/coms.v(127[12] 300[6])
    defparam i11398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11399_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n11643), 
            .I3(GND_net), .O(n15938));   // verilog/coms.v(127[12] 300[6])
    defparam i11399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11400_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n11643), 
            .I3(GND_net), .O(n15939));   // verilog/coms.v(127[12] 300[6])
    defparam i11400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25557_2_lut (.I0(displacement[7]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31143));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25557_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11401_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n11643), 
            .I3(GND_net), .O(n15940));   // verilog/coms.v(127[12] 300[6])
    defparam i11401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_Mux_7_i1_3_lut (.I0(encoder0_position[7]), .I1(encoder1_position[7]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4815));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_7_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11402_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n11643), 
            .I3(GND_net), .O(n15941));   // verilog/coms.v(127[12] 300[6])
    defparam i11402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25549_2_lut (.I0(displacement[15]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31135));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25549_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14748_4_lut (.I0(n1_adj_4815), .I1(n29773), .I2(n31143), 
            .I3(control_mode[1]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14748_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_652_Mux_15_i1_3_lut (.I0(encoder0_position[15]), .I1(encoder1_position[15]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4807));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11403_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n11643), 
            .I3(GND_net), .O(n15942));   // verilog/coms.v(127[12] 300[6])
    defparam i11403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14740_4_lut (.I0(n1_adj_4807), .I1(n29773), .I2(n31135), 
            .I3(control_mode[1]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14740_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11404_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n11643), 
            .I3(GND_net), .O(n15943));   // verilog/coms.v(127[12] 300[6])
    defparam i11404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11405_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n11643), 
            .I3(GND_net), .O(n15944));   // verilog/coms.v(127[12] 300[6])
    defparam i11405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11244_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n4725), .I3(GND_net), .O(n15783));   // verilog/coms.v(127[12] 300[6])
    defparam i11244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11406_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n11643), 
            .I3(GND_net), .O(n15945));   // verilog/coms.v(127[12] 300[6])
    defparam i11406_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF h1_38 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_LUT4 i11407_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n11643), 
            .I3(GND_net), .O(n15946));   // verilog/coms.v(127[12] 300[6])
    defparam i11407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_24_lut (.I0(duty[22]), .I1(n31935), .I2(n3), .I3(n23506), 
            .O(pwm_setpoint_22__N_3[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i25548_2_lut (.I0(displacement[16]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31134));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25548_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_16_i1_3_lut (.I0(encoder0_position[16]), .I1(encoder1_position[16]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4806));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_16_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_IO SCL_pad (.PACKAGE_PIN(SCL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCL_pad.PIN_TYPE = 6'b011001;
    defparam SCL_pad.PULLUP = 1'b0;
    defparam SCL_pad.NEG_TRIGGER = 1'b0;
    defparam SCL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i11408_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n11643), 
            .I3(GND_net), .O(n15947));   // verilog/coms.v(127[12] 300[6])
    defparam i11408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14739_4_lut (.I0(n1_adj_4806), .I1(n29773), .I2(n31134), 
            .I3(control_mode[1]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14739_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11409_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n11643), 
            .I3(GND_net), .O(n15948));   // verilog/coms.v(127[12] 300[6])
    defparam i11409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11410_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n11643), 
            .I3(GND_net), .O(n15949));   // verilog/coms.v(127[12] 300[6])
    defparam i11410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25547_2_lut (.I0(displacement[17]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31133));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25547_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_17_i1_3_lut (.I0(encoder0_position[17]), .I1(encoder1_position[17]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4805));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14738_4_lut (.I0(n1_adj_4805), .I1(n29773), .I2(n31133), 
            .I3(control_mode[1]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14738_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i25546_2_lut (.I0(displacement[18]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31132));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25546_2_lut.LUT_INIT = 16'h2222;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_534_23_lut (.I0(duty[21]), .I1(n31935), .I2(n4), .I3(n23505), 
            .O(pwm_setpoint_22__N_3[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4758));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11411_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n11643), 
            .I3(GND_net), .O(n15950));   // verilog/coms.v(127[12] 300[6])
    defparam i11411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11412_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n11643), 
            .I3(GND_net), .O(n15951));   // verilog/coms.v(127[12] 300[6])
    defparam i11412_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_534_23 (.CI(n23505), .I0(n31935), .I1(n4), .CO(n23506));
    SB_LUT4 i11413_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n11643), 
            .I3(GND_net), .O(n15952));   // verilog/coms.v(127[12] 300[6])
    defparam i11413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11414_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n11643), .I3(GND_net), .O(n15953));   // verilog/coms.v(127[12] 300[6])
    defparam i11414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11415_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n11643), .I3(GND_net), .O(n15954));   // verilog/coms.v(127[12] 300[6])
    defparam i11415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11416_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n11643), .I3(GND_net), .O(n15955));   // verilog/coms.v(127[12] 300[6])
    defparam i11416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11417_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n11643), .I3(GND_net), .O(n15956));   // verilog/coms.v(127[12] 300[6])
    defparam i11417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11418_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n11643), .I3(GND_net), .O(n15957));   // verilog/coms.v(127[12] 300[6])
    defparam i11418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11419_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n11643), .I3(GND_net), .O(n15958));   // verilog/coms.v(127[12] 300[6])
    defparam i11419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_Mux_18_i1_3_lut (.I0(encoder0_position[18]), .I1(encoder1_position[18]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4804));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_18_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14737_4_lut (.I0(n1_adj_4804), .I1(n29773), .I2(n31132), 
            .I3(control_mode[1]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14737_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i25545_2_lut (.I0(displacement[19]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31131));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25545_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_19_i1_3_lut (.I0(encoder0_position[19]), .I1(encoder1_position[19]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4803));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_19_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14736_4_lut (.I0(n1_adj_4803), .I1(n29773), .I2(n31131), 
            .I3(control_mode[1]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14736_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11420_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n11643), .I3(GND_net), .O(n15959));   // verilog/coms.v(127[12] 300[6])
    defparam i11420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25544_2_lut (.I0(displacement[20]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31130));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25544_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11421_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n11643), .I3(GND_net), .O(n15960));   // verilog/coms.v(127[12] 300[6])
    defparam i11421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11422_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n11643), .I3(GND_net), .O(n15961));   // verilog/coms.v(127[12] 300[6])
    defparam i11422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_Mux_20_i1_3_lut (.I0(encoder0_position[20]), .I1(encoder1_position[20]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4802));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_20_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14735_4_lut (.I0(n1_adj_4802), .I1(n29773), .I2(n31130), 
            .I3(control_mode[1]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14735_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11423_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n11643), .I3(GND_net), .O(n15962));   // verilog/coms.v(127[12] 300[6])
    defparam i11423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11424_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n11643), .I3(GND_net), .O(n15963));   // verilog/coms.v(127[12] 300[6])
    defparam i11424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11425_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n11643), .I3(GND_net), .O(n15964));   // verilog/coms.v(127[12] 300[6])
    defparam i11425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25543_2_lut (.I0(displacement[21]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31129));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25543_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_21_i1_3_lut (.I0(encoder0_position[21]), .I1(encoder1_position[21]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4801));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14734_4_lut (.I0(n1_adj_4801), .I1(n29773), .I2(n31129), 
            .I3(control_mode[1]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14734_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11426_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n11643), .I3(GND_net), .O(n15965));   // verilog/coms.v(127[12] 300[6])
    defparam i11426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25542_2_lut (.I0(displacement[22]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31128));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25542_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11427_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n11643), .I3(GND_net), .O(n15966));   // verilog/coms.v(127[12] 300[6])
    defparam i11427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11428_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n11643), .I3(GND_net), .O(n15967));   // verilog/coms.v(127[12] 300[6])
    defparam i11428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_Mux_22_i1_3_lut (.I0(encoder0_position[22]), .I1(encoder1_position[22]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4800));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14733_4_lut (.I0(n1_adj_4800), .I1(n29773), .I2(n31128), 
            .I3(control_mode[1]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14733_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11429_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n11643), .I3(GND_net), .O(n15968));   // verilog/coms.v(127[12] 300[6])
    defparam i11429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11430_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n11643), .I3(GND_net), .O(n15969));   // verilog/coms.v(127[12] 300[6])
    defparam i11430_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[0]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_LUT4 i11431_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n11643), .I3(GND_net), .O(n15970));   // verilog/coms.v(127[12] 300[6])
    defparam i11431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11432_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n11643), .I3(GND_net), .O(n15971));   // verilog/coms.v(127[12] 300[6])
    defparam i11432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11433_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n11643), .I3(GND_net), .O(n15972));   // verilog/coms.v(127[12] 300[6])
    defparam i11433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11434_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n11643), .I3(GND_net), .O(n15973));   // verilog/coms.v(127[12] 300[6])
    defparam i11434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11435_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n11643), .I3(GND_net), .O(n15974));   // verilog/coms.v(127[12] 300[6])
    defparam i11435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11436_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n11643), .I3(GND_net), .O(n15975));   // verilog/coms.v(127[12] 300[6])
    defparam i11436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11437_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n11643), .I3(GND_net), .O(n15976));   // verilog/coms.v(127[12] 300[6])
    defparam i11437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11438_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n11643), .I3(GND_net), .O(n15977));   // verilog/coms.v(127[12] 300[6])
    defparam i11438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11439_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n11643), .I3(GND_net), .O(n15978));   // verilog/coms.v(127[12] 300[6])
    defparam i11439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11440_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n11643), .I3(GND_net), .O(n15979));   // verilog/coms.v(127[12] 300[6])
    defparam i11440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11441_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n11643), .I3(GND_net), .O(n15980));   // verilog/coms.v(127[12] 300[6])
    defparam i11441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_22_lut (.I0(duty[20]), .I1(n31935), .I2(n5_adj_4758), 
            .I3(n23504), .O(pwm_setpoint_22__N_3[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_22 (.CI(n23504), .I0(n31935), .I1(n5_adj_4758), .CO(n23505));
    SB_LUT4 i11442_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n11643), .I3(GND_net), .O(n15981));   // verilog/coms.v(127[12] 300[6])
    defparam i11442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11443_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n11643), .I3(GND_net), .O(n15982));   // verilog/coms.v(127[12] 300[6])
    defparam i11443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11444_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n11643), .I3(GND_net), .O(n15983));   // verilog/coms.v(127[12] 300[6])
    defparam i11444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11445_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n11643), .I3(GND_net), .O(n15984));   // verilog/coms.v(127[12] 300[6])
    defparam i11445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25556_2_lut (.I0(displacement[8]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31142));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25556_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_534_21_lut (.I0(duty[19]), .I1(n31935), .I2(n6), .I3(n23503), 
            .O(pwm_setpoint_22__N_3[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_21 (.CI(n23503), .I0(n31935), .I1(n6), .CO(n23504));
    SB_LUT4 add_534_20_lut (.I0(duty[18]), .I1(n31935), .I2(n7), .I3(n23502), 
            .O(pwm_setpoint_22__N_3[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i4_4_lut (.I0(control_mode[5]), .I1(control_mode[7]), .I2(control_mode[4]), 
            .I3(control_mode[6]), .O(n10_adj_4761));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[3]), .I1(n10_adj_4761), .I2(control_mode[2]), 
            .I3(GND_net), .O(n29773));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i25537_2_lut (.I0(displacement[23]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31127));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25537_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_23_i1_3_lut (.I0(encoder0_position[23]), .I1(encoder1_position[23]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4799));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_23_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14732_4_lut (.I0(n1_adj_4799), .I1(n29773), .I2(n31127), 
            .I3(control_mode[1]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14732_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_534_20 (.CI(n23502), .I0(n31935), .I1(n7), .CO(n23503));
    SB_LUT4 i11446_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n11643), .I3(GND_net), .O(n15985));   // verilog/coms.v(127[12] 300[6])
    defparam i11446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11447_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n11643), .I3(GND_net), .O(n15986));   // verilog/coms.v(127[12] 300[6])
    defparam i11447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11448_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n11643), .I3(GND_net), .O(n15987));   // verilog/coms.v(127[12] 300[6])
    defparam i11448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_Mux_8_i1_3_lut (.I0(encoder0_position[8]), .I1(encoder1_position[8]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4814));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_8_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11449_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n11643), .I3(GND_net), .O(n15988));   // verilog/coms.v(127[12] 300[6])
    defparam i11449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11450_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n11643), .I3(GND_net), .O(n15989));   // verilog/coms.v(127[12] 300[6])
    defparam i11450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11451_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n11643), .I3(GND_net), .O(n15990));   // verilog/coms.v(127[12] 300[6])
    defparam i11451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11452_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n11643), .I3(GND_net), .O(n15991));   // verilog/coms.v(127[12] 300[6])
    defparam i11452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11453_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n11643), .I3(GND_net), .O(n15992));   // verilog/coms.v(127[12] 300[6])
    defparam i11453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11454_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n11643), .I3(GND_net), .O(n15993));   // verilog/coms.v(127[12] 300[6])
    defparam i11454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11455_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n11643), .I3(GND_net), .O(n15994));   // verilog/coms.v(127[12] 300[6])
    defparam i11455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11456_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n11643), .I3(GND_net), .O(n15995));   // verilog/coms.v(127[12] 300[6])
    defparam i11456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_19_lut (.I0(duty[17]), .I1(n31935), .I2(n8), .I3(n23501), 
            .O(pwm_setpoint_22__N_3[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14747_4_lut (.I0(n1_adj_4814), .I1(n29773), .I2(n31142), 
            .I3(control_mode[1]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14747_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_534_19 (.CI(n23501), .I0(n31935), .I1(n8), .CO(n23502));
    SB_LUT4 add_534_18_lut (.I0(duty[16]), .I1(n31935), .I2(n9), .I3(n23500), 
            .O(pwm_setpoint_22__N_3[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11457_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n11643), .I3(GND_net), .O(n15996));   // verilog/coms.v(127[12] 300[6])
    defparam i11457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11458_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n11643), .I3(GND_net), .O(n15997));   // verilog/coms.v(127[12] 300[6])
    defparam i11458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11459_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n11643), .I3(GND_net), .O(n15998));   // verilog/coms.v(127[12] 300[6])
    defparam i11459_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_534_18 (.CI(n23500), .I0(n31935), .I1(n9), .CO(n23501));
    SB_LUT4 add_534_17_lut (.I0(duty[15]), .I1(n31935), .I2(n10), .I3(n23499), 
            .O(pwm_setpoint_22__N_3[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_17 (.CI(n23499), .I0(n31935), .I1(n10), .CO(n23500));
    SB_LUT4 add_534_16_lut (.I0(duty[14]), .I1(n31935), .I2(n11), .I3(n23498), 
            .O(pwm_setpoint_22__N_3[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11460_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n11643), .I3(GND_net), .O(n15999));   // verilog/coms.v(127[12] 300[6])
    defparam i11460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11461_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n11643), .I3(GND_net), .O(n16000));   // verilog/coms.v(127[12] 300[6])
    defparam i11461_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_534_16 (.CI(n23498), .I0(n31935), .I1(n11), .CO(n23499));
    SB_LUT4 add_534_15_lut (.I0(duty[13]), .I1(n31935), .I2(n12), .I3(n23497), 
            .O(pwm_setpoint_22__N_3[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_15 (.CI(n23497), .I0(n31935), .I1(n12), .CO(n23498));
    SB_LUT4 i11462_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n4727), .I3(GND_net), .O(n16001));   // verilog/coms.v(127[12] 300[6])
    defparam i11462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11463_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n4727), .I3(GND_net), .O(n16002));   // verilog/coms.v(127[12] 300[6])
    defparam i11463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11464_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n4727), .I3(GND_net), .O(n16003));   // verilog/coms.v(127[12] 300[6])
    defparam i11464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11465_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n4727), .I3(GND_net), .O(n16004));   // verilog/coms.v(127[12] 300[6])
    defparam i11465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11466_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n4727), .I3(GND_net), .O(n16005));   // verilog/coms.v(127[12] 300[6])
    defparam i11466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11467_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n4727), .I3(GND_net), .O(n16006));   // verilog/coms.v(127[12] 300[6])
    defparam i11467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11468_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n4727), .I3(GND_net), .O(n16007));   // verilog/coms.v(127[12] 300[6])
    defparam i11468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_14_lut (.I0(duty[12]), .I1(n31935), .I2(n13), .I3(n23496), 
            .O(pwm_setpoint_22__N_3[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11469_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n4727), .I3(GND_net), .O(n16008));   // verilog/coms.v(127[12] 300[6])
    defparam i11469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11470_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n4727), .I3(GND_net), .O(n16009));   // verilog/coms.v(127[12] 300[6])
    defparam i11470_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_534_14 (.CI(n23496), .I0(n31935), .I1(n13), .CO(n23497));
    SB_LUT4 add_534_13_lut (.I0(duty[11]), .I1(n31935), .I2(n14), .I3(n23495), 
            .O(pwm_setpoint_22__N_3[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11471_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n4727), .I3(GND_net), .O(n16010));   // verilog/coms.v(127[12] 300[6])
    defparam i11471_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_534_13 (.CI(n23495), .I0(n31935), .I1(n14), .CO(n23496));
    SB_LUT4 add_534_12_lut (.I0(duty[10]), .I1(n31935), .I2(n15), .I3(n23494), 
            .O(pwm_setpoint_22__N_3[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11472_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n4727), .I3(GND_net), .O(n16011));   // verilog/coms.v(127[12] 300[6])
    defparam i11472_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_534_12 (.CI(n23494), .I0(n31935), .I1(n15), .CO(n23495));
    SB_LUT4 add_534_11_lut (.I0(duty[9]), .I1(n31935), .I2(n16), .I3(n23493), 
            .O(pwm_setpoint_22__N_3[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11473_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n4727), .I3(GND_net), .O(n16012));   // verilog/coms.v(127[12] 300[6])
    defparam i11473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11474_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n4727), .I3(GND_net), .O(n16013));   // verilog/coms.v(127[12] 300[6])
    defparam i11474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11475_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n4727), .I3(GND_net), .O(n16014));   // verilog/coms.v(127[12] 300[6])
    defparam i11475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_534_11 (.CI(n23493), .I0(n31935), .I1(n16), .CO(n23494));
    SB_LUT4 add_534_10_lut (.I0(duty[8]), .I1(n31935), .I2(n17), .I3(n23492), 
            .O(pwm_setpoint_22__N_3[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_10 (.CI(n23492), .I0(n31935), .I1(n17), .CO(n23493));
    SB_LUT4 i11242_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n4725), .I3(GND_net), .O(n15781));   // verilog/coms.v(127[12] 300[6])
    defparam i11242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11243_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n4725), .I3(GND_net), .O(n15782));   // verilog/coms.v(127[12] 300[6])
    defparam i11243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_9_lut (.I0(duty[7]), .I1(n31935), .I2(n18), .I3(n23491), 
            .O(pwm_setpoint_22__N_3[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_9 (.CI(n23491), .I0(n31935), .I1(n18), .CO(n23492));
    SB_LUT4 i11476_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n4727), .I3(GND_net), .O(n16015));   // verilog/coms.v(127[12] 300[6])
    defparam i11476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_8_lut (.I0(duty[6]), .I1(n31935), .I2(n19), .I3(n23490), 
            .O(pwm_setpoint_22__N_3[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_8 (.CI(n23490), .I0(n31935), .I1(n19), .CO(n23491));
    SB_LUT4 i11477_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n4727), .I3(GND_net), .O(n16016));   // verilog/coms.v(127[12] 300[6])
    defparam i11477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11478_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n4727), .I3(GND_net), .O(n16017));   // verilog/coms.v(127[12] 300[6])
    defparam i11478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11479_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n4727), .I3(GND_net), .O(n16018));   // verilog/coms.v(127[12] 300[6])
    defparam i11479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11230_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n4725), .I3(GND_net), .O(n15769));   // verilog/coms.v(127[12] 300[6])
    defparam i11230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11480_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n4727), .I3(GND_net), .O(n16019));   // verilog/coms.v(127[12] 300[6])
    defparam i11480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11231_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n4725), .I3(GND_net), .O(n15770));   // verilog/coms.v(127[12] 300[6])
    defparam i11231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_7_lut (.I0(duty[5]), .I1(n31935), .I2(n20), .I3(n23489), 
            .O(pwm_setpoint_22__N_3[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_7 (.CI(n23489), .I0(n31935), .I1(n20), .CO(n23490));
    SB_LUT4 i11481_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n4727), .I3(GND_net), .O(n16020));   // verilog/coms.v(127[12] 300[6])
    defparam i11481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11482_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n4727), .I3(GND_net), .O(n16021));   // verilog/coms.v(127[12] 300[6])
    defparam i11482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_534_6_lut (.I0(duty[4]), .I1(n31935), .I2(n21), .I3(n23488), 
            .O(pwm_setpoint_22__N_3[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11483_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n4727), .I3(GND_net), .O(n16022));   // verilog/coms.v(127[12] 300[6])
    defparam i11483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25555_2_lut (.I0(displacement[9]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31141));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25555_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11484_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n4727), .I3(GND_net), .O(n16023));   // verilog/coms.v(127[12] 300[6])
    defparam i11484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11232_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n4725), .I3(GND_net), .O(n15771));   // verilog/coms.v(127[12] 300[6])
    defparam i11232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25403_2_lut (.I0(displacement[0]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31082));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25403_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_0_i1_3_lut (.I0(encoder0_position[0]), .I1(encoder1_position[0]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14595_4_lut (.I0(n1), .I1(n29773), .I2(n31082), .I3(control_mode[1]), 
            .O(motor_state[0]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14595_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11241_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n4725), .I3(GND_net), .O(n15780));   // verilog/coms.v(127[12] 300[6])
    defparam i11241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25563_2_lut (.I0(displacement[1]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31149));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25563_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_1_i1_3_lut (.I0(encoder0_position[1]), .I1(encoder1_position[1]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4821));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_1_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14754_4_lut (.I0(n1_adj_4821), .I1(n29773), .I2(n31149), 
            .I3(control_mode[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14754_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i25562_2_lut (.I0(displacement[2]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31148));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25562_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_2_i1_3_lut (.I0(encoder0_position[2]), .I1(encoder1_position[2]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4820));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_2_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14753_4_lut (.I0(n1_adj_4820), .I1(n29773), .I2(n31148), 
            .I3(control_mode[1]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14753_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_534_6 (.CI(n23488), .I0(n31935), .I1(n21), .CO(n23489));
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(144[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4790));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_26[23]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_26[22]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_26[21]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_26[20]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_26[19]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_26[18]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_26[17]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_26[16]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_26[15]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_26[14]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_26[13]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_26[12]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_26[11]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_26[10]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_26[9]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_26[8]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_26[7]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_26[6]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_26[5]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_26[4]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_26[3]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_26[2]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_26[1]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[22]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[21]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[20]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[19]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[18]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[17]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[16]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[15]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[14]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[13]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[12]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[11]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[10]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[9]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[8]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[7]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[6]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[5]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[4]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[3]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[2]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[1]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_LUT4 add_534_5_lut (.I0(duty[3]), .I1(n31935), .I2(n22), .I3(n23487), 
            .O(pwm_setpoint_22__N_3[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i25561_2_lut (.I0(displacement[3]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31147));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25561_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_534_5 (.CI(n23487), .I0(n31935), .I1(n22), .CO(n23488));
    SB_LUT4 add_534_4_lut (.I0(duty[2]), .I1(n31935), .I2(n23), .I3(n23486), 
            .O(pwm_setpoint_22__N_3[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_652_Mux_3_i1_3_lut (.I0(encoder0_position[3]), .I1(encoder1_position[3]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4819));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_Mux_9_i1_3_lut (.I0(encoder0_position[9]), .I1(encoder1_position[9]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4813));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_9_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14746_4_lut (.I0(n1_adj_4813), .I1(n29773), .I2(n31141), 
            .I3(control_mode[1]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14746_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i14752_4_lut (.I0(n1_adj_4819), .I1(n29773), .I2(n31147), 
            .I3(control_mode[1]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14752_4_lut.LUT_INIT = 16'h3022;
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_534_4 (.CI(n23486), .I0(n31935), .I1(n23), .CO(n23487));
    SB_LUT4 i11233_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n4725), .I3(GND_net), .O(n15772));   // verilog/coms.v(127[12] 300[6])
    defparam i11233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11234_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n4725), .I3(GND_net), .O(n15773));   // verilog/coms.v(127[12] 300[6])
    defparam i11234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11235_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n4725), .I3(GND_net), .O(n15774));   // verilog/coms.v(127[12] 300[6])
    defparam i11235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11236_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n4725), .I3(GND_net), .O(n15775));   // verilog/coms.v(127[12] 300[6])
    defparam i11236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11237_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n4725), .I3(GND_net), .O(n15776));   // verilog/coms.v(127[12] 300[6])
    defparam i11237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11238_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n4725), .I3(GND_net), .O(n15777));   // verilog/coms.v(127[12] 300[6])
    defparam i11238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11239_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n4725), .I3(GND_net), .O(n15778));   // verilog/coms.v(127[12] 300[6])
    defparam i11239_3_lut.LUT_INIT = 16'hcaca;
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i11240_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n4725), .I3(GND_net), .O(n15779));   // verilog/coms.v(127[12] 300[6])
    defparam i11240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25560_2_lut (.I0(displacement[4]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31146));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25560_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_4_i1_3_lut (.I0(encoder0_position[4]), .I1(encoder1_position[4]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4818));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_4_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22820_2_lut_3_lut_4_lut (.I0(n14295), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n771), .O(n28639));
    defparam i22820_2_lut_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i1_4_lut_4_lut (.I0(n14309), .I1(n63), .I2(n771), .I3(n27831), 
            .O(n5_adj_4795));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hcc04;
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n2), .I3(n23722), .O(displacement_23__N_26[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25554_2_lut (.I0(displacement[10]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31140));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25554_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i25552_2_lut (.I0(displacement[12]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31138));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25552_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4790), .I3(n23721), .O(displacement_23__N_26[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n23721), .I0(encoder1_position[22]), 
            .I1(n3_adj_4790), .CO(n23722));
    SB_LUT4 mux_652_Mux_10_i1_3_lut (.I0(encoder0_position[10]), .I1(encoder1_position[10]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4812));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_10_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14745_4_lut (.I0(n1_adj_4812), .I1(n29773), .I2(n31140), 
            .I3(control_mode[1]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14745_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_652_Mux_12_i1_3_lut (.I0(encoder0_position[12]), .I1(encoder1_position[12]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4810));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_12_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n4_adj_4789), .I3(n23720), .O(displacement_23__N_26[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n23720), .I0(encoder1_position[21]), 
            .I1(n4_adj_4789), .CO(n23721));
    SB_LUT4 i14743_4_lut (.I0(n1_adj_4810), .I1(n29773), .I2(n31138), 
            .I3(control_mode[1]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14743_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_534_3_lut (.I0(duty[1]), .I1(n31935), .I2(n24), .I3(n23485), 
            .O(pwm_setpoint_22__N_3[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_3 (.CI(n23485), .I0(n31935), .I1(n24), .CO(n23486));
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5), .I3(n23719), .O(displacement_23__N_26[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n23719), .I0(encoder1_position[20]), 
            .I1(n5), .CO(n23720));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4770));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_534_2_lut (.I0(duty[0]), .I1(n31935), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_3[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_534_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_534_2 (.CI(VCC_net), .I0(n31935), .I1(n25), .CO(n23485));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4764), .I3(n23718), .O(displacement_23__N_26[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n23718), .I0(encoder1_position[19]), 
            .I1(n6_adj_4764), .CO(n23719));
    SB_LUT4 i25553_2_lut (.I0(displacement[11]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31139));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i25553_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_652_Mux_11_i1_3_lut (.I0(encoder0_position[11]), .I1(encoder1_position[11]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4811));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_652_Mux_11_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4765), .I3(n23717), .O(displacement_23__N_26[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n23717), .I0(encoder1_position[18]), 
            .I1(n7_adj_4765), .CO(n23718));
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4766), .I3(n23716), .O(displacement_23__N_26[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n23716), .I0(encoder1_position[17]), 
            .I1(n8_adj_4766), .CO(n23717));
    SB_LUT4 i14744_4_lut (.I0(n1_adj_4811), .I1(n29773), .I2(n31139), 
            .I3(control_mode[1]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14744_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11660_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4725), .I3(GND_net), .O(n16199));   // verilog/coms.v(127[12] 300[6])
    defparam i11660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11664_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4763), 
            .I3(n14282), .O(n16203));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11664_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11665_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4725), .I3(GND_net), .O(n16204));   // verilog/coms.v(127[12] 300[6])
    defparam i11665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11666_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4725), .I3(GND_net), .O(n16205));   // verilog/coms.v(127[12] 300[6])
    defparam i11666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11667_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4725), .I3(GND_net), .O(n16206));   // verilog/coms.v(127[12] 300[6])
    defparam i11667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11668_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4725), .I3(GND_net), .O(n16207));   // verilog/coms.v(127[12] 300[6])
    defparam i11668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11669_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4725), .I3(GND_net), .O(n16208));   // verilog/coms.v(127[12] 300[6])
    defparam i11669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11670_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4725), .I3(GND_net), .O(n16209));   // verilog/coms.v(127[12] 300[6])
    defparam i11670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4767), .I3(n23715), .O(displacement_23__N_26[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n23715), .I0(encoder1_position[16]), 
            .I1(n9_adj_4767), .CO(n23716));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4768), .I3(n23714), .O(displacement_23__N_26[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11671_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n4725), .I3(GND_net), .O(n16210));   // verilog/coms.v(127[12] 300[6])
    defparam i11671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11672_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n4725), .I3(GND_net), .O(n16211));   // verilog/coms.v(127[12] 300[6])
    defparam i11672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11673_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n4725), .I3(GND_net), .O(n16212));   // verilog/coms.v(127[12] 300[6])
    defparam i11673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3422[2]), 
            .I3(r_SM_Main[0]), .O(n15488));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n15488), 
            .I3(rx_data_ready), .O(n27405));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i26069_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n27820));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i26069_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n23714), .I0(encoder1_position[15]), 
            .I1(n10_adj_4768), .CO(n23715));
    SB_LUT4 i11674_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n4725), .I3(GND_net), .O(n16213));   // verilog/coms.v(127[12] 300[6])
    defparam i11674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4769), .I3(n23713), .O(displacement_23__N_26[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11675_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n4725), .I3(GND_net), .O(n16214));   // verilog/coms.v(127[12] 300[6])
    defparam i11675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11676_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n4725), .I3(GND_net), .O(n16215));   // verilog/coms.v(127[12] 300[6])
    defparam i11676_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_26[0]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n23713), .I0(encoder1_position[14]), 
            .I1(n11_adj_4769), .CO(n23714));
    SB_LUT4 i11677_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n4725), .I3(GND_net), .O(n16216));   // verilog/coms.v(127[12] 300[6])
    defparam i11677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4770), .I3(n23712), .O(displacement_23__N_26[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11678_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n4725), .I3(GND_net), .O(n16217));   // verilog/coms.v(127[12] 300[6])
    defparam i11678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11679_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n4725), .I3(GND_net), .O(n16218));   // verilog/coms.v(127[12] 300[6])
    defparam i11679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11680_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n4725), .I3(GND_net), .O(n16219));   // verilog/coms.v(127[12] 300[6])
    defparam i11680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11681_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n4725), .I3(GND_net), .O(n16220));   // verilog/coms.v(127[12] 300[6])
    defparam i11681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4769));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11682_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n4725), .I3(GND_net), .O(n16221));   // verilog/coms.v(127[12] 300[6])
    defparam i11682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11683_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n4725), .I3(GND_net), .O(n16222));   // verilog/coms.v(127[12] 300[6])
    defparam i11683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11684_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n4725), .I3(GND_net), .O(n16223));   // verilog/coms.v(127[12] 300[6])
    defparam i11684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11685_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n4725), .I3(GND_net), .O(n16224));   // verilog/coms.v(127[12] 300[6])
    defparam i11685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11686_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n4725), .I3(GND_net), .O(n16225));   // verilog/coms.v(127[12] 300[6])
    defparam i11686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11687_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n4725), .I3(GND_net), .O(n16226));   // verilog/coms.v(127[12] 300[6])
    defparam i11687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11688_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n4725), .I3(GND_net), .O(n16227));   // verilog/coms.v(127[12] 300[6])
    defparam i11688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11689_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n4725), .I3(GND_net), .O(n16228));   // verilog/coms.v(127[12] 300[6])
    defparam i11689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11690_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n4725), .I3(GND_net), .O(n16229));   // verilog/coms.v(127[12] 300[6])
    defparam i11690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11691_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n4725), .I3(GND_net), .O(n16230));   // verilog/coms.v(127[12] 300[6])
    defparam i11691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11692_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n4725), .I3(GND_net), .O(n16231));   // verilog/coms.v(127[12] 300[6])
    defparam i11692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11693_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n4725), .I3(GND_net), .O(n16232));   // verilog/coms.v(127[12] 300[6])
    defparam i11693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1623 (.I0(n27831), .I1(n14328), .I2(n23_adj_4822), 
            .I3(n4452), .O(n27755));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1623.LUT_INIT = 16'hafbf;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n23712), .I0(encoder1_position[13]), 
            .I1(n12_adj_4770), .CO(n23713));
    SB_LUT4 i1_3_lut (.I0(n123), .I1(n27755), .I2(n63), .I3(GND_net), 
            .O(n7_adj_4759));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut.LUT_INIT = 16'h8c8c;
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4771), .I3(n23711), .O(displacement_23__N_26[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n23711), .I0(encoder1_position[12]), 
            .I1(n13_adj_4771), .CO(n23712));
    SB_LUT4 i2_4_lut_adj_1624 (.I0(n7_adj_4759), .I1(n123), .I2(n14309), 
            .I3(n8515), .O(n6_adj_4823));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1624.LUT_INIT = 16'haeaf;
    SB_LUT4 i3_4_lut (.I0(n63_adj_4788), .I1(n6_adj_4823), .I2(n14318), 
            .I3(\FRAME_MATCHER.state_31__N_2668 [1]), .O(n32532));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hdfdd;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_4867[1]), .I1(r_SM_Main_adj_4867[0]), 
            .I2(r_SM_Main_adj_4867[2]), .I3(r_SM_Main_2__N_3493[1]), .O(n32553));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4772), .I3(n23710), .O(displacement_23__N_26[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1625 (.I0(n5_adj_4798), .I1(n122), .I2(n23_adj_4822), 
            .I3(n63), .O(n6_adj_4760));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'haeaa;
    SB_LUT4 i3_4_lut_adj_1626 (.I0(n32898), .I1(n6_adj_4760), .I2(n14328), 
            .I3(n4452), .O(n8_adj_4824));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1626.LUT_INIT = 16'hcfce;
    SB_LUT4 i4_4_lut_adj_1627 (.I0(n122), .I1(n8_adj_4824), .I2(n63_adj_4788), 
            .I3(n5_adj_4795), .O(n32531));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1627.LUT_INIT = 16'hefcf;
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n23710), .I0(encoder1_position[11]), 
            .I1(n14_adj_4772), .CO(n23711));
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4773), .I3(n23709), .O(displacement_23__N_26[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25565_3_lut (.I0(start), .I1(n28731), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n31069));   // verilog/neopixel.v(35[12] 117[6])
    defparam i25565_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i18_4_lut (.I0(n31069), .I1(n29426), .I2(state[1]), .I3(start), 
            .O(n26505));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i11698_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n30174), 
            .I3(GND_net), .O(n16237));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11698_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11225_3_lut (.I0(n15643), .I1(r_Bit_Index[0]), .I2(n15548), 
            .I3(GND_net), .O(n15764));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11225_3_lut.LUT_INIT = 16'h1414;
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n23709), .I0(encoder1_position[10]), 
            .I1(n15_adj_4773), .CO(n23710));
    SB_LUT4 i11700_3_lut (.I0(quadA_debounced_adj_4785), .I1(reg_B_adj_4879[1]), 
            .I2(n29458), .I3(GND_net), .O(n16239));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11700_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11191_3_lut (.I0(n28775), .I1(r_Bit_Index_adj_4869[0]), .I2(n28749), 
            .I3(GND_net), .O(n15730));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11191_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i11702_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1138), .I3(GND_net), .O(n16241));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11703_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1138), .I3(GND_net), .O(n16242));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11704_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1138), .I3(GND_net), .O(n16243));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11705_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1138), .I3(GND_net), .O(n16244));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11706_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1138), .I3(GND_net), .O(n16245));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11707_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1138), .I3(GND_net), .O(n16246));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11708_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1138), .I3(GND_net), .O(n16247));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4774), .I3(n23708), .O(displacement_23__N_26[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n23708), .I0(encoder1_position[9]), 
            .I1(n16_adj_4774), .CO(n23709));
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    GND i1 (.Y(GND_net));
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced_adj_4785, 
            quadB_debounced_adj_4786}), .reg_B({reg_B_adj_4879}), .n29458(n29458), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n16239(n16239), .n15723(n15723)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(195[15] 200[4])
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4775), .I3(n23707), .O(displacement_23__N_26[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n23707), .I0(encoder1_position[8]), 
            .I1(n17_adj_4775), .CO(n23708));
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4776), .I3(n23706), .O(displacement_23__N_26[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n23706), .I0(encoder1_position[7]), 
            .I1(n18_adj_4776), .CO(n23707));
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4777), .I3(n23705), .O(displacement_23__N_26[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n23705), .I0(encoder1_position[6]), 
            .I1(n19_adj_4777), .CO(n23706));
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4778), .I3(n23704), .O(displacement_23__N_26[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n23704), .I0(encoder1_position[5]), 
            .I1(n20_adj_4778), .CO(n23705));
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4779), .I3(n23703), .O(displacement_23__N_26[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n23703), .I0(encoder1_position[4]), 
            .I1(n21_adj_4779), .CO(n23704));
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4780), .I3(n23702), .O(displacement_23__N_26[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n23702), .I0(encoder1_position[3]), 
            .I1(n22_adj_4780), .CO(n23703));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4781), .I3(n23701), .O(displacement_23__N_26[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n23701), .I0(encoder1_position[2]), 
            .I1(n23_adj_4781), .CO(n23702));
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4782), .I3(n23700), .O(displacement_23__N_26[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n23700), .I0(encoder1_position[1]), 
            .I1(n24_adj_4782), .CO(n23701));
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4783), .I3(VCC_net), .O(displacement_23__N_26[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4783), .CO(n23700));
    motorControl control (.setpoint({setpoint}), .GND_net(GND_net), .\Kp[12] (Kp[12]), 
            .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[13] (Ki[13]), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
            .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), 
            .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .motor_state({motor_state}), 
            .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .VCC_net(VCC_net), .\Ki[11] (Ki[11]), 
            .\Ki[12] (Ki[12]), .PWMLimit({PWMLimit}), .IntegralLimit({IntegralLimit}), 
            .duty({duty}), .clk32MHz(clk32MHz), .n25(n25), .n31935(n31935)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(172[16] 184[4])
    SB_LUT4 i11245_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n4725), .I3(GND_net), .O(n15784));   // verilog/coms.v(127[12] 300[6])
    defparam i11245_3_lut.LUT_INIT = 16'hcaca;
    coms neopxl_color_23__I_0 (.\data_out_frame[11] ({\data_out_frame[11] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .GND_net(GND_net), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .rx_data({rx_data}), 
         .rx_data_ready(rx_data_ready), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .n15783(n15783), .IntegralLimit({IntegralLimit}), .clk32MHz(clk32MHz), 
         .n15782(n15782), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n15781(n15781), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n15780(n15780), .n15779(n15779), .n15778(n15778), .n15777(n15777), 
         .n15776(n15776), .n15775(n15775), .\FRAME_MATCHER.state[1] (\FRAME_MATCHER.state [1]), 
         .n14318(n14318), .n63(n63), .n3303(n3303), .n15774(n15774), 
         .n15773(n15773), .n15772(n15772), .n4452(n4452), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n14295(n14295), .n23(n23_adj_4822), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .\data_in[3][3] (\data_in[3] [3]), 
         .\data_in[0] ({\data_in[0] }), .\data_in[2] ({\data_in[2] }), .\data_in[3][6] (\data_in[3] [6]), 
         .\data_in[3][1] (\data_in[3] [1]), .\data_in[1] ({\data_in[1] }), 
         .\data_in[3][0] (\data_in[3] [0]), .\data_in[3][4] (\data_in[3] [4]), 
         .\data_in[3][2] (\data_in[3] [2]), .\data_in[3][7] (\data_in[3] [7]), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .n771(n771), .n15771(n15771), 
         .n15770(n15770), .n15769(n15769), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .setpoint({setpoint}), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .n11643(n11643), .\data_in_frame[3] ({\data_in_frame[3] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n4727(n4727), .\data_in_frame[13] ({\data_in_frame[13] }), .n15768(n15768), 
         .n15767(n15767), .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .n15766(n15766), .n15765(n15765), 
         .n4725(n4725), .n29573(n29573), .n63_adj_3(n63_adj_4788), .n14309(n14309), 
         .n123(n123), .DE_c(DE_c), .LED_c(LED_c), .n14328(n14328), .n32531(n32531), 
         .n32532(n32532), .n16232(n16232), .PWMLimit({PWMLimit}), .n16231(n16231), 
         .n16230(n16230), .n16229(n16229), .n16228(n16228), .n16227(n16227), 
         .n16226(n16226), .n16225(n16225), .n16224(n16224), .n16223(n16223), 
         .n16222(n16222), .n16221(n16221), .n16220(n16220), .n16219(n16219), 
         .n16218(n16218), .n16217(n16217), .n16216(n16216), .n16215(n16215), 
         .n16214(n16214), .n16213(n16213), .n16212(n16212), .n16211(n16211), 
         .n16210(n16210), .n16209(n16209), .control_mode({control_mode}), 
         .n16208(n16208), .n16207(n16207), .n16206(n16206), .n16205(n16205), 
         .n16204(n16204), .n16199(n16199), .tx_active(tx_active), .n27831(n27831), 
         .n16023(n16023), .neopxl_color({neopxl_color}), .n16022(n16022), 
         .n16021(n16021), .n16020(n16020), .n16019(n16019), .n16018(n16018), 
         .n16017(n16017), .n16016(n16016), .n16015(n16015), .n16014(n16014), 
         .n16013(n16013), .n16012(n16012), .n16011(n16011), .n16010(n16010), 
         .n16009(n16009), .n16008(n16008), .n16007(n16007), .n16006(n16006), 
         .n16005(n16005), .n16004(n16004), .n16003(n16003), .n16002(n16002), 
         .n16001(n16001), .n16000(n16000), .n15999(n15999), .n15998(n15998), 
         .n15997(n15997), .n15996(n15996), .n15995(n15995), .n15994(n15994), 
         .n15993(n15993), .n15992(n15992), .n15991(n15991), .n15990(n15990), 
         .n15989(n15989), .n15988(n15988), .n15987(n15987), .n15986(n15986), 
         .n15985(n15985), .n15984(n15984), .n15983(n15983), .n15982(n15982), 
         .n15981(n15981), .n15980(n15980), .n15979(n15979), .n15978(n15978), 
         .n15977(n15977), .n15976(n15976), .n15975(n15975), .n15974(n15974), 
         .n15973(n15973), .n15972(n15972), .n15971(n15971), .n15970(n15970), 
         .n15969(n15969), .n15968(n15968), .n15967(n15967), .n15966(n15966), 
         .n15965(n15965), .n15964(n15964), .n15963(n15963), .n15962(n15962), 
         .n15961(n15961), .n15960(n15960), .n15959(n15959), .n15958(n15958), 
         .n15957(n15957), .n15956(n15956), .n15955(n15955), .n15954(n15954), 
         .n15953(n15953), .n15952(n15952), .n15951(n15951), .n15950(n15950), 
         .n15949(n15949), .n15948(n15948), .n15947(n15947), .n15946(n15946), 
         .n15945(n15945), .n15944(n15944), .n15943(n15943), .n15942(n15942), 
         .n15941(n15941), .n15940(n15940), .n15939(n15939), .n15938(n15938), 
         .n15937(n15937), .n15936(n15936), .n15935(n15935), .n15934(n15934), 
         .n15933(n15933), .n15932(n15932), .n15931(n15931), .n15930(n15930), 
         .n15929(n15929), .n15928(n15928), .n15927(n15927), .n15926(n15926), 
         .n15925(n15925), .n15924(n15924), .n15923(n15923), .n15922(n15922), 
         .n15921(n15921), .n15920(n15920), .n15919(n15919), .n15918(n15918), 
         .n15917(n15917), .n15916(n15916), .n15915(n15915), .n15914(n15914), 
         .n15913(n15913), .n15912(n15912), .n15911(n15911), .n15910(n15910), 
         .n15909(n15909), .n15908(n15908), .n15907(n15907), .n15906(n15906), 
         .n15905(n15905), .n15904(n15904), .n15903(n15903), .n15902(n15902), 
         .n15901(n15901), .\FRAME_MATCHER.state_31__N_2668[1] (\FRAME_MATCHER.state_31__N_2668 [1]), 
         .n15900(n15900), .n15899(n15899), .n15898(n15898), .n15897(n15897), 
         .n15896(n15896), .n15895(n15895), .n8515(n8515), .n122(n122), 
         .n5(n5_adj_4798), .n32898(n32898), .n30290(n30290), .n27243(n27243), 
         .n15719(n15719), .n15894(n15894), .n15893(n15893), .n15892(n15892), 
         .n15891(n15891), .n15890(n15890), .n15889(n15889), .n15888(n15888), 
         .n15887(n15887), .n15886(n15886), .n15885(n15885), .n15884(n15884), 
         .n15883(n15883), .n15882(n15882), .n15881(n15881), .n15880(n15880), 
         .n15879(n15879), .n15878(n15878), .n15877(n15877), .n15876(n15876), 
         .n15875(n15875), .n15874(n15874), .n15873(n15873), .n15872(n15872), 
         .n15871(n15871), .n15870(n15870), .n15869(n15869), .n15868(n15868), 
         .n15867(n15867), .n15866(n15866), .n15865(n15865), .n15864(n15864), 
         .n15863(n15863), .n15862(n15862), .n15718(n15718), .n15716(n15716), 
         .n15715(n15715), .\Ki[0] (Ki[0]), .n15714(n15714), .\Kp[0] (Kp[0]), 
         .n15713(n15713), .n15861(n15861), .n15860(n15860), .n15859(n15859), 
         .n15858(n15858), .n15857(n15857), .n15856(n15856), .n15855(n15855), 
         .n15705(n15705), .n15854(n15854), .n15853(n15853), .n15852(n15852), 
         .n15851(n15851), .n15850(n15850), .n15849(n15849), .n15848(n15848), 
         .\Ki[15] (Ki[15]), .n15847(n15847), .\Ki[14] (Ki[14]), .n15846(n15846), 
         .\Ki[13] (Ki[13]), .n15845(n15845), .\Ki[12] (Ki[12]), .n15844(n15844), 
         .\Ki[11] (Ki[11]), .n15843(n15843), .\Ki[10] (Ki[10]), .n15842(n15842), 
         .\Ki[9] (Ki[9]), .n15841(n15841), .\Ki[8] (Ki[8]), .n15840(n15840), 
         .\Ki[7] (Ki[7]), .n15839(n15839), .\Ki[6] (Ki[6]), .n15838(n15838), 
         .\Ki[5] (Ki[5]), .n15837(n15837), .\Ki[4] (Ki[4]), .n15836(n15836), 
         .\Ki[3] (Ki[3]), .n15835(n15835), .\Ki[2] (Ki[2]), .n15834(n15834), 
         .\Ki[1] (Ki[1]), .n15833(n15833), .\Kp[15] (Kp[15]), .n15832(n15832), 
         .\Kp[14] (Kp[14]), .n15831(n15831), .\Kp[13] (Kp[13]), .n15830(n15830), 
         .\Kp[12] (Kp[12]), .n15829(n15829), .\Kp[11] (Kp[11]), .n15828(n15828), 
         .\Kp[10] (Kp[10]), .n15827(n15827), .\Kp[9] (Kp[9]), .n15826(n15826), 
         .\Kp[8] (Kp[8]), .n15825(n15825), .\Kp[7] (Kp[7]), .n15824(n15824), 
         .\Kp[6] (Kp[6]), .n15823(n15823), .\Kp[5] (Kp[5]), .n15822(n15822), 
         .\Kp[4] (Kp[4]), .n15821(n15821), .\Kp[3] (Kp[3]), .n15820(n15820), 
         .\Kp[2] (Kp[2]), .n15819(n15819), .\Kp[1] (Kp[1]), .n15818(n15818), 
         .n15817(n15817), .n15815(n15815), .n15814(n15814), .n15813(n15813), 
         .n15812(n15812), .n15811(n15811), .n15810(n15810), .n15809(n15809), 
         .n15807(n15807), .n15806(n15806), .n15805(n15805), .n15804(n15804), 
         .n15803(n15803), .n15802(n15802), .n15801(n15801), .n15800(n15800), 
         .n15799(n15799), .n15798(n15798), .n15797(n15797), .n15796(n15796), 
         .n15795(n15795), .n15794(n15794), .n15793(n15793), .n15792(n15792), 
         .n15791(n15791), .n15790(n15790), .n15789(n15789), .n15788(n15788), 
         .n15787(n15787), .n15786(n15786), .n15785(n15785), .n15784(n15784), 
         .n28749(n28749), .n28775(n28775), .VCC_net(VCC_net), .r_SM_Main({r_SM_Main_adj_4867}), 
         .n8353(n8353), .tx_o(tx_o), .\r_SM_Main_2__N_3493[1] (r_SM_Main_2__N_3493[1]), 
         .\r_Bit_Index[0] (r_Bit_Index_adj_4869[0]), .n4(n4_adj_4762), .n15730(n15730), 
         .n32553(n32553), .n15722(n15722), .tx_enable(tx_enable), .n15548(n15548), 
         .n15643(n15643), .\r_SM_Main_2__N_3422[2] (r_SM_Main_2__N_3422[2]), 
         .r_SM_Main_adj_11({r_SM_Main}), .n27820(n27820), .r_Rx_Data(r_Rx_Data), 
         .n19238(n19238), .n4_adj_7(n4_adj_4784), .n4_adj_8(n4_adj_4787), 
         .\r_Bit_Index[0]_adj_9 (r_Bit_Index[0]), .n14287(n14287), .RX_N_2(RX_N_2), 
         .n14282(n14282), .n4_adj_10(n4_adj_4763), .n27405(n27405), .n15764(n15764), 
         .n16203(n16203), .n15712(n15712), .n15711(n15711), .n15710(n15710), 
         .n15709(n15709), .n15708(n15708), .n15707(n15707), .n15706(n15706)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(138[8] 161[4])
    SB_LUT4 i11246_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n4725), .I3(GND_net), .O(n15785));   // verilog/coms.v(127[12] 300[6])
    defparam i11246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11247_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n4725), .I3(GND_net), .O(n15786));   // verilog/coms.v(127[12] 300[6])
    defparam i11247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11248_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n4725), .I3(GND_net), .O(n15787));   // verilog/coms.v(127[12] 300[6])
    defparam i11248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11249_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15788));   // verilog/coms.v(127[12] 300[6])
    defparam i11249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11250_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15789));   // verilog/coms.v(127[12] 300[6])
    defparam i11250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4768));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11251_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15790));   // verilog/coms.v(127[12] 300[6])
    defparam i11251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11252_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15791));   // verilog/coms.v(127[12] 300[6])
    defparam i11252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11253_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15792));   // verilog/coms.v(127[12] 300[6])
    defparam i11253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4767));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11254_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15793));   // verilog/coms.v(127[12] 300[6])
    defparam i11254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11255_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15794));   // verilog/coms.v(127[12] 300[6])
    defparam i11255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11256_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15795));   // verilog/coms.v(127[12] 300[6])
    defparam i11256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11257_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15796));   // verilog/coms.v(127[12] 300[6])
    defparam i11257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11258_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15797));   // verilog/coms.v(127[12] 300[6])
    defparam i11258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11259_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15798));   // verilog/coms.v(127[12] 300[6])
    defparam i11259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11260_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15799));   // verilog/coms.v(127[12] 300[6])
    defparam i11260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11261_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15800));   // verilog/coms.v(127[12] 300[6])
    defparam i11261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11262_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15801));   // verilog/coms.v(127[12] 300[6])
    defparam i11262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11263_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15802));   // verilog/coms.v(127[12] 300[6])
    defparam i11263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11264_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15803));   // verilog/coms.v(127[12] 300[6])
    defparam i11264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11265_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15804));   // verilog/coms.v(127[12] 300[6])
    defparam i11265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11266_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15805));   // verilog/coms.v(127[12] 300[6])
    defparam i11266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11267_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15806));   // verilog/coms.v(127[12] 300[6])
    defparam i11267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11268_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15807));   // verilog/coms.v(127[12] 300[6])
    defparam i11268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11270_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15809));   // verilog/coms.v(127[12] 300[6])
    defparam i11270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11192_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n26593), .I3(GND_net), .O(n15731));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11271_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15810));   // verilog/coms.v(127[12] 300[6])
    defparam i11271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11272_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15811));   // verilog/coms.v(127[12] 300[6])
    defparam i11272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4783));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11193_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n26593), .I3(GND_net), .O(n15732));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11193_3_lut.LUT_INIT = 16'hacac;
    \pwm(32000000,20000,32000000,23,1)  PWM (.INHA_c_0(INHA_c_0), .CLK_c(CLK_c), 
            .pwm_setpoint({pwm_setpoint}), .GND_net(GND_net), .\half_duty_new[0] (half_duty_new[0]), 
            .n1138(n1138), .VCC_net(VCC_net), .\half_duty[0][0] (\half_duty[0] [0]), 
            .\half_duty[0][1] (\half_duty[0] [1]), .\half_duty[0][2] (\half_duty[0] [2]), 
            .\half_duty[0][3] (\half_duty[0] [3]), .\half_duty[0][4] (\half_duty[0] [4]), 
            .\half_duty[0][5] (\half_duty[0] [5]), .\half_duty[0][6] (\half_duty[0] [6]), 
            .\half_duty[0][7] (\half_duty[0] [7]), .\half_duty_new[1] (half_duty_new[1]), 
            .\half_duty_new[2] (half_duty_new[2]), .\half_duty_new[3] (half_duty_new[3]), 
            .\half_duty_new[4] (half_duty_new[4]), .\half_duty_new[5] (half_duty_new[5]), 
            .\half_duty_new[6] (half_duty_new[6]), .\half_duty_new[7] (half_duty_new[7]), 
            .n16247(n16247), .n16246(n16246), .n16245(n16245), .n16244(n16244), 
            .n16243(n16243), .n16242(n16242), .n16241(n16241), .n15724(n15724));   // verilog/TinyFPGA_B.v(90[43] 96[3])
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4782));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11273_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15812));   // verilog/coms.v(127[12] 300[6])
    defparam i11273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11274_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15813));   // verilog/coms.v(127[12] 300[6])
    defparam i11274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11194_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n26593), .I3(GND_net), .O(n15733));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11275_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15814));   // verilog/coms.v(127[12] 300[6])
    defparam i11275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11276_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15815));   // verilog/coms.v(127[12] 300[6])
    defparam i11276_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, GND_net, clk32MHz, 
            data_o, reg_B, n30174, ENCODER0_B_c_0, n16237, ENCODER0_A_c_1, 
            n15721) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output [1:0]reg_B;
    output n30174;
    input ENCODER0_B_c_0;
    input n16237;
    input ENCODER0_A_c_1;
    input n15721;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2849;
    
    wire count_direction, n23550, n23551, n2845, count_enable, B_delayed, 
        A_delayed, n23573, n23572, n23571, n23570, n23569, n23568, 
        n23567, n23566, n23565, n23564, n23563, n23562, n23561, 
        n23560, n23559, n23558, n23557, n23556, n23555, n23554, 
        n23553, n23552;
    
    SB_LUT4 add_603_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n23550), .O(n2849[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_2 (.CI(n23550), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n23551));
    SB_CARRY add_603_1 (.CI(GND_net), .I0(n2845), .I1(n2845), .CO(n23550));
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_603_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2845), 
            .I3(n23573), .O(n2849[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_603_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2845), 
            .I3(n23572), .O(n2849[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_24 (.CI(n23572), .I0(encoder0_position[22]), .I1(n2845), 
            .CO(n23573));
    SB_LUT4 add_603_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2845), 
            .I3(n23571), .O(n2849[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i898_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2845));   // quad.v(37[5] 40[8])
    defparam i898_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2849[23]));   // quad.v(35[10] 41[6])
    SB_CARRY add_603_23 (.CI(n23571), .I0(encoder0_position[21]), .I1(n2845), 
            .CO(n23572));
    SB_LUT4 add_603_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2845), 
            .I3(n23570), .O(n2849[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_22 (.CI(n23570), .I0(encoder0_position[20]), .I1(n2845), 
            .CO(n23571));
    SB_LUT4 add_603_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2845), 
            .I3(n23569), .O(n2849[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_21 (.CI(n23569), .I0(encoder0_position[19]), .I1(n2845), 
            .CO(n23570));
    SB_LUT4 add_603_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2845), 
            .I3(n23568), .O(n2849[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_20 (.CI(n23568), .I0(encoder0_position[18]), .I1(n2845), 
            .CO(n23569));
    SB_LUT4 add_603_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2845), 
            .I3(n23567), .O(n2849[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_19 (.CI(n23567), .I0(encoder0_position[17]), .I1(n2845), 
            .CO(n23568));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_603_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2845), 
            .I3(n23566), .O(n2849[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_18 (.CI(n23566), .I0(encoder0_position[16]), .I1(n2845), 
            .CO(n23567));
    SB_LUT4 add_603_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2845), 
            .I3(n23565), .O(n2849[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_17 (.CI(n23565), .I0(encoder0_position[15]), .I1(n2845), 
            .CO(n23566));
    SB_LUT4 add_603_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2845), 
            .I3(n23564), .O(n2849[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_16 (.CI(n23564), .I0(encoder0_position[14]), .I1(n2845), 
            .CO(n23565));
    SB_LUT4 add_603_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2845), 
            .I3(n23563), .O(n2849[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_15 (.CI(n23563), .I0(encoder0_position[13]), .I1(n2845), 
            .CO(n23564));
    SB_LUT4 add_603_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2845), 
            .I3(n23562), .O(n2849[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_14 (.CI(n23562), .I0(encoder0_position[12]), .I1(n2845), 
            .CO(n23563));
    SB_LUT4 add_603_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2845), 
            .I3(n23561), .O(n2849[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_13 (.CI(n23561), .I0(encoder0_position[11]), .I1(n2845), 
            .CO(n23562));
    SB_LUT4 add_603_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2845), 
            .I3(n23560), .O(n2849[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_12 (.CI(n23560), .I0(encoder0_position[10]), .I1(n2845), 
            .CO(n23561));
    SB_LUT4 add_603_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2845), 
            .I3(n23559), .O(n2849[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_11 (.CI(n23559), .I0(encoder0_position[9]), .I1(n2845), 
            .CO(n23560));
    SB_LUT4 add_603_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2845), 
            .I3(n23558), .O(n2849[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_10 (.CI(n23558), .I0(encoder0_position[8]), .I1(n2845), 
            .CO(n23559));
    SB_LUT4 add_603_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2845), 
            .I3(n23557), .O(n2849[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_9 (.CI(n23557), .I0(encoder0_position[7]), .I1(n2845), 
            .CO(n23558));
    SB_LUT4 add_603_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2845), 
            .I3(n23556), .O(n2849[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_8 (.CI(n23556), .I0(encoder0_position[6]), .I1(n2845), 
            .CO(n23557));
    SB_LUT4 add_603_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2845), 
            .I3(n23555), .O(n2849[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_7 (.CI(n23555), .I0(encoder0_position[5]), .I1(n2845), 
            .CO(n23556));
    SB_LUT4 add_603_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2845), 
            .I3(n23554), .O(n2849[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_6 (.CI(n23554), .I0(encoder0_position[4]), .I1(n2845), 
            .CO(n23555));
    SB_LUT4 add_603_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2845), 
            .I3(n23553), .O(n2849[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_5 (.CI(n23553), .I0(encoder0_position[3]), .I1(n2845), 
            .CO(n23554));
    SB_LUT4 add_603_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2845), 
            .I3(n23552), .O(n2849[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_4 (.CI(n23552), .I0(encoder0_position[2]), .I1(n2845), 
            .CO(n23553));
    SB_LUT4 add_603_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2845), 
            .I3(n23551), .O(n2849[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_603_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_603_3 (.CI(n23551), .I0(encoder0_position[1]), .I1(n2845), 
            .CO(n23552));
    \grp_debouncer(2,5)_U0  debounce (.reg_B({reg_B}), .GND_net(GND_net), 
            .n30174(n30174), .clk32MHz(clk32MHz), .ENCODER0_B_c_0(ENCODER0_B_c_0), 
            .n16237(n16237), .data_o({data_o}), .ENCODER0_A_c_1(ENCODER0_A_c_1), 
            .n15721(n15721));   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (reg_B, GND_net, n30174, clk32MHz, ENCODER0_B_c_0, 
            n16237, data_o, ENCODER0_A_c_1, n15721);
    output [1:0]reg_B;
    input GND_net;
    output n30174;
    input clk32MHz;
    input ENCODER0_B_c_0;
    input n16237;
    output [1:0]data_o;
    input ENCODER0_A_c_1;
    input n15721;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3732;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n1;
    wire [2:0]n17;
    
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n30174), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i1405_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(170[42:59])
    defparam i1405_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18623_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i18623_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i18616_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i18616_2_lut.LUT_INIT = 16'h6666;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1198__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n1), .R(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n16237));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i2_3_lut_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[2]), 
            .I3(GND_net), .O(n30174));
    defparam i2_3_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n15721));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1198__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1198__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (GND_net, timer, \neo_pixel_transmitter.done , clk32MHz, 
            \state[1] , start, n28731, n26593, VCC_net, n28597, 
            n15451, \state_3__N_372[1] , \neo_pixel_transmitter.t0 , neopxl_color, 
            LED_c, NEOPXL_c, n15761, n15760, n15759, n15758, n15757, 
            n15756, n15755, n15754, n15753, n15752, n15751, n15750, 
            n15749, n15748, n15747, n15746, n15745, n15744, n15743, 
            n15742, n15741, n15740, n15739, n15738, n15737, n15736, 
            n15735, n15734, n15733, n15732, n15731, n26505, n29426, 
            n15726, n15704) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [31:0]timer;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output \state[1] ;
    output start;
    output n28731;
    output n26593;
    input VCC_net;
    output n28597;
    output n15451;
    output \state_3__N_372[1] ;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input [23:0]neopxl_color;
    input LED_c;
    output NEOPXL_c;
    input n15761;
    input n15760;
    input n15759;
    input n15758;
    input n15757;
    input n15756;
    input n15755;
    input n15754;
    input n15753;
    input n15752;
    input n15751;
    input n15750;
    input n15749;
    input n15748;
    input n15747;
    input n15746;
    input n15745;
    input n15744;
    input n15743;
    input n15742;
    input n15741;
    input n15740;
    input n15739;
    input n15738;
    input n15737;
    input n15736;
    input n15735;
    input n15734;
    input n15733;
    input n15732;
    input n15731;
    input n26505;
    output n29426;
    input n15726;
    input n15704;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]n133;
    
    wire n23951, n24214, n3090, n3116, n24215, n2001, n2008, n1994, 
        n1995, n27;
    wire [31:0]n255;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n23473, n2398, n2299, n2324, n23445, n23952, \neo_pixel_transmitter.done_N_580 , 
        n32240, n15508, n15621, n24147, n2906, n2918, n24148, 
        n2701, n2602, n2621, n24082, n47, n3091, n24213, n3006, 
        n2907, n24146, n1304, n1305, n10, n24083, n1306, n1309, 
        n12, n2702, n2603, n24081, n1302, n1303, n1308, n16, 
        n23950, n1307, n1301, n1334, n1928, n31927, n1829, n31942, 
        n1037, n31943, n3007, n2908, n24145, n23949, n14186, n28657, 
        n24851;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire n28723, n23948, n2703, n2604, n24080, n7, n14300, n23947, 
        n23946, n2704, n2605, n24079, n23945, n23944, n23472, 
        n23943, n23471, n23470, n23446, n23942, n2406, n2307, 
        n23437, n2399, n2300, n23444, n45, n3092, n24212, n3008, 
        n2909, n31922, n24144, n2705, n2606, n24078, n23941, n2291, 
        n2192, n2225, n23675, n2292, n2193, n23674, n23940, n2293, 
        n2194, n23673, n2294, n2195, n23672, n23939, n2295, n2196, 
        n23671, n2296, n2197, n23670, n23938, n2297, n2198, n23669, 
        n2706, n2607, n24077, n2298, n2199, n23668, n23937, n2200, 
        n23667, n2201, n23666, n2301, n2202, n23665, n23469, n2302, 
        n2203, n23664, n1202, n1235, n23936, n23438, n2400, n23443, 
        n2303, n2204, n23663, n1203, n23935, n23468, n2304, n2205, 
        n23662, n23467, n2305, n2206, n23661, n3009, n2707, n2608, 
        n24076, n1204, n23934, n1895, n23816, n2306, n2207, n23660, 
        n1896, n23815, n2208, n23659, n1996, n1897, n23814, n1205, 
        n23933, n2308, n2209, n31925, n23658, n1997, n1898, n23813, 
        n2309, n1998, n1899, n23812, n1206, n23932, n1999, n1900, 
        n23811, n2000, n1901, n23810, n1207, n23931, n1902, n23809, 
        n2002, n1903, n23808, n2708, n2609, n31923, n24075, n1208, 
        n23930, n2003, n1904, n23807, n2004, n1905, n23806, n1209, 
        n31926, n23929, n2005, n1906, n23805, n2006, n1907, n23804, 
        n2007, n1908, n23803, n23466, n1909, n23802, n1400, n23928, 
        n2009, n1401, n23927, n2407, n23436, n2093, n2027, n23801, 
        n43, n3093, n24211, n2885, n2786, n2819, n24143, n2709, 
        n2094, n23800, n1402, n23926, n2095, n23799, n2096, n23798, 
        n1403, n23925, n2097, n23797, n2098, n23796, n1404, n23924, 
        n2099, n23795, n2100, n23794, n1405, n23923, n2101, n23793, 
        n2886, n2787, n24142, n2588, n2489, n2522, n24074, n2102, 
        n23792, n1406, n23922, n2103, n23791, n2104, n23790, n1407, 
        n23921, n2105, n23789, n2589, n2490, n24073, n2106, n23788, 
        n2401, n23442, n1408, n31928, n23920, n2107, n23787, n23465, 
        n2402, n23441, n23464, n2108, n31929, n23786, n2423, n31938, 
        n1109, n19749, n1105, n1103, n1108, n12_adj_4609, n1107, 
        n1106, n1104, n1136, n1806, n1803, n1798, n1805, n24, 
        n1808, n1804, n1802, n1807, n22, n1800, n1799, n1797, 
        n1801, n23, n1796, n1809, n21, n31941, n1409, n2109, 
        n23463, n2;
    wire [31:0]n971;
    
    wire n1007, n2126, n23785, n23784, n31408, n2408, n31924, 
        n23435, n41, n3094, n24210, n31068, n19831, n28727, n31409, 
        n28787, \neo_pixel_transmitter.done_N_586 , n35, n27_adj_4610, 
        n25, n63, n28, n51, n59, n11, n26, n57, n33, n29, 
        n27_adj_4611, n49, n15, n61, n25_adj_4612, n30044, n3209, 
        n19727, n17, n19, n37, n29685, n31, n55, n16_adj_4613, 
        n23_adj_4614, n39, n53, n17_adj_4615, n21_adj_4616, n13, 
        n24935, n25270, n1006, n1499, n1433, n23919, n1009, n12921, 
        n1008, n906, n1005, n15566, n905, n28613, n8, n30359, 
        n6, n4, n1730, n31937, n23462;
    wire [31:0]one_wire_N_523;
    
    wire n14323, n1135, n12074;
    wire [4:0]color_bit_N_566;
    
    wire n32020, n32122, n31090, n32098;
    wire [3:0]state_3__N_372;
    
    wire n2887, n2788, n24141, n2590, n2491, n24072, n2403, n23440, 
        n23783, n3095, n24209, n1500, n23918, n2888, n2789, n24140, 
        n2591, n2492, n24071, n23782, n1501, n23917, n2693, n28_adj_4617, 
        n2699, n2694, n2691, n38, n19737, n2696, n2697, n36, 
        n2700, n42, n2690, n2689, n40, n2687, n2695, n41_adj_4618, 
        n2688, n2698, n2692, n39_adj_4619, n2720, n31930, n3000, 
        n30, n2990, n3003, n2997, n42_adj_4620, n3004, n3002, 
        n2994, n2993, n40_adj_4621, n3001, n3005, n2996, n2988, 
        n45_adj_4622, n23781, n2986, n2984, n2995, n2989, n44, 
        n2999, n2992, n2998, n43_adj_4623, n2991, n47_adj_4624, 
        n2985, n2987, n49_adj_4625, n3017, n31921, n2409, n27_adj_4626, 
        n2390, n2391, n2397, n2394, n33_adj_4627, n2392, n2405, 
        n32, n2396, n31_adj_4628, n2393, n2395, n35_adj_4629, n2404, 
        n37_adj_4630, n31931, n1699, n1709, n17_adj_4631, n1698, 
        n1707, n1703, n1705, n21_adj_4632, n1704, n1701, n1708, 
        n20, n1702, n1697, n24_adj_4633, n1700, n1706, n1532, 
        n31934, n1631, n31936;
    wire [31:0]n1;
    
    wire n1608, n1606, n1604, n1603, n20_adj_4647, n1602, n1609, 
        n13_adj_4648, n1598, n1600, n18, n1605, n1599, n22_adj_4649, 
        n1601, n1607, n1502, n23916, n23780, n2889, n2790, n24139, 
        n838, n2592, n2493, n24070, n23779, n1503, n23915, n23778, 
        n2593, n2494, n24069, n23777, n1504, n23914, n18_adj_4655, 
        n25_adj_4656, n2890, n2791, n24138, n23461, n1505, n23913, 
        n23776, n1506, n23912, n23775, n2594, n2495, n24068, n3096, 
        n24208, n23774, n23773, n2891, n2792, n24137, n1507, n23911, 
        n23772, n23771, n1508, n31933, n23910, n23770, n2595, 
        n2496, n24067, n31932, n23769, n1509, n2892, n2793, n24136, 
        n3097, n24207, n23909, n2596, n2497, n24066, n2893, n2794, 
        n24135, n23460, n31940, n807, n60, n23908, n3098, n24206, 
        n2894, n2795, n24134, n3099, n24205, n2597, n2498, n24065, 
        n23459, n2895, n2796, n24133, n23907, n23458, n3100, n24204, 
        n27_adj_4659, n23611, n23906, n22_adj_4661, n23610, n2601, 
        n36_adj_4662, n25_adj_4663, n2600, n34, n739, n12895, n608, 
        n708, n28641, n19721, n23_adj_4665, n23609, n23457, n25284, 
        n28587, n2896, n2797, n24132, n23456, n28_adj_4668, n23608, 
        n2598, n2499, n24064, n23905, n26_adj_4669, n23607, n40_adj_4671, 
        n21_adj_4672, n23606, n23904, n3101, n24203, n2897, n2798, 
        n24131, n2599, n2500, n24063, n23605, n23903, n23604, 
        n2501, n24062, n23902, n29_adj_4675, n23603, n23901, n23602, 
        n30_adj_4676, n23601, n26_adj_4677, n19_adj_4678, n16_adj_4679, 
        n24_adj_4680, n28_adj_4681, n26_adj_4682, n28_adj_4683, n24_adj_4684, 
        n23600, n25_adj_4685, n23599, n23900, n23598, n2898, n2799, 
        n24130, n23597, n23899, n23596, n23595, n23594, n2502, 
        n24061, n14_adj_4687, n9_adj_4688, n23593, n23898, n23592, 
        n23455, n23897, n28_adj_4689, n32_adj_4690, n30_adj_4691, 
        n31_adj_4692, n29_adj_4693, n23591, n38_adj_4694, n23590, 
        n23439, n23454, n23896, n2503, n24060, n23589, n23895, 
        n23588, n23587, n23894, n9_adj_4695, n23586, n23585, n23893, 
        n23584, n23583, n23892, n23582, n2899, n2800, n24129, 
        n2504, n24059, n24931, n23581, n4_adj_4696, n23891, n23890, 
        n23453, n39_adj_4697, n23889, n3102, n24202, n2900, n2801, 
        n24128, n23888, n23452, n23451, n3103, n24201, n2901, 
        n2802, n24127, n2505, n24058, n23450, n2506, n24057, n23887, 
        n2507, n24056, n23886, n23885, n2902, n2803, n24126, n3104, 
        n24200, n2508, n24055, n18_adj_4698, n17_adj_4699, n19_adj_4700, 
        n2903, n2804, n24125, n2509, n24054, n3105, n24199, n23884, 
        n23883, n3106, n24198, n2904, n2805, n24124, n2905, n2806, 
        n24123, n24053, n23882, n24052, n3107, n24197, n23881, 
        n3108, n24196, n3109, n24195, n2807, n24122, n23449, n2808, 
        n24121, n24051, n23880, n3083, n24194, n2809, n24120, 
        n3084, n24193, n24050, n24119, n24049, n23879, n23878, 
        n3085, n24192, n24118, n3086, n24191, n37_adj_4701, n24117, 
        n24048, n3087, n24190, n3088, n24189, n3089, n24188, n24047, 
        n24046, n33_adj_4702, n24187, n41_adj_4703, n24186, n24116, 
        n38_adj_4704, n43_adj_4705, n40_adj_4706, n46, n24185, n39_adj_4707, 
        n24115, n47_adj_4708, n18_adj_4709, n24045, n20_adj_4710, 
        n19_adj_4711, n24_adj_4712, n34_adj_4713, n19755, n16_adj_4714, 
        n17_adj_4715, n22_adj_4716, n18_adj_4717, n19765, n30_adj_4718, 
        n28_adj_4719, n29_adj_4720, n27_adj_4721, n38_adj_4722, n36_adj_4723, 
        n37_adj_4724, n35_adj_4725, n20_adj_4726, n19_adj_4727, n32_adj_4728, 
        n30_adj_4729, n31_adj_4730, n29_adj_4731, n32233, n30363, 
        n14_adj_4732, n1121, n19684, n4607, n32173, n30471, n32167, 
        n30474, n32119, n32095, n31960, n32017, n24114, n31156, 
        n36_adj_4733, n37_adj_4734, n28653, n27865, n111, n116, 
        n16_adj_4735, n18_adj_4736, n23877, n24184, n24044, n23974, 
        n24113, n23973, n23876, n24183, n24043, n24112, n24182, 
        n24181, n24111, n24042, n23972, n23875, n24041, n24180, 
        n24110, n24179, n24109, n24108, n24107, n24178, n24040, 
        n24177, n24039, n24038, n24176, n24106, n23971, n23874, 
        n23970, n24175, n24105, n24037, n23475, n23476, n24104, 
        n24036, n30218, n24174, n23969, n24173, n24172, n24103, 
        n24035, n23968, n23873, n23872, n24034, n24102, n24171, 
        n24101, n23871, n24170, n24100, n23967, n23870, n31957, 
        n24099, n40_adj_4737, n31939, n24169, n38_adj_4738, n22_adj_4739, 
        n30_adj_4740, n34_adj_4741, n32_adj_4742, n33_adj_4743, n31_adj_4744, 
        n42_adj_4745, n46_adj_4746, n44_adj_4747, n45_adj_4748, n43_adj_4749, 
        n40_adj_4750, n48, n52, n39_adj_4751, n23484, n23448, n23483, 
        n24098, n23966, n23482, n24168, n23869, n24167, n39_adj_4752, 
        n24033, n24032, n23868, n24097, n37_adj_4753, n23481, n23965, 
        n24166, n34_adj_4754, n42_adj_4755, n24165, n24031, n23480, 
        n46_adj_4756, n23964, n23867, n24030, n24096, n23963, n24095, 
        n23866, n33_adj_4757, n24164, n24094, n23962, n24093, n24029, 
        n24163, n24092, n23961, n24162, n23865, n24161, n24160, 
        n23960, n23479, n24159, n24028, n24091, n23959, n24158, 
        n24090, n24027, n24157, n23958, n24156, n24026, n24089, 
        n24088, n24155, n24025, n23957, n23864, n23447, n24154, 
        n24024, n24221, n24220, n23478, n23956, n24219, n24153, 
        n24087, n23863, n23955, n24152, n24023, n24218, n24086, 
        n24151, n23477, n24217, n24150, n24085, n23862, n23954, 
        n23861, n24149, n24084, n24216, n23860, n23953, n23474;
    
    SB_LUT4 timer_1191_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n23951), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_22 (.CI(n24214), .I0(n3090), .I1(n3116), .CO(n24215));
    SB_LUT4 i11_4_lut (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n23473), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n23445), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_17 (.CI(n23951), .I0(GND_net), .I1(timer[15]), 
            .CO(n23952));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n32240), .D(\neo_pixel_transmitter.done_N_580 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n15508), 
            .D(n255[1]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2009_6 (.CI(n24147), .I0(n2906), .I1(n2918), .CO(n24148));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n24082), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n24213), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n24146), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1808_10 (.CI(n24082), .I0(n2602), .I1(n2621), .CO(n24083));
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1306), .I2(n1309), .I3(GND_net), 
            .O(n12));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n24081), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut (.I0(n1302), .I1(n1303), .I2(n1308), .I3(n10), 
            .O(n16));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1191_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n23950), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(n1307), .I1(n16), .I2(n12), .I3(n1301), .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26096_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31927));
    defparam i26096_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_5 (.CI(n24146), .I0(n2907), .I1(n2918), .CO(n24147));
    SB_CARRY timer_1191_add_4_16 (.CI(n23950), .I0(GND_net), .I1(timer[14]), 
            .CO(n23951));
    SB_LUT4 i26111_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31942));
    defparam i26111_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26112_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31943));
    defparam i26112_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n24145), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n23949), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_9 (.CI(n24081), .I0(n2603), .I1(n2621), .CO(n24082));
    SB_LUT4 i22902_4_lut (.I0(n14186), .I1(n28657), .I2(n24851), .I3(state[0]), 
            .O(n28723));
    defparam i22902_4_lut.LUT_INIT = 16'hfaee;
    SB_CARRY timer_1191_add_4_15 (.CI(n23949), .I0(GND_net), .I1(timer[13]), 
            .CO(n23950));
    SB_LUT4 timer_1191_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n23948), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n24080), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_14 (.CI(n23948), .I0(GND_net), .I1(timer[12]), 
            .CO(n23949));
    SB_CARRY mod_5_add_1808_8 (.CI(n24080), .I0(n2604), .I1(n2621), .CO(n24081));
    SB_LUT4 i20_4_lut (.I0(n28723), .I1(\state[1] ), .I2(start), .I3(\neo_pixel_transmitter.done ), 
            .O(n7));
    defparam i20_4_lut.LUT_INIT = 16'hcfcd;
    SB_CARRY mod_5_add_2143_21 (.CI(n24213), .I0(n3091), .I1(n3116), .CO(n24214));
    SB_LUT4 i1_4_lut (.I0(n28731), .I1(n7), .I2(n14300), .I3(\state[1] ), 
            .O(n26593));
    defparam i1_4_lut.LUT_INIT = 16'hccc4;
    SB_LUT4 timer_1191_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n23947), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1191_add_4_13 (.CI(n23947), .I0(GND_net), .I1(timer[11]), 
            .CO(n23948));
    SB_LUT4 timer_1191_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n23946), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n24145), .I0(n2908), .I1(n2918), .CO(n24146));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n24079), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_12 (.CI(n23946), .I0(GND_net), .I1(timer[10]), 
            .CO(n23947));
    SB_LUT4 timer_1191_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n23945), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1191_add_4_11 (.CI(n23945), .I0(GND_net), .I1(timer[9]), 
            .CO(n23946));
    SB_LUT4 timer_1191_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n23944), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_7 (.CI(n24079), .I0(n2605), .I1(n2621), .CO(n24080));
    SB_CARRY timer_1191_add_4_10 (.CI(n23944), .I0(GND_net), .I1(timer[8]), 
            .CO(n23945));
    SB_CARRY add_21_21 (.CI(n23472), .I0(bit_ctr[19]), .I1(GND_net), .CO(n23473));
    SB_LUT4 timer_1191_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n23943), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n23471), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_20 (.CI(n23471), .I0(bit_ctr[18]), .I1(GND_net), .CO(n23472));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n23470), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_19 (.CI(n23470), .I0(bit_ctr[17]), .I1(GND_net), .CO(n23471));
    SB_CARRY timer_1191_add_4_9 (.CI(n23943), .I0(GND_net), .I1(timer[7]), 
            .CO(n23944));
    SB_CARRY mod_5_add_1607_13 (.CI(n23445), .I0(n2299), .I1(n2324), .CO(n23446));
    SB_LUT4 timer_1191_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n23942), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n23437), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n23444), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n23472), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n24212), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n31922), 
            .I3(n24144), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n24078), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_8 (.CI(n23942), .I0(GND_net), .I1(timer[6]), 
            .CO(n23943));
    SB_LUT4 timer_1191_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n23941), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1191_add_4_7 (.CI(n23941), .I0(GND_net), .I1(timer[5]), 
            .CO(n23942));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n23675), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n23674), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n23940), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_19 (.CI(n23674), .I0(n2193), .I1(n2225), .CO(n23675));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n23673), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n24078), .I0(n2606), .I1(n2621), .CO(n24079));
    SB_CARRY timer_1191_add_4_6 (.CI(n23940), .I0(GND_net), .I1(timer[4]), 
            .CO(n23941));
    SB_CARRY mod_5_add_1540_18 (.CI(n23673), .I0(n2194), .I1(n2225), .CO(n23674));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n23672), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n23939), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_17 (.CI(n23672), .I0(n2195), .I1(n2225), .CO(n23673));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n23671), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_5 (.CI(n23939), .I0(GND_net), .I1(timer[3]), 
            .CO(n23940));
    SB_CARRY mod_5_add_1540_16 (.CI(n23671), .I0(n2196), .I1(n2225), .CO(n23672));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n23670), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n23938), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_15 (.CI(n23670), .I0(n2197), .I1(n2225), .CO(n23671));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n23669), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_3 (.CI(n24144), .I0(n2909), .I1(n31922), .CO(n24145));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n24077), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_4 (.CI(n23938), .I0(GND_net), .I1(timer[2]), 
            .CO(n23939));
    SB_CARRY mod_5_add_1540_14 (.CI(n23669), .I0(n2198), .I1(n2225), .CO(n23670));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n23668), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n23937), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_13 (.CI(n23668), .I0(n2199), .I1(n2225), .CO(n23669));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n23667), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_3 (.CI(n23937), .I0(GND_net), .I1(timer[1]), 
            .CO(n23938));
    SB_CARRY mod_5_add_1540_12 (.CI(n23667), .I0(n2200), .I1(n2225), .CO(n23668));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n23666), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_11 (.CI(n23666), .I0(n2201), .I1(n2225), .CO(n23667));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n23665), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n24077), .I0(n2607), .I1(n2621), .CO(n24078));
    SB_CARRY timer_1191_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n23937));
    SB_CARRY mod_5_add_1540_10 (.CI(n23665), .I0(n2202), .I1(n2225), .CO(n23666));
    SB_CARRY mod_5_add_1607_12 (.CI(n23444), .I0(n2300), .I1(n2324), .CO(n23445));
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n23469), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n23664), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n23936), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n23664), .I0(n2203), .I1(n2225), .CO(n23665));
    SB_CARRY mod_5_add_1607_5 (.CI(n23437), .I0(n2307), .I1(n2324), .CO(n23438));
    SB_CARRY add_21_18 (.CI(n23469), .I0(bit_ctr[16]), .I1(GND_net), .CO(n23470));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n23443), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n23663), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n23935), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n23663), .I0(n2204), .I1(n2225), .CO(n23664));
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n23468), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_17 (.CI(n23468), .I0(bit_ctr[15]), .I1(GND_net), .CO(n23469));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n23662), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n23935), .I0(n1203), .I1(n1235), .CO(n23936));
    SB_CARRY mod_5_add_1540_7 (.CI(n23662), .I0(n2205), .I1(n2225), .CO(n23663));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n23467), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_16 (.CI(n23467), .I0(bit_ctr[14]), .I1(GND_net), .CO(n23468));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n23661), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n24212), .I0(n3092), .I1(n3116), .CO(n24213));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n31922), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n24076), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n23934), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n23816), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n23661), .I0(n2206), .I1(n2225), .CO(n23662));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n23660), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n23815), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n23934), .I0(n1204), .I1(n1235), .CO(n23935));
    SB_CARRY mod_5_add_1339_16 (.CI(n23815), .I0(n1896), .I1(n1928), .CO(n23816));
    SB_CARRY mod_5_add_1540_5 (.CI(n23660), .I0(n2207), .I1(n2225), .CO(n23661));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n23659), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n23814), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n23933), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n23814), .I0(n1897), .I1(n1928), .CO(n23815));
    SB_CARRY mod_5_add_1540_4 (.CI(n23659), .I0(n2208), .I1(n2225), .CO(n23660));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n31925), 
            .I3(n23658), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n23813), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n23933), .I0(n1205), .I1(n1235), .CO(n23934));
    SB_CARRY mod_5_add_1339_14 (.CI(n23813), .I0(n1898), .I1(n1928), .CO(n23814));
    SB_CARRY mod_5_add_1540_3 (.CI(n23658), .I0(n2209), .I1(n31925), .CO(n23659));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n31925), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n23812), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n24076), .I0(n2608), .I1(n2621), .CO(n24077));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n23932), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n23812), .I0(n1899), .I1(n1928), .CO(n23813));
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n31925), 
            .CO(n23658));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n23811), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n23932), .I0(n1206), .I1(n1235), .CO(n23933));
    SB_CARRY mod_5_add_1339_12 (.CI(n23811), .I0(n1900), .I1(n1928), .CO(n23812));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n23810), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n23931), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n23810), .I0(n1901), .I1(n1928), .CO(n23811));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n23809), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n23931), .I0(n1207), .I1(n1235), .CO(n23932));
    SB_CARRY mod_5_add_1339_10 (.CI(n23809), .I0(n1902), .I1(n1928), .CO(n23810));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n23808), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n31922), 
            .CO(n24144));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n31923), 
            .I3(n24075), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n23930), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n23808), .I0(n1903), .I1(n1928), .CO(n23809));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n23807), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n23930), .I0(n1208), .I1(n1235), .CO(n23931));
    SB_CARRY mod_5_add_1339_8 (.CI(n23807), .I0(n1904), .I1(n1928), .CO(n23808));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n23806), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n31926), 
            .I3(n23929), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_7 (.CI(n23806), .I0(n1905), .I1(n1928), .CO(n23807));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n23805), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_3 (.CI(n23929), .I0(n1209), .I1(n31926), .CO(n23930));
    SB_CARRY mod_5_add_1339_6 (.CI(n23805), .I0(n1906), .I1(n1928), .CO(n23806));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n23804), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_3 (.CI(n24075), .I0(n2609), .I1(n31923), .CO(n24076));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n31926), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_5 (.CI(n23804), .I0(n1907), .I1(n1928), .CO(n23805));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n23803), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n31926), 
            .CO(n23929));
    SB_CARRY mod_5_add_1339_4 (.CI(n23803), .I0(n1908), .I1(n1928), .CO(n23804));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n23466), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_11 (.CI(n23443), .I0(n2301), .I1(n2324), .CO(n23444));
    SB_CARRY add_21_15 (.CI(n23466), .I0(bit_ctr[13]), .I1(GND_net), .CO(n23467));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n31927), 
            .I3(n23802), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n23928), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_3 (.CI(n23802), .I0(n1909), .I1(n31927), .CO(n23803));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n31927), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n23927), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n31927), 
            .CO(n23802));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n23436), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n23801), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n24211), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n24143), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n31923), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_10 (.CI(n23927), .I0(n1302), .I1(n1334), .CO(n23928));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n23800), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n23800), .I0(n1995), .I1(n2027), .CO(n23801));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n23926), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n23799), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n23799), .I0(n1996), .I1(n2027), .CO(n23800));
    SB_CARRY mod_5_add_937_9 (.CI(n23926), .I0(n1303), .I1(n1334), .CO(n23927));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n23798), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n23798), .I0(n1997), .I1(n2027), .CO(n23799));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n23925), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n23797), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n23797), .I0(n1998), .I1(n2027), .CO(n23798));
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n31923), 
            .CO(n24075));
    SB_CARRY mod_5_add_937_8 (.CI(n23925), .I0(n1304), .I1(n1334), .CO(n23926));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n23796), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n23796), .I0(n1999), .I1(n2027), .CO(n23797));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n23924), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n23795), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n23795), .I0(n2000), .I1(n2027), .CO(n23796));
    SB_CARRY mod_5_add_937_7 (.CI(n23924), .I0(n1305), .I1(n1334), .CO(n23925));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n23794), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n23794), .I0(n2001), .I1(n2027), .CO(n23795));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n23923), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n23793), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n23793), .I0(n2002), .I1(n2027), .CO(n23794));
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n24142), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n24074), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n23923), .I0(n1306), .I1(n1334), .CO(n23924));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n23792), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n23792), .I0(n2003), .I1(n2027), .CO(n23793));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n23922), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n23791), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n23791), .I0(n2004), .I1(n2027), .CO(n23792));
    SB_CARRY mod_5_add_937_5 (.CI(n23922), .I0(n1307), .I1(n1334), .CO(n23923));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n23790), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n23790), .I0(n2005), .I1(n2027), .CO(n23791));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n23921), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n23789), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n23789), .I0(n2006), .I1(n2027), .CO(n23790));
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n24073), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n23921), .I0(n1308), .I1(n1334), .CO(n23922));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n23788), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n23442), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_5 (.CI(n23788), .I0(n2007), .I1(n2027), .CO(n23789));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n31928), 
            .I3(n23920), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n23787), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n23465), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n23442), .I0(n2302), .I1(n2324), .CO(n23443));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n23441), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n23787), .I0(n2008), .I1(n2027), .CO(n23788));
    SB_CARRY add_21_14 (.CI(n23465), .I0(bit_ctr[12]), .I1(GND_net), .CO(n23466));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n23464), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_4 (.CI(n23436), .I0(n2308), .I1(n2324), .CO(n23437));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n31929), 
            .I3(n23786), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n23920), .I0(n1309), .I1(n31928), .CO(n23921));
    SB_CARRY mod_5_add_1406_3 (.CI(n23786), .I0(n2009), .I1(n31929), .CO(n23787));
    SB_LUT4 i26107_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31938));
    defparam i26107_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n15508), 
            .D(n255[31]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n15508), 
            .D(n255[30]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i15208_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n19749));
    defparam i15208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n19749), .I2(n1103), .I3(n1108), 
            .O(n12_adj_4609));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1107), .I1(n12_adj_4609), .I2(n1106), .I3(n1104), 
            .O(n1136));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1489 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22));
    defparam i8_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n21));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut (.I0(n21), .I1(n23), .I2(n22), .I3(n24), .O(n1829));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26110_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31941));
    defparam i26110_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n31928), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_9 (.CI(n23441), .I0(n2303), .I1(n2324), .CO(n23442));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n31929), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_13 (.CI(n23464), .I0(bit_ctr[11]), .I1(GND_net), .CO(n23465));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n23463), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_19 (.CI(n24211), .I0(n3093), .I1(n3116), .CO(n24212));
    SB_CARRY mod_5_add_1942_25 (.CI(n24142), .I0(n2787), .I1(n2819), .CO(n24143));
    SB_CARRY mod_5_add_1741_22 (.CI(n24073), .I0(n2490), .I1(n2522), .CO(n24074));
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n31929), 
            .CO(n23786));
    SB_LUT4 i26046_2_lut (.I0(n2), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i26046_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n23785), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n31928), 
            .CO(n23920));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n23784), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25757_4_lut (.I0(n24851), .I1(n28657), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n31408));
    defparam i25757_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n31924), 
            .I3(n23435), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n24210), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25505_2_lut (.I0(n28657), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n31068));
    defparam i25505_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53_4_lut (.I0(n31068), .I1(n19831), .I2(\state[1] ), .I3(n14186), 
            .O(n28727));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n28727), .I1(n31409), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n28787));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_586 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut (.I0(n35), .I1(n27_adj_4610), .I2(n25), .I3(n63), 
            .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1490 (.I0(n51), .I1(n59), .I2(n11), .I3(n47), 
            .O(n26));
    defparam i10_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1491 (.I0(n57), .I1(n33), .I2(n43), .I3(n29), 
            .O(n27_adj_4611));
    defparam i11_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1492 (.I0(n49), .I1(n15), .I2(n41), .I3(n61), 
            .O(n25_adj_4612));
    defparam i9_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25_adj_4612), .I1(n27_adj_4611), .I2(n26), 
            .I3(n28), .O(n30044));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15186_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n19727));
    defparam i15186_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(n17), .I1(n19), .I2(n37), .I3(n45), .O(n29685));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1493 (.I0(n31), .I1(n19727), .I2(n30044), .I3(n55), 
            .O(n16_adj_4613));
    defparam i6_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1494 (.I0(n23_adj_4614), .I1(n39), .I2(n29685), 
            .I3(n53), .O(n17_adj_4615));
    defparam i7_4_lut_adj_1494.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1495 (.I0(n17_adj_4615), .I1(n21_adj_4616), .I2(n16_adj_4613), 
            .I3(n13), .O(n24935));
    defparam i9_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1496 (.I0(bit_ctr[3]), .I1(n24935), .I2(GND_net), 
            .I3(GND_net), .O(n25270));
    defparam i1_2_lut_adj_1496.LUT_INIT = 16'h6666;
    SB_LUT4 i26044_2_lut (.I0(n2), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i26044_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n23919), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n23784), .I0(n2094), .I1(n2126), .CO(n23785));
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n12921), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_3_lut_adj_1497 (.I0(n15566), .I1(n905), .I2(n28613), .I3(GND_net), 
            .O(n8));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut_adj_1497.LUT_INIT = 16'h0101;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n8), .I2(n906), .I3(n12921), 
            .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h040c;
    SB_LUT4 i24528_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n30359));
    defparam i24528_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut_adj_1498 (.I0(n2), .I1(n6), .I2(n1005), .I3(n30359), 
            .O(n1037));
    defparam i3_4_lut_adj_1498.LUT_INIT = 16'hfdfc;
    SB_LUT4 i26062_2_lut (.I0(n2), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4));   // verilog/neopixel.v(22[26:36])
    defparam i26062_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i26106_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31937));
    defparam i26106_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_12 (.CI(n23463), .I0(bit_ctr[10]), .I1(GND_net), .CO(n23464));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n23462), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22907_4_lut (.I0(n14186), .I1(n24851), .I2(n28657), .I3(state[0]), 
            .O(n28731));
    defparam i22907_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i15289_4_lut (.I0(one_wire_N_523[9]), .I1(n14323), .I2(one_wire_N_523[11]), 
            .I3(one_wire_N_523[10]), .O(n19831));
    defparam i15289_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i233_2_lut (.I0(n19831), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1135));   // verilog/neopixel.v(103[9] 111[12])
    defparam i233_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1499 (.I0(n12074), .I1(n1135), .I2(\state[1] ), 
            .I3(state[0]), .O(n28597));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1499.LUT_INIT = 16'h0535;
    SB_LUT4 i1_4_lut_adj_1500 (.I0(state[0]), .I1(n12074), .I2(n1135), 
            .I3(\state[1] ), .O(n15451));
    defparam i1_4_lut_adj_1500.LUT_INIT = 16'haf33;
    SB_LUT4 mod_5_i2239_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n24935), 
            .I3(GND_net), .O(color_bit_N_566[4]));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2239_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i25751_4_lut (.I0(n32020), .I1(n25270), .I2(n32122), .I3(bit_ctr[2]), 
            .O(n31090));
    defparam i25751_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i14649_4_lut (.I0(n32098), .I1(\state_3__N_372[1] ), .I2(n31090), 
            .I3(color_bit_N_566[4]), .O(state_3__N_372[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i14649_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_21_11 (.CI(n23462), .I0(bit_ctr[9]), .I1(GND_net), .CO(n23463));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n24141), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n24072), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n24210), .I0(n3094), .I1(n3116), .CO(n24211));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n23440), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n24141), .I0(n2788), .I1(n2819), .CO(n24142));
    SB_CARRY mod_5_add_1741_21 (.CI(n24072), .I0(n2491), .I1(n2522), .CO(n24073));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n23783), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n15508), 
            .D(n255[29]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n24209), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n23918), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n24140), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n24071), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n23918), .I0(n1401), .I1(n1433), .CO(n23919));
    SB_CARRY mod_5_add_1473_17 (.CI(n23783), .I0(n2095), .I1(n2126), .CO(n23784));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n23782), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n23917), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n23782), .I0(n2096), .I1(n2126), .CO(n23783));
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n15508), 
            .D(n255[28]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n15508), 
            .D(n255[27]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n15508), 
            .D(n255[26]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4617));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1501 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38));
    defparam i15_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i15196_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n19737));
    defparam i15196_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1502 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n19737), 
            .O(n36));
    defparam i13_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n2700), .I1(n38), .I2(n28_adj_4617), .I3(n2705), 
            .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n2687), .I1(n36), .I2(n2703), .I3(n2695), 
            .O(n41_adj_4618));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4619));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_4619), .I1(n41_adj_4618), .I2(n40), 
            .I3(n42), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26099_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31930));
    defparam i26099_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut (.I0(n3000), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n30));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i16_4_lut_adj_1503 (.I0(n2990), .I1(n3003), .I2(n2997), .I3(n3006), 
            .O(n42_adj_4620));
    defparam i16_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n3004), .I1(n3002), .I2(n2994), .I3(n2993), 
            .O(n40_adj_4621));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1504 (.I0(n3001), .I1(n3005), .I2(n2996), .I3(n2988), 
            .O(n45_adj_4622));
    defparam i19_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n23781), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18_4_lut_adj_1505 (.I0(n2986), .I1(n2984), .I2(n2995), .I3(n2989), 
            .O(n44));
    defparam i18_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1506 (.I0(n2999), .I1(n2992), .I2(n2998), .I3(n3008), 
            .O(n43_adj_4623));
    defparam i17_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n2991), .I1(n42_adj_4620), .I2(n30), .I3(n3007), 
            .O(n47_adj_4624));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n45_adj_4622), .I1(n2985), .I2(n40_adj_4621), 
            .I3(n2987), .O(n49_adj_4625));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n49_adj_4625), .I1(n47_adj_4624), .I2(n43_adj_4623), 
            .I3(n44), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26090_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31921));
    defparam i26090_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_3_lut_adj_1507 (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), 
            .I3(GND_net), .O(n27_adj_4626));
    defparam i7_3_lut_adj_1507.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1508 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4627));
    defparam i13_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1509 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32));
    defparam i12_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1510 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4628));
    defparam i11_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1511 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4629));
    defparam i15_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1512 (.I0(n33_adj_4627), .I1(n27_adj_4626), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4630));
    defparam i17_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1513 (.I0(n37_adj_4630), .I1(n35_adj_4629), .I2(n31_adj_4628), 
            .I3(n32), .O(n2423));
    defparam i19_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i26100_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31931));
    defparam i26100_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1514 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_4631));
    defparam i4_3_lut_adj_1514.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1515 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4632));
    defparam i8_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1516 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20));
    defparam i7_3_lut_adj_1516.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1517 (.I0(n21_adj_4632), .I1(n17_adj_4631), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4633));
    defparam i11_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1518 (.I0(n1700), .I1(n24_adj_4633), .I2(n20), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i26103_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31934));
    defparam i26103_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26105_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31936));
    defparam i26105_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1004_10 (.CI(n23917), .I0(n1402), .I1(n1433), .CO(n23918));
    SB_LUT4 i8_4_lut_adj_1519 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4647));
    defparam i8_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), .I3(GND_net), 
            .O(n13_adj_4648));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1520 (.I0(n13_adj_4648), .I1(n20_adj_4647), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4649));
    defparam i10_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1521 (.I0(n1601), .I1(n22_adj_4649), .I2(n18), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_23 (.CI(n24140), .I0(n2789), .I1(n2819), .CO(n24141));
    SB_CARRY mod_5_add_1741_20 (.CI(n24071), .I0(n2492), .I1(n2522), .CO(n24072));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n23916), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_17 (.CI(n24209), .I0(n3095), .I1(n3116), .CO(n24210));
    SB_CARRY mod_5_add_1473_15 (.CI(n23781), .I0(n2097), .I1(n2126), .CO(n23782));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n23780), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n24139), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1522 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n12921));
    defparam i1_2_lut_adj_1522.LUT_INIT = 16'h9999;
    SB_CARRY mod_5_add_1942_22 (.CI(n24139), .I0(n2790), .I1(n2819), .CO(n24140));
    SB_CARRY mod_5_add_1473_14 (.CI(n23780), .I0(n2098), .I1(n2126), .CO(n23781));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n24070), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n24070), .I0(n2493), .I1(n2522), .CO(n24071));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n23779), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n23916), .I0(n1403), .I1(n1433), .CO(n23917));
    SB_CARRY mod_5_add_1473_13 (.CI(n23779), .I0(n2099), .I1(n2126), .CO(n23780));
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n23915), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n23778), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n23778), .I0(n2100), .I1(n2126), .CO(n23779));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n24069), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1004_8 (.CI(n23915), .I0(n1404), .I1(n1433), .CO(n23916));
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n15508), 
            .D(n255[8]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n23777), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n23914), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_4_lut_adj_1523 (.I0(bit_ctr[15]), .I1(n18_adj_4655), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4656));
    defparam i9_4_lut_adj_1523.LUT_INIT = 16'hfefc;
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n15508), 
            .D(n255[25]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n24138), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n15508), 
            .D(n255[7]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_7 (.CI(n23914), .I0(n1405), .I1(n1433), .CO(n23915));
    SB_CARRY mod_5_add_1741_18 (.CI(n24069), .I0(n2494), .I1(n2522), .CO(n24070));
    SB_CARRY mod_5_add_1473_11 (.CI(n23777), .I0(n2101), .I1(n2126), .CO(n23778));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n23461), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n23913), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n24138), .I0(n2791), .I1(n2819), .CO(n24139));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n23776), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_10 (.CI(n23461), .I0(bit_ctr[8]), .I1(GND_net), .CO(n23462));
    SB_CARRY mod_5_add_1473_10 (.CI(n23776), .I0(n2102), .I1(n2126), .CO(n23777));
    SB_CARRY mod_5_add_1004_6 (.CI(n23913), .I0(n1406), .I1(n1433), .CO(n23914));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n23912), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n23775), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n24068), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n24208), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n23775), .I0(n2103), .I1(n2126), .CO(n23776));
    SB_CARRY mod_5_add_1004_5 (.CI(n23912), .I0(n1407), .I1(n1433), .CO(n23913));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n23774), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n23774), .I0(n2104), .I1(n2126), .CO(n23775));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n23773), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n24137), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n24068), .I0(n2495), .I1(n2522), .CO(n24069));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n23911), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n23773), .I0(n2105), .I1(n2126), .CO(n23774));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n23772), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n23911), .I0(n1408), .I1(n1433), .CO(n23912));
    SB_CARRY mod_5_add_1473_6 (.CI(n23772), .I0(n2106), .I1(n2126), .CO(n23773));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n23771), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n31933), 
            .I3(n23910), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_5 (.CI(n23771), .I0(n2107), .I1(n2126), .CO(n23772));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n23770), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_3 (.CI(n23910), .I0(n1409), .I1(n31933), .CO(n23911));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n24067), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n23770), .I0(n2108), .I1(n2126), .CO(n23771));
    SB_CARRY mod_5_add_1942_20 (.CI(n24137), .I0(n2792), .I1(n2819), .CO(n24138));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n31932), 
            .I3(n23769), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n31933), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n24136), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n31933), 
            .CO(n23910));
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_16 (.CI(n24208), .I0(n3096), .I1(n3116), .CO(n24209));
    SB_CARRY mod_5_add_1473_3 (.CI(n23769), .I0(n2109), .I1(n31932), .CO(n23770));
    SB_CARRY mod_5_add_1741_16 (.CI(n24067), .I0(n2496), .I1(n2522), .CO(n24068));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n24207), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n31932), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n23909), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n31932), 
            .CO(n23769));
    SB_CARRY mod_5_add_1942_19 (.CI(n24136), .I0(n2793), .I1(n2819), .CO(n24137));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n24066), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n24135), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n23460), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26109_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31940));
    defparam i26109_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_15 (.CI(n24207), .I0(n3097), .I1(n3116), .CO(n24208));
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n23908), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n24206), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n24135), .I0(n2794), .I1(n2819), .CO(n24136));
    SB_CARRY mod_5_add_2143_14 (.CI(n24206), .I0(n3098), .I1(n3116), .CO(n24207));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n24134), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n15508), 
            .D(n255[24]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_15 (.CI(n24066), .I0(n2497), .I1(n2522), .CO(n24067));
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n15508), 
            .D(n255[23]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n24205), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n24134), .I0(n2795), .I1(n2819), .CO(n24135));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n24065), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_9 (.CI(n23460), .I0(bit_ctr[7]), .I1(GND_net), .CO(n23461));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n23459), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_13 (.CI(n24205), .I0(n3099), .I1(n3116), .CO(n24206));
    SB_CARRY mod_5_add_1741_14 (.CI(n24065), .I0(n2498), .I1(n2522), .CO(n24066));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n24133), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n23908), .I0(n1500), .I1(n1532), .CO(n23909));
    SB_CARRY add_21_8 (.CI(n23459), .I0(bit_ctr[6]), .I1(GND_net), .CO(n23460));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n23907), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n23458), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_11 (.CI(n23907), .I0(n1501), .I1(n1532), .CO(n23908));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n24204), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_523[16]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n23611), .O(n27_adj_4659)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n23906), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_523[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n23610), .O(n22_adj_4661)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i14_4_lut_adj_1524 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4662));
    defparam i14_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1525 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4663));
    defparam i3_3_lut_adj_1525.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1526 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34));
    defparam i12_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_7 (.CI(n23458), .I0(bit_ctr[5]), .I1(GND_net), .CO(n23459));
    SB_CARRY sub_14_add_2_32 (.CI(n23610), .I0(timer[30]), .I1(n1[30]), 
            .CO(n23611));
    SB_CARRY mod_5_add_1071_10 (.CI(n23906), .I0(n1502), .I1(n1532), .CO(n23907));
    SB_LUT4 i1_2_lut_adj_1527 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n12895));
    defparam i1_2_lut_adj_1527.LUT_INIT = 16'h6666;
    SB_LUT4 i15136_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i15136_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i26095_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31926));
    defparam i26095_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n608), .I2(n28641), .I3(n19721), 
            .O(n739));
    defparam i2_4_lut.LUT_INIT = 16'h0105;
    SB_CARRY mod_5_add_1942_16 (.CI(n24133), .I0(n2796), .I1(n2819), .CO(n24134));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_523[22]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n23609), .O(n23_adj_4665)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n23457), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_6 (.CI(n23457), .I0(bit_ctr[4]), .I1(GND_net), .CO(n23458));
    SB_LUT4 i25575_3_lut (.I0(n25284), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n28587));
    defparam i25575_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n28641), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n24132), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n23456), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_31 (.CI(n23609), .I0(timer[29]), .I1(n1[29]), 
            .CO(n23610));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26092_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31923));
    defparam i26092_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_12 (.CI(n24204), .I0(n3100), .I1(n3116), .CO(n24205));
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_523[18]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n23608), .O(n28_adj_4668)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1942_15 (.CI(n24132), .I0(n2797), .I1(n2819), .CO(n24133));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n24064), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n23905), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_30 (.CI(n23608), .I0(timer[28]), .I1(n1[28]), 
            .CO(n23609));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_523[25]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n23607), .O(n26_adj_4669)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1071_9 (.CI(n23905), .I0(n1503), .I1(n1532), .CO(n23906));
    SB_CARRY mod_5_add_1741_13 (.CI(n24064), .I0(n2499), .I1(n2522), .CO(n24065));
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n15508), 
            .D(n255[22]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n15508), 
            .D(n255[21]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i18_4_lut_adj_1528 (.I0(n25_adj_4663), .I1(n36_adj_4662), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4671));
    defparam i18_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_29 (.CI(n23607), .I0(timer[27]), .I1(n1[27]), 
            .CO(n23608));
    SB_LUT4 sub_14_add_2_28_lut (.I0(one_wire_N_523[17]), .I1(timer[26]), 
            .I2(n1[26]), .I3(n23606), .O(n21_adj_4672)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n23904), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_28 (.CI(n23606), .I0(timer[26]), .I1(n1[26]), 
            .CO(n23607));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n24203), .O(n27_adj_4610)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n23904), .I0(n1504), .I1(n1532), .CO(n23905));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n24131), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n24131), .I0(n2798), .I1(n2819), .CO(n24132));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n24063), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n23605), .O(one_wire_N_523[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n23903), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_27 (.CI(n23605), .I0(timer[25]), .I1(n1[25]), 
            .CO(n23606));
    SB_CARRY mod_5_add_1741_12 (.CI(n24063), .I0(n2500), .I1(n2522), .CO(n24064));
    SB_CARRY mod_5_add_1071_7 (.CI(n23903), .I0(n1505), .I1(n1532), .CO(n23904));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n23604), .O(one_wire_N_523[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_26 (.CI(n23604), .I0(timer[24]), .I1(n1[24]), 
            .CO(n23605));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n24062), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n23902), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_523[14]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n23603), .O(n29_adj_4675)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_5 (.CI(n23456), .I0(bit_ctr[3]), .I1(GND_net), .CO(n23457));
    SB_CARRY sub_14_add_2_25 (.CI(n23603), .I0(timer[23]), .I1(n1[23]), 
            .CO(n23604));
    SB_CARRY mod_5_add_1071_6 (.CI(n23902), .I0(n1506), .I1(n1532), .CO(n23903));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n23901), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n1[22]), 
            .I3(n23602), .O(one_wire_N_523[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_24 (.CI(n23602), .I0(timer[22]), .I1(n1[22]), 
            .CO(n23603));
    SB_CARRY mod_5_add_1071_5 (.CI(n23901), .I0(n1507), .I1(n1532), .CO(n23902));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_523[15]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n23601), .O(n30_adj_4676)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i26094_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31925));
    defparam i26094_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_4_lut_adj_1529 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4677));
    defparam i11_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1530 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19_adj_4678));
    defparam i4_3_lut_adj_1530.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4679));
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1532 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4680));
    defparam i9_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1533 (.I0(n19_adj_4678), .I1(n26_adj_4677), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4681));
    defparam i13_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1534 (.I0(n1896), .I1(n28_adj_4681), .I2(n24_adj_4680), 
            .I3(n16_adj_4679), .O(n1928));
    defparam i14_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1535 (.I0(n25_adj_4656), .I1(n27), .I2(n26_adj_4682), 
            .I3(n28_adj_4683), .O(n2027));
    defparam i15_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_23 (.CI(n23601), .I0(timer[21]), .I1(n1[21]), 
            .CO(n23602));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_523[12]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n23600), .O(n24_adj_4684)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n23600), .I0(timer[20]), .I1(n1[20]), 
            .CO(n23601));
    SB_LUT4 sub_14_add_2_21_lut (.I0(one_wire_N_523[13]), .I1(timer[19]), 
            .I2(n1[19]), .I3(n23599), .O(n25_adj_4685)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n23900), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_21 (.CI(n23599), .I0(timer[19]), .I1(n1[19]), 
            .CO(n23600));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n23598), .O(one_wire_N_523[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n24130), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n24062), .I0(n2501), .I1(n2522), .CO(n24063));
    SB_CARRY mod_5_add_1071_4 (.CI(n23900), .I0(n1508), .I1(n1532), .CO(n23901));
    SB_CARRY sub_14_add_2_20 (.CI(n23598), .I0(timer[18]), .I1(n1[18]), 
            .CO(n23599));
    SB_LUT4 sub_14_add_2_19_lut (.I0(GND_net), .I1(timer[17]), .I2(n1[17]), 
            .I3(n23597), .O(one_wire_N_523[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n31934), 
            .I3(n23899), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_19 (.CI(n23597), .I0(timer[17]), .I1(n1[17]), 
            .CO(n23598));
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n23596), .O(one_wire_N_523[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n23596), .I0(timer[16]), .I1(n1[16]), 
            .CO(n23597));
    SB_CARRY mod_5_add_1071_3 (.CI(n23899), .I0(n1509), .I1(n31934), .CO(n23900));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n23595), .O(one_wire_N_523[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_17 (.CI(n23595), .I0(timer[15]), .I1(n1[15]), 
            .CO(n23596));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n31934), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n23594), .O(one_wire_N_523[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_16 (.CI(n23594), .I0(timer[14]), .I1(n1[14]), 
            .CO(n23595));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n24061), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n24061), .I0(n2502), .I1(n2522), .CO(n24062));
    SB_LUT4 i6_4_lut_adj_1536 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4687));
    defparam i6_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n31934), 
            .CO(n23899));
    SB_LUT4 i1_3_lut_adj_1537 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4688));
    defparam i1_3_lut_adj_1537.LUT_INIT = 16'hecec;
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n23593), .O(one_wire_N_523[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_15 (.CI(n23593), .I0(timer[13]), .I1(n1[13]), 
            .CO(n23594));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n23898), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n23592), .O(one_wire_N_523[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n23455), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_8 (.CI(n23440), .I0(n2304), .I1(n2324), .CO(n23441));
    SB_CARRY sub_14_add_2_14 (.CI(n23592), .I0(timer[12]), .I1(n1[12]), 
            .CO(n23593));
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n23897), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n15508), 
            .D(n255[0]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1538 (.I0(n9_adj_4688), .I1(n14_adj_4687), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1539 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4689));
    defparam i10_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1540 (.I0(n2203), .I1(n28_adj_4689), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4690));
    defparam i14_4_lut_adj_1540.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1541 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4691));
    defparam i12_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1542 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4692));
    defparam i13_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1543 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4693));
    defparam i11_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1544 (.I0(n29_adj_4693), .I1(n31_adj_4692), .I2(n30_adj_4691), 
            .I3(n32_adj_4690), .O(n2225));
    defparam i17_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i26091_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31922));
    defparam i26091_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n23591), .O(one_wire_N_523[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_adj_1545 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4694));
    defparam i16_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_4 (.CI(n23455), .I0(bit_ctr[2]), .I1(GND_net), .CO(n23456));
    SB_CARRY mod_5_add_1607_3 (.CI(n23435), .I0(n2309), .I1(n31924), .CO(n23436));
    SB_CARRY sub_14_add_2_13 (.CI(n23591), .I0(timer[11]), .I1(n1[11]), 
            .CO(n23592));
    SB_CARRY mod_5_add_1138_13 (.CI(n23897), .I0(n1599), .I1(n1631), .CO(n23898));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n23590), .O(one_wire_N_523[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n23439), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n23454), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_3 (.CI(n23454), .I0(bit_ctr[1]), .I1(GND_net), .CO(n23455));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n23896), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n23454));
    SB_CARRY sub_14_add_2_12 (.CI(n23590), .I0(timer[10]), .I1(n1[10]), 
            .CO(n23591));
    SB_CARRY mod_5_add_2143_11 (.CI(n24203), .I0(n3101), .I1(n3116), .CO(n24204));
    SB_CARRY mod_5_add_1942_13 (.CI(n24130), .I0(n2799), .I1(n2819), .CO(n24131));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n24060), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n23896), .I0(n1600), .I1(n1631), .CO(n23897));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n23589), .O(one_wire_N_523[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n23589), .I0(timer[9]), .I1(n1[9]), 
            .CO(n23590));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n23895), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n23588), .O(one_wire_N_523[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n23588), .I0(timer[8]), .I1(n1[8]), 
            .CO(n23589));
    SB_CARRY mod_5_add_1138_11 (.CI(n23895), .I0(n1601), .I1(n1631), .CO(n23896));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n23587), .O(one_wire_N_523[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n23587), .I0(timer[7]), .I1(n1[7]), .CO(n23588));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n23894), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_523[9]), .I1(timer[6]), .I2(n1[6]), 
            .I3(n23586), .O(n9_adj_4695)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_8 (.CI(n23586), .I0(timer[6]), .I1(n1[6]), .CO(n23587));
    SB_CARRY mod_5_add_1741_9 (.CI(n24060), .I0(n2503), .I1(n2522), .CO(n24061));
    SB_CARRY mod_5_add_1138_10 (.CI(n23894), .I0(n1602), .I1(n1631), .CO(n23895));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n23585), .O(one_wire_N_523[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n23585), .I0(timer[5]), .I1(n1[5]), .CO(n23586));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n23893), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n23584), .O(one_wire_N_523[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n23584), .I0(timer[4]), .I1(n1[4]), .CO(n23585));
    SB_CARRY mod_5_add_1138_9 (.CI(n23893), .I0(n1603), .I1(n1631), .CO(n23894));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n23583), .O(one_wire_N_523[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n23583), .I0(timer[3]), .I1(n1[3]), .CO(n23584));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n23892), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n23582), .O(one_wire_N_523[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n23582), .I0(timer[2]), .I1(n1[2]), .CO(n23583));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n24129), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n24059), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n23892), .I0(n1604), .I1(n1631), .CO(n23893));
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4696), .I1(timer[1]), .I2(n1[1]), 
            .I3(n23581), .O(n24931)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_3 (.CI(n23581), .I0(timer[1]), .I1(n1[1]), .CO(n23582));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n23891), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_523[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_adj_4696)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n23581));
    SB_CARRY mod_5_add_1138_7 (.CI(n23891), .I0(n1605), .I1(n1631), .CO(n23892));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n23890), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n24059), .I0(n2504), .I1(n2522), .CO(n24060));
    SB_CARRY mod_5_add_1138_6 (.CI(n23890), .I0(n1606), .I1(n1631), .CO(n23891));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n23453), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4697));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n23889), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n24202), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_12 (.CI(n24129), .I0(n2800), .I1(n2819), .CO(n24130));
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_10 (.CI(n24202), .I0(n3102), .I1(n3116), .CO(n24203));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n24128), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n23889), .I0(n1607), .I1(n1631), .CO(n23890));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n23888), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n23452), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n23439), .I0(n2305), .I1(n2324), .CO(n23440));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n23438), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n23452), .I0(n2292), .I1(n2324), .CO(n23453));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n23451), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n23451), .I0(n2293), .I1(n2324), .CO(n23452));
    SB_CARRY mod_5_add_1942_11 (.CI(n24128), .I0(n2801), .I1(n2819), .CO(n24129));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n24201), .O(n23_adj_4614)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n24127), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n24058), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n23888), .I0(n1608), .I1(n1631), .CO(n23889));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n23450), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n31924), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_7 (.CI(n24058), .I0(n2505), .I1(n2522), .CO(n24059));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n24057), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n24057), .I0(n2506), .I1(n2522), .CO(n24058));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n31936), 
            .I3(n23887), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n23887), .I0(n1609), .I1(n31936), .CO(n23888));
    SB_CARRY mod_5_add_1942_10 (.CI(n24127), .I0(n2802), .I1(n2819), .CO(n24128));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n31936), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n24056), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n31936), 
            .CO(n23887));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n23886), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n23885), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n24126), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n24201), .I0(n3103), .I1(n3116), .CO(n24202));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n24200), .O(n21_adj_4616)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n24056), .I0(n2507), .I1(n2522), .CO(n24057));
    SB_CARRY mod_5_add_1942_9 (.CI(n24126), .I0(n2803), .I1(n2819), .CO(n24127));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n24055), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1546 (.I0(n1499), .I1(n1504), .I2(n1503), .I3(n1505), 
            .O(n18_adj_4698));
    defparam i7_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1547 (.I0(bit_ctr[20]), .I1(n1508), .I2(n1509), 
            .I3(n1507), .O(n17_adj_4699));
    defparam i6_4_lut_adj_1547.LUT_INIT = 16'hffec;
    SB_LUT4 i8_4_lut_adj_1548 (.I0(n1502), .I1(n1506), .I2(n1501), .I3(n1500), 
            .O(n19_adj_4700));
    defparam i8_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_3_lut (.I0(n19_adj_4700), .I1(n17_adj_4699), .I2(n18_adj_4698), 
            .I3(GND_net), .O(n1532));
    defparam i10_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i26101_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31932));
    defparam i26101_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26102_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31933));
    defparam i26102_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n24125), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n24125), .I0(n2804), .I1(n2819), .CO(n24126));
    SB_CARRY mod_5_add_1741_4 (.CI(n24055), .I0(n2508), .I1(n2522), .CO(n24056));
    SB_CARRY mod_5_add_1205_14 (.CI(n23885), .I0(n1698), .I1(n1730), .CO(n23886));
    SB_CARRY mod_5_add_2143_8 (.CI(n24200), .I0(n3104), .I1(n3116), .CO(n24201));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n31931), 
            .I3(n24054), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n24199), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n23884), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n23884), .I0(n1699), .I1(n1730), .CO(n23885));
    SB_CARRY mod_5_add_2143_7 (.CI(n24199), .I0(n3105), .I1(n3116), .CO(n24200));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n23883), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n15508), 
            .D(n255[20]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1191__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n24198), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_3 (.CI(n24054), .I0(n2509), .I1(n31931), .CO(n24055));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n24124), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n31931), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_12 (.CI(n23883), .I0(n1700), .I1(n1730), .CO(n23884));
    SB_CARRY mod_5_add_1942_7 (.CI(n24124), .I0(n2805), .I1(n2819), .CO(n24125));
    SB_CARRY mod_5_add_2143_6 (.CI(n24198), .I0(n3106), .I1(n3116), .CO(n24199));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n24123), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n31931), 
            .CO(n24054));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n24053), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n23882), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n24052), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n24197), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n23438), .I0(n2306), .I1(n2324), .CO(n23439));
    SB_CARRY mod_5_add_1205_11 (.CI(n23882), .I0(n1701), .I1(n1730), .CO(n23883));
    SB_CARRY mod_5_add_2143_5 (.CI(n24197), .I0(n3107), .I1(n3116), .CO(n24198));
    SB_CARRY mod_5_add_1942_6 (.CI(n24123), .I0(n2806), .I1(n2819), .CO(n24124));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n23881), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n24196), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n24196), .I0(n3108), .I1(n3116), .CO(n24197));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n31921), 
            .I3(n24195), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n24122), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n23881), .I0(n1702), .I1(n1730), .CO(n23882));
    SB_CARRY mod_5_add_1942_5 (.CI(n24122), .I0(n2807), .I1(n2819), .CO(n24123));
    SB_CARRY mod_5_add_1674_21 (.CI(n24052), .I0(n2391), .I1(n2423), .CO(n24053));
    SB_CARRY mod_5_add_1607_18 (.CI(n23450), .I0(n2294), .I1(n2324), .CO(n23451));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n23449), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n24121), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_3 (.CI(n24195), .I0(n3109), .I1(n31921), .CO(n24196));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n31921), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n24051), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n31921), 
            .CO(n24195));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n23880), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n24194), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n24121), .I0(n2808), .I1(n2819), .CO(n24122));
    SB_CARRY mod_5_add_1674_20 (.CI(n24051), .I0(n2392), .I1(n2423), .CO(n24052));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n31930), 
            .I3(n24120), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n24120), .I0(n2809), .I1(n31930), .CO(n24121));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n31930), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n31930), 
            .CO(n24120));
    SB_CARRY mod_5_add_1205_9 (.CI(n23880), .I0(n1703), .I1(n1730), .CO(n23881));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n24193), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n24050), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n24119), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n24050), .I0(n2393), .I1(n2423), .CO(n24051));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n24049), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n23879), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n23879), .I0(n1704), .I1(n1730), .CO(n23880));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n23878), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n24193), .I0(n2985), .I1(n3017), .CO(n24194));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n24192), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n24192), .I0(n2986), .I1(n3017), .CO(n24193));
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n24118), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n24049), .I0(n2394), .I1(n2423), .CO(n24050));
    SB_CARRY mod_5_add_1875_24 (.CI(n24118), .I0(n2688), .I1(n2720), .CO(n24119));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n24191), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1549 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4701));
    defparam i15_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n24117), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n24048), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n24191), .I0(n2987), .I1(n3017), .CO(n24192));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n24190), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n24190), .I0(n2988), .I1(n3017), .CO(n24191));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n24189), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i21_4_lut_adj_1550 (.I0(n37_adj_4701), .I1(n39_adj_4697), .I2(n38_adj_4694), 
            .I3(n40_adj_4671), .O(n2621));
    defparam i21_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_23 (.CI(n24189), .I0(n2989), .I1(n3017), .CO(n24190));
    SB_LUT4 i3_4_lut_4_lut (.I0(n28587), .I1(n12895), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_CARRY mod_5_add_1674_17 (.CI(n24048), .I0(n2395), .I1(n2423), .CO(n24049));
    SB_CARRY mod_5_add_1875_23 (.CI(n24117), .I0(n2689), .I1(n2720), .CO(n24118));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n24188), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n24047), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n24047), .I0(n2396), .I1(n2423), .CO(n24048));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n24046), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n23878), .I0(n1705), .I1(n1730), .CO(n23879));
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4702));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_2076_22 (.CI(n24188), .I0(n2990), .I1(n3017), .CO(n24189));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n24187), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1551 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_4703));
    defparam i16_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i26006_3_lut_4_lut (.I0(n12895), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n28587), .O(n28613));   // verilog/neopixel.v(22[26:36])
    defparam i26006_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n15508), 
            .D(n255[19]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2076_21 (.CI(n24187), .I0(n2991), .I1(n3017), .CO(n24188));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n24186), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n24116), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n24116), .I0(n2690), .I1(n2720), .CO(n24117));
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_4704));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1552 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43_adj_4705));
    defparam i18_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1553 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_4706));
    defparam i15_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1554 (.I0(n41_adj_4703), .I1(n33_adj_4702), .I2(n2889), 
            .I3(n2901), .O(n46));
    defparam i21_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_15 (.CI(n24046), .I0(n2397), .I1(n2423), .CO(n24047));
    SB_CARRY mod_5_add_2076_20 (.CI(n24186), .I0(n2992), .I1(n3017), .CO(n24187));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n24185), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1555 (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39_adj_4707));
    defparam i14_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n24115), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i22_4_lut_adj_1556 (.I0(n43_adj_4705), .I1(n2904), .I2(n38_adj_4704), 
            .I3(n2893), .O(n47_adj_4708));
    defparam i22_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_4708), .I1(n39_adj_4707), .I2(n46), 
            .I3(n40_adj_4706), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1557 (.I0(bit_ctr[6]), .I1(bit_ctr[15]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[9]), .O(n18_adj_4709));
    defparam i7_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_21 (.CI(n24115), .I0(n2691), .I1(n2720), .CO(n24116));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n24045), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_4_lut_adj_1558 (.I0(bit_ctr[18]), .I1(n18_adj_4709), .I2(bit_ctr[13]), 
            .I3(bit_ctr[11]), .O(n20_adj_4710));
    defparam i9_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1559 (.I0(bit_ctr[8]), .I1(bit_ctr[10]), .I2(bit_ctr[27]), 
            .I3(bit_ctr[26]), .O(n19_adj_4711));
    defparam i8_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_19 (.CI(n24185), .I0(n2993), .I1(n3017), .CO(n24186));
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4712));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1560 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4713));
    defparam i13_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i15214_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n19755));
    defparam i15214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1561 (.I0(n1405), .I1(n19755), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4714));
    defparam i6_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1562 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4715));
    defparam i7_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1563 (.I0(n17_adj_4715), .I1(n1408), .I2(n16_adj_4714), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i26093_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31924));
    defparam i26093_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1564 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4716));
    defparam i1_3_lut_adj_1564.LUT_INIT = 16'hecec;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4717));
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'heeee;
    SB_LUT4 i15224_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n19765));
    defparam i15224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1566 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_4717), 
            .O(n30_adj_4718));
    defparam i13_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1567 (.I0(n2098), .I1(n19765), .I2(n2094), .I3(n2099), 
            .O(n28_adj_4719));
    defparam i11_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1568 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4720));
    defparam i12_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1569 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4721));
    defparam i10_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1570 (.I0(n27_adj_4721), .I1(n29_adj_4720), .I2(n28_adj_4719), 
            .I3(n30_adj_4718), .O(n2126));
    defparam i16_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1571 (.I0(n2490), .I1(n34_adj_4713), .I2(n24_adj_4712), 
            .I3(n2494), .O(n38_adj_4722));
    defparam i17_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1572 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4723));
    defparam i15_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1573 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4716), 
            .O(n37_adj_4724));
    defparam i16_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1574 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4725));
    defparam i14_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1575 (.I0(n35_adj_4725), .I1(n37_adj_4724), .I2(n36_adj_4723), 
            .I3(n38_adj_4722), .O(n2522));
    defparam i20_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 i26098_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31929));
    defparam i26098_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4726));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26097_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31928));
    defparam i26097_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1576 (.I0(bit_ctr[3]), .I1(n19_adj_4711), .I2(bit_ctr[4]), 
            .I3(n20_adj_4710), .O(n19_adj_4727));
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'hffec;
    SB_LUT4 i14_4_lut_adj_1577 (.I0(bit_ctr[20]), .I1(n19_adj_4727), .I2(bit_ctr[24]), 
            .I3(n20_adj_4726), .O(n32_adj_4728));
    defparam i14_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1578 (.I0(bit_ctr[23]), .I1(bit_ctr[5]), .I2(bit_ctr[29]), 
            .I3(bit_ctr[25]), .O(n30_adj_4729));
    defparam i12_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1579 (.I0(bit_ctr[30]), .I1(bit_ctr[7]), .I2(bit_ctr[14]), 
            .I3(bit_ctr[16]), .O(n31_adj_4730));
    defparam i13_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1580 (.I0(bit_ctr[28]), .I1(bit_ctr[31]), .I2(bit_ctr[21]), 
            .I3(bit_ctr[12]), .O(n29_adj_4731));
    defparam i11_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n32233));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n32233_bdd_4_lut (.I0(n32233), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n30363));
    defparam n32233_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i17_4_lut_adj_1581 (.I0(n29_adj_4731), .I1(n31_adj_4730), .I2(n30_adj_4729), 
            .I3(n32_adj_4728), .O(\state_3__N_372[1] ));
    defparam i17_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1582 (.I0(one_wire_N_523[3]), .I1(one_wire_N_523[4]), 
            .I2(one_wire_N_523[2]), .I3(GND_net), .O(n24851));
    defparam i2_3_lut_adj_1582.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1583 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n14300));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_2_lut_adj_1583.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_3_lut_adj_1584 (.I0(n24931), .I1(one_wire_N_523[4]), .I2(one_wire_N_523[3]), 
            .I3(GND_net), .O(n28657));
    defparam i1_3_lut_adj_1584.LUT_INIT = 16'hecec;
    SB_LUT4 i6_4_lut_adj_1585 (.I0(n14323), .I1(one_wire_N_523[5]), .I2(one_wire_N_523[10]), 
            .I3(one_wire_N_523[7]), .O(n14_adj_4732));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1586 (.I0(n9_adj_4695), .I1(n14_adj_4732), .I2(one_wire_N_523[8]), 
            .I3(one_wire_N_523[11]), .O(n14186));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i219_2_lut (.I0(LED_c), .I1(\state_3__N_372[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1121));   // verilog/neopixel.v(40[18] 45[12])
    defparam i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_1587 (.I0(n14186), .I1(n28657), .I2(GND_net), 
            .I3(GND_net), .O(n19684));
    defparam i2_2_lut_adj_1587.LUT_INIT = 16'heeee;
    SB_LUT4 i1633_4_lut (.I0(n19684), .I1(n1121), .I2(\state[1] ), .I3(n14300), 
            .O(n4607));
    defparam i1633_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 bit_ctr_0__bdd_4_lut_26351 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n32173));
    defparam bit_ctr_0__bdd_4_lut_26351.LUT_INIT = 16'he4aa;
    SB_LUT4 n32173_bdd_4_lut (.I0(n32173), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n30471));
    defparam n32173_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_26301 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n32167));
    defparam bit_ctr_0__bdd_4_lut_26301.LUT_INIT = 16'he4aa;
    SB_LUT4 n32167_bdd_4_lut (.I0(n32167), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n30474));
    defparam n32167_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_26296 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n32119));
    defparam bit_ctr_0__bdd_4_lut_26296.LUT_INIT = 16'he4aa;
    SB_LUT4 n32119_bdd_4_lut (.I0(n32119), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n32122));
    defparam n32119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n30471), .I2(n30474), 
            .I3(n25270), .O(n32095));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n32095_bdd_4_lut (.I0(n32095), .I1(n31960), .I2(n30363), .I3(n25270), 
            .O(n32098));
    defparam n32095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_26257 (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n32017));
    defparam bit_ctr_0__bdd_4_lut_26257.LUT_INIT = 16'he4aa;
    SB_LUT4 n32017_bdd_4_lut (.I0(n32017), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n32020));
    defparam n32017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n24114), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i26025_4_lut (.I0(\state[1] ), .I1(n31156), .I2(state[0]), 
            .I3(n4607), .O(n15508));
    defparam i26025_4_lut.LUT_INIT = 16'h01f1;
    SB_LUT4 i16_4_lut_adj_1588 (.I0(n21_adj_4672), .I1(n23_adj_4665), .I2(n22_adj_4661), 
            .I3(n24_adj_4684), .O(n36_adj_4733));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1589 (.I0(n25_adj_4685), .I1(n27_adj_4659), .I2(n26_adj_4669), 
            .I3(n28_adj_4668), .O(n37_adj_4734));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1590 (.I0(n37_adj_4734), .I1(n29_adj_4675), .I2(n36_adj_4733), 
            .I3(n30_adj_4676), .O(n14323));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i22834_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n28653));
    defparam i22834_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26005_2_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n27865));
    defparam i26005_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1591 (.I0(one_wire_N_523[4]), .I1(one_wire_N_523[3]), 
            .I2(n27865), .I3(n24931), .O(n111));
    defparam i1_4_lut_adj_1591.LUT_INIT = 16'h5155;
    SB_LUT4 i1_4_lut_adj_1592 (.I0(n111), .I1(n27865), .I2(one_wire_N_523[2]), 
            .I3(one_wire_N_523[3]), .O(n116));
    defparam i1_4_lut_adj_1592.LUT_INIT = 16'haeee;
    SB_LUT4 i6_4_lut_adj_1593 (.I0(one_wire_N_523[8]), .I1(one_wire_N_523[10]), 
            .I2(n28653), .I3(n116), .O(n16_adj_4735));
    defparam i6_4_lut_adj_1593.LUT_INIT = 16'h0100;
    SB_LUT4 i8_3_lut_adj_1594 (.I0(one_wire_N_523[5]), .I1(n16_adj_4735), 
            .I2(n14323), .I3(GND_net), .O(n18_adj_4736));
    defparam i8_3_lut_adj_1594.LUT_INIT = 16'h0404;
    SB_LUT4 i3_4_lut_adj_1595 (.I0(n9_adj_4695), .I1(one_wire_N_523[11]), 
            .I2(n18_adj_4736), .I3(one_wire_N_523[7]), .O(n32240));
    defparam i3_4_lut_adj_1595.LUT_INIT = 16'hffef;
    SB_LUT4 i25573_3_lut_4_lut (.I0(n24851), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n14186), .O(n31156));
    defparam i25573_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_372[1] ), .O(n15621));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY mod_5_add_1674_14 (.CI(n24045), .I0(n2398), .I1(n2423), .CO(n24046));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n23877), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n23877), .I0(n1706), .I1(n1730), .CO(n23878));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n24184), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n24044), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n19721), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[29]), .O(n25284));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ba;
    SB_LUT4 mod_5_i471_3_lut_4_lut_4_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(bit_ctr[29]), .I3(n19721), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'hd262;
    SB_LUT4 i3380_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n28587), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i3380_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n23974), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n24114), .I0(n2692), .I1(n2720), .CO(n24115));
    SB_CARRY mod_5_add_2076_18 (.CI(n24184), .I0(n2994), .I1(n3017), .CO(n24185));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n24113), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n24044), .I0(n2399), .I1(n2423), .CO(n24045));
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n23973), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n23876), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n24183), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n24113), .I0(n2693), .I1(n2720), .CO(n24114));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n24043), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n23973), .I0(n1104), .I1(n1136), .CO(n23974));
    SB_CARRY mod_5_add_1674_12 (.CI(n24043), .I0(n2400), .I1(n2423), .CO(n24044));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n24112), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n24112), .I0(n2694), .I1(n2720), .CO(n24113));
    SB_CARRY mod_5_add_2076_17 (.CI(n24183), .I0(n2995), .I1(n3017), .CO(n24184));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n24182), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n24182), .I0(n2996), .I1(n3017), .CO(n24183));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n24181), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n23876), .I0(n1707), .I1(n1730), .CO(n23877));
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n15508), 
            .D(n255[18]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n24111), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n24042), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n23972), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n24042), .I0(n2401), .I1(n2423), .CO(n24043));
    SB_CARRY mod_5_add_2076_15 (.CI(n24181), .I0(n2997), .I1(n3017), .CO(n24182));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n23875), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n24111), .I0(n2695), .I1(n2720), .CO(n24112));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n24041), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n24180), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n24180), .I0(n2998), .I1(n3017), .CO(n24181));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n24110), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n24041), .I0(n2402), .I1(n2423), .CO(n24042));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n24179), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n24110), .I0(n2696), .I1(n2720), .CO(n24111));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n24109), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n24109), .I0(n2697), .I1(n2720), .CO(n24110));
    SB_CARRY mod_5_add_2076_13 (.CI(n24179), .I0(n2999), .I1(n3017), .CO(n24180));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n24108), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n24108), .I0(n2698), .I1(n2720), .CO(n24109));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n24107), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n24178), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n24178), .I0(n3000), .I1(n3017), .CO(n24179));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n24040), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n24177), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk32MHz), .E(n15451), .D(state_3__N_372[0]), 
            .S(n28597));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_9 (.CI(n24040), .I0(n2403), .I1(n2423), .CO(n24041));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n24039), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n24107), .I0(n2699), .I1(n2720), .CO(n24108));
    SB_CARRY mod_5_add_1674_8 (.CI(n24039), .I0(n2404), .I1(n2423), .CO(n24040));
    SB_CARRY mod_5_add_803_7 (.CI(n23972), .I0(n1105), .I1(n1136), .CO(n23973));
    SB_CARRY mod_5_add_1205_4 (.CI(n23875), .I0(n1708), .I1(n1730), .CO(n23876));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n24038), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n24177), .I0(n3001), .I1(n3017), .CO(n24178));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n24176), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n24106), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n24106), .I0(n2700), .I1(n2720), .CO(n24107));
    SB_CARRY mod_5_add_1674_7 (.CI(n24038), .I0(n2405), .I1(n2423), .CO(n24039));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n23971), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n31937), 
            .I3(n23874), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_17 (.CI(n23449), .I0(n2295), .I1(n2324), .CO(n23450));
    SB_CARRY mod_5_add_2076_10 (.CI(n24176), .I0(n3002), .I1(n3017), .CO(n24177));
    SB_CARRY mod_5_add_803_6 (.CI(n23971), .I0(n1106), .I1(n1136), .CO(n23972));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n23970), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_3 (.CI(n23874), .I0(n1709), .I1(n31937), .CO(n23875));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n24175), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n24105), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n24105), .I0(n2701), .I1(n2720), .CO(n24106));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n24037), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n23970), .I0(n1107), .I1(n1136), .CO(n23971));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n31937), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_24 (.CI(n23475), .I0(bit_ctr[22]), .I1(GND_net), .CO(n23476));
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n15508), 
            .D(n255[6]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2076_9 (.CI(n24175), .I0(n3003), .I1(n3017), .CO(n24176));
    SB_CARRY mod_5_add_1674_6 (.CI(n24037), .I0(n2406), .I1(n2423), .CO(n24038));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n24104), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n15508), 
            .D(n255[5]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n15508), 
            .D(n255[17]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n15508), 
            .D(n255[16]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n15508), 
            .D(n255[4]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i22822_2_lut_4_lut (.I0(bit_ctr[28]), .I1(n19721), .I2(n608), 
            .I3(bit_ctr[29]), .O(n28641));
    defparam i22822_2_lut_4_lut.LUT_INIT = 16'h02a8;
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n24036), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15181_2_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n19721));
    defparam i15181_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mux_635_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_580 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_635_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n15508), 
            .D(n255[3]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n15508), 
            .D(n255[15]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n28787), .D(\neo_pixel_transmitter.done_N_586 ), 
            .R(n30218));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n24174), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n24174), .I0(n3004), .I1(n3017), .CO(n24175));
    SB_CARRY mod_5_add_1875_10 (.CI(n24104), .I0(n2702), .I1(n2720), .CO(n24105));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n23969), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n24036), .I0(n2407), .I1(n2423), .CO(n24037));
    SB_CARRY mod_5_add_803_4 (.CI(n23969), .I0(n1108), .I1(n1136), .CO(n23970));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n24173), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n31937), 
            .CO(n23874));
    SB_CARRY mod_5_add_2076_7 (.CI(n24173), .I0(n3005), .I1(n3017), .CO(n24174));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n24172), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n24103), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n24103), .I0(n2703), .I1(n2720), .CO(n24104));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n24035), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n24035), .I0(n2408), .I1(n2423), .CO(n24036));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n31941), 
            .I3(n23968), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n23873), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n23872), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n31938), 
            .I3(n24034), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_6 (.CI(n24172), .I0(n3006), .I1(n3017), .CO(n24173));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n24102), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_3 (.CI(n24034), .I0(n2409), .I1(n31938), .CO(n24035));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n24171), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n24102), .I0(n2704), .I1(n2720), .CO(n24103));
    SB_CARRY mod_5_add_2076_5 (.CI(n24171), .I0(n3007), .I1(n3017), .CO(n24172));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n24101), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n23872), .I0(n1797), .I1(n1829), .CO(n23873));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n23871), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n24101), .I0(n2705), .I1(n2720), .CO(n24102));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n31938), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n23968), .I0(n1109), .I1(n31941), .CO(n23969));
    SB_CARRY mod_5_add_1272_14 (.CI(n23871), .I0(n1798), .I1(n1829), .CO(n23872));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n31941), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n24170), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n24170), .I0(n3008), .I1(n3017), .CO(n24171));
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n31941), 
            .CO(n23968));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n24100), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n24100), .I0(n2706), .I1(n2720), .CO(n24101));
    SB_LUT4 timer_1191_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n23967), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n23870), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n15761));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i25678_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n15566));
    defparam i25678_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_CARRY mod_5_add_1272_13 (.CI(n23870), .I0(n1799), .I1(n1829), .CO(n23871));
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n15760));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n15759));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n15758));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n15757));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n15756));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n15755));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n15754));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n15753));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n15752));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n15751));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n15750));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n15749));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n15748));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n15747));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n15746));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n15745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n15744));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n15743));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n15742));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n15741));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n15740));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n15739));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n15738));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n15737));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n15736));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n15735));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n15734));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n15733));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n15732));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n15731));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n15508), 
            .D(n255[2]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 bit_ctr_0__bdd_4_lut_26174 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n31957));
    defparam bit_ctr_0__bdd_4_lut_26174.LUT_INIT = 16'he4aa;
    SB_LUT4 n31957_bdd_4_lut (.I0(n31957), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n31960));
    defparam n31957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n15508), 
            .D(n255[14]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n24099), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1596 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4737));
    defparam i16_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n31939), 
            .I3(n24169), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n24169), .I0(n3009), .I1(n31939), .CO(n24170));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n31939), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_5 (.CI(n24099), .I0(n2707), .I1(n2720), .CO(n24100));
    SB_LUT4 i14_4_lut_adj_1597 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4738));
    defparam i14_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut_adj_1598 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4739));
    defparam i3_2_lut_adj_1598.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1599 (.I0(bit_ctr[12]), .I1(n22_adj_4739), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4740));
    defparam i11_4_lut_adj_1599.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1600 (.I0(n2294), .I1(n30_adj_4740), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4741));
    defparam i15_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1601 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4742));
    defparam i13_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1602 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4743));
    defparam i14_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1603 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4744));
    defparam i12_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1604 (.I0(n31_adj_4744), .I1(n33_adj_4743), .I2(n32_adj_4742), 
            .I3(n34_adj_4741), .O(n2324));
    defparam i18_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1605 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42_adj_4745));
    defparam i15_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1606 (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46_adj_4746));
    defparam i19_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1607 (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44_adj_4747));
    defparam i17_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1608 (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45_adj_4748));
    defparam i18_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1609 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43_adj_4749));
    defparam i16_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut_adj_1610 (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), 
            .I3(GND_net), .O(n40_adj_4750));
    defparam i13_3_lut_adj_1610.LUT_INIT = 16'hecec;
    SB_LUT4 i21_4_lut_adj_1611 (.I0(n3107), .I1(n42_adj_4745), .I2(n3087), 
            .I3(n3086), .O(n48));
    defparam i21_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1612 (.I0(n43_adj_4749), .I1(n45_adj_4748), .I2(n44_adj_4747), 
            .I3(n46_adj_4746), .O(n52));
    defparam i25_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3095), .I1(n3084), .I2(GND_net), .I3(GND_net), 
            .O(n39_adj_4751));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26_4_lut (.I0(n39_adj_4751), .I1(n52), .I2(n48), .I3(n40_adj_4750), 
            .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n23484), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n23448), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n26505));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n31938), 
            .CO(n24034));
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n23483), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_32 (.CI(n23483), .I0(bit_ctr[30]), .I1(GND_net), .CO(n23484));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n31939), 
            .CO(n24169));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n24098), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n23966), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n23482), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n24168), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n23869), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n24098), .I0(n2708), .I1(n2720), .CO(n24099));
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n24167), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1191__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i15_4_lut_adj_1613 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4752));
    defparam i15_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n24033), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1191_add_4_32 (.CI(n23966), .I0(GND_net), .I1(timer[30]), 
            .CO(n23967));
    SB_CARRY mod_5_add_1272_12 (.CI(n23869), .I0(n1800), .I1(n1829), .CO(n23870));
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n24032), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n23868), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n31940), 
            .I3(n24097), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i13_4_lut_adj_1614 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4753));
    defparam i13_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_26 (.CI(n24167), .I0(n2886), .I1(n2918), .CO(n24168));
    SB_CARRY mod_5_add_669_6 (.CI(n24032), .I0(n906), .I1(VCC_net), .CO(n24033));
    SB_CARRY add_21_31 (.CI(n23482), .I0(bit_ctr[29]), .I1(GND_net), .CO(n23483));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n23481), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1191_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n23965), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n24166), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4754));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n15508), 
            .D(n255[13]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i18_4_lut_adj_1615 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4755));
    defparam i18_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n15508), 
            .D(n255[12]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n15508), 
            .D(n255[11]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n15508), 
            .D(n255[10]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2009_25 (.CI(n24166), .I0(n2887), .I1(n2918), .CO(n24167));
    SB_CARRY add_21_30 (.CI(n23481), .I0(bit_ctr[28]), .I1(GND_net), .CO(n23482));
    SB_CARRY mod_5_add_1875_3 (.CI(n24097), .I0(n2709), .I1(n31940), .CO(n24098));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n24165), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n31940), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n28613), .I2(VCC_net), 
            .I3(n24031), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n24031), .I0(n28613), .I1(VCC_net), 
            .CO(n24032));
    SB_CARRY timer_1191_add_4_31 (.CI(n23965), .I0(GND_net), .I1(timer[29]), 
            .CO(n23966));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n23480), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_11 (.CI(n23868), .I0(n1801), .I1(n1829), .CO(n23869));
    SB_LUT4 i22_4_lut_adj_1616 (.I0(n37_adj_4753), .I1(n39_adj_4752), .I2(n38_adj_4738), 
            .I3(n40_adj_4737), .O(n46_adj_4756));
    defparam i22_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1191_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n23964), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_16 (.CI(n23448), .I0(n2296), .I1(n2324), .CO(n23449));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n23867), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n31940), 
            .CO(n24097));
    SB_LUT4 i2_3_lut_adj_1617 (.I0(n19831), .I1(state[0]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n29426));   // verilog/neopixel.v(36[4] 116[11])
    defparam i2_3_lut_adj_1617.LUT_INIT = 16'hfdfd;
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n15566), .I2(VCC_net), 
            .I3(n24030), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_24 (.CI(n24165), .I0(n2888), .I1(n2918), .CO(n24166));
    SB_CARRY timer_1191_add_4_30 (.CI(n23964), .I0(GND_net), .I1(timer[28]), 
            .CO(n23965));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n24096), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_4 (.CI(n24030), .I0(n15566), .I1(VCC_net), 
            .CO(n24031));
    SB_LUT4 timer_1191_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n23963), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n24095), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n23867), .I0(n1802), .I1(n1829), .CO(n23868));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n23866), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4757));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n24164), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_29 (.CI(n23963), .I0(GND_net), .I1(timer[27]), 
            .CO(n23964));
    SB_CARRY mod_5_add_1808_23 (.CI(n24095), .I0(n2589), .I1(n2621), .CO(n24096));
    SB_CARRY add_21_29 (.CI(n23480), .I0(bit_ctr[27]), .I1(GND_net), .CO(n23481));
    SB_LUT4 i1_2_lut_3_lut (.I0(n28731), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n12074));   // verilog/neopixel.v(36[4] 116[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n24094), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n24094), .I0(n2590), .I1(n2621), .CO(n24095));
    SB_LUT4 timer_1191_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n23962), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n15508), 
            .D(n255[9]), .R(n15621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n24093), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n24164), .I0(n2889), .I1(n2918), .CO(n24165));
    SB_DFF timer_1191__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n12921), .I2(GND_net), 
            .I3(n24029), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1191_add_4_28 (.CI(n23962), .I0(GND_net), .I1(timer[26]), 
            .CO(n23963));
    SB_CARRY mod_5_add_1808_21 (.CI(n24093), .I0(n2591), .I1(n2621), .CO(n24094));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n24163), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_3 (.CI(n24029), .I0(n12921), .I1(GND_net), 
            .CO(n24030));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n24092), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n23866), .I0(n1803), .I1(n1829), .CO(n23867));
    SB_LUT4 i25576_3_lut_4_lut (.I0(n14186), .I1(n31408), .I2(start), 
            .I3(\state[1] ), .O(n31409));
    defparam i25576_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_22 (.CI(n24163), .I0(n2890), .I1(n2918), .CO(n24164));
    SB_LUT4 timer_1191_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n23961), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n24162), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_27 (.CI(n23961), .I0(GND_net), .I1(timer[25]), 
            .CO(n23962));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n23865), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_4_lut_4_lut_adj_1618 (.I0(n19831), .I1(\state[1] ), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n30218));
    defparam i3_4_lut_4_lut_adj_1618.LUT_INIT = 16'h0004;
    SB_CARRY mod_5_add_1808_20 (.CI(n24092), .I0(n2592), .I1(n2621), .CO(n24093));
    SB_CARRY mod_5_add_2009_21 (.CI(n24162), .I0(n2891), .I1(n2918), .CO(n24163));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n24161), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n24161), .I0(n2892), .I1(n2918), .CO(n24162));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n24160), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1191_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n23960), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_8 (.CI(n23865), .I0(n1804), .I1(n1829), .CO(n23866));
    SB_DFF timer_1191__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1191__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i23_4_lut_adj_1619 (.I0(n33_adj_4757), .I1(n46_adj_4756), .I2(n42_adj_4755), 
            .I3(n34_adj_4754), .O(n2819));
    defparam i23_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n15726));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n15704));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n24029));
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n23479), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_19 (.CI(n24160), .I0(n2893), .I1(n2918), .CO(n24161));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n24159), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4), .I1(n4), .I2(n1037), .I3(n24028), 
            .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n24091), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_26 (.CI(n23960), .I0(GND_net), .I1(timer[24]), 
            .CO(n23961));
    SB_CARRY mod_5_add_1808_19 (.CI(n24091), .I0(n2593), .I1(n2621), .CO(n24092));
    SB_CARRY mod_5_add_2009_18 (.CI(n24159), .I0(n2894), .I1(n2918), .CO(n24160));
    SB_LUT4 timer_1191_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n23959), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1191_add_4_25 (.CI(n23959), .I0(GND_net), .I1(timer[23]), 
            .CO(n23960));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n24158), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n24090), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n24027), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n24158), .I0(n2895), .I1(n2918), .CO(n24159));
    SB_CARRY mod_5_add_736_7 (.CI(n24027), .I0(n1005), .I1(n1037), .CO(n24028));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n24157), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_2_lut_adj_1620 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4655));
    defparam i2_2_lut_adj_1620.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1621 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4683));
    defparam i12_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_16 (.CI(n24157), .I0(n2896), .I1(n2918), .CO(n24158));
    SB_LUT4 timer_1191_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n23958), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n24156), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n24090), .I0(n2594), .I1(n2621), .CO(n24091));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n24026), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n24089), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_24 (.CI(n23958), .I0(GND_net), .I1(timer[22]), 
            .CO(n23959));
    SB_CARRY mod_5_add_2009_15 (.CI(n24156), .I0(n2897), .I1(n2918), .CO(n24157));
    SB_CARRY mod_5_add_1808_17 (.CI(n24089), .I0(n2595), .I1(n2621), .CO(n24090));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n24088), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n24155), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n24026), .I0(n1006), .I1(n1037), .CO(n24027));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n24025), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n24155), .I0(n2898), .I1(n2918), .CO(n24156));
    SB_LUT4 timer_1191_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n23957), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n23864), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n23447), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n24154), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_23 (.CI(n23957), .I0(GND_net), .I1(timer[21]), 
            .CO(n23958));
    SB_CARRY mod_5_add_2009_13 (.CI(n24154), .I0(n2899), .I1(n2918), .CO(n24155));
    SB_CARRY mod_5_add_1272_7 (.CI(n23864), .I0(n1805), .I1(n1829), .CO(n23865));
    SB_CARRY mod_5_add_736_5 (.CI(n24025), .I0(n1007), .I1(n1037), .CO(n24026));
    SB_CARRY mod_5_add_1808_16 (.CI(n24088), .I0(n2596), .I1(n2621), .CO(n24089));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n24024), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_28 (.CI(n23479), .I0(bit_ctr[26]), .I1(GND_net), .CO(n23480));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n24221), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n24220), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n24220), .I0(n3084), .I1(n3116), .CO(n24221));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n23478), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1191_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n23956), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_15 (.CI(n23447), .I0(n2297), .I1(n2324), .CO(n23448));
    SB_CARRY add_21_27 (.CI(n23478), .I0(bit_ctr[25]), .I1(GND_net), .CO(n23479));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n24219), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n31924), 
            .CO(n23435));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n24153), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n24087), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n24153), .I0(n2900), .I1(n2918), .CO(n24154));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n23863), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_22 (.CI(n23956), .I0(GND_net), .I1(timer[20]), 
            .CO(n23957));
    SB_LUT4 timer_1191_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n23955), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_27 (.CI(n24219), .I0(n3085), .I1(n3116), .CO(n24220));
    SB_CARRY mod_5_add_1272_6 (.CI(n23863), .I0(n1806), .I1(n1829), .CO(n23864));
    SB_CARRY mod_5_add_736_4 (.CI(n24024), .I0(n1008), .I1(n1037), .CO(n24025));
    SB_CARRY mod_5_add_1808_15 (.CI(n24087), .I0(n2597), .I1(n2621), .CO(n24088));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n24152), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n24152), .I0(n2901), .I1(n2918), .CO(n24153));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n31943), 
            .I3(n24023), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n24218), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n24086), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_3 (.CI(n24023), .I0(n1009), .I1(n31943), .CO(n24024));
    SB_CARRY mod_5_add_2143_26 (.CI(n24218), .I0(n3086), .I1(n3116), .CO(n24219));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n24151), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n24086), .I0(n2598), .I1(n2621), .CO(n24087));
    SB_CARRY mod_5_add_2009_10 (.CI(n24151), .I0(n2902), .I1(n2918), .CO(n24152));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n23477), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n31943), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n24217), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n24150), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n24085), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n31943), 
            .CO(n24023));
    SB_CARRY timer_1191_add_4_21 (.CI(n23955), .I0(GND_net), .I1(timer[19]), 
            .CO(n23956));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n23862), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n23862), .I0(n1807), .I1(n1829), .CO(n23863));
    SB_LUT4 i10_4_lut_adj_1622 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4682));
    defparam i10_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_26 (.CI(n23477), .I0(bit_ctr[24]), .I1(GND_net), .CO(n23478));
    SB_CARRY mod_5_add_2009_9 (.CI(n24150), .I0(n2903), .I1(n2918), .CO(n24151));
    SB_CARRY mod_5_add_1808_13 (.CI(n24085), .I0(n2599), .I1(n2621), .CO(n24086));
    SB_LUT4 timer_1191_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n23954), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n23861), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n24217), .I0(n3087), .I1(n3116), .CO(n24218));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n24149), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n24084), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n24216), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1191_add_4_20 (.CI(n23954), .I0(GND_net), .I1(timer[18]), 
            .CO(n23955));
    SB_CARRY mod_5_add_1272_4 (.CI(n23861), .I0(n1808), .I1(n1829), .CO(n23862));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n31942), 
            .I3(n23860), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1191_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n23953), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_3 (.CI(n23860), .I0(n1809), .I1(n31942), .CO(n23861));
    SB_CARRY mod_5_add_2009_8 (.CI(n24149), .I0(n2904), .I1(n2918), .CO(n24150));
    SB_CARRY mod_5_add_1808_12 (.CI(n24084), .I0(n2600), .I1(n2621), .CO(n24085));
    SB_CARRY mod_5_add_2143_24 (.CI(n24216), .I0(n3088), .I1(n3116), .CO(n24217));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n23476), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n24148), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n24083), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n24215), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n24148), .I0(n2905), .I1(n2918), .CO(n24149));
    SB_CARRY mod_5_add_2143_23 (.CI(n24215), .I0(n3089), .I1(n3116), .CO(n24216));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n24147), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_25 (.CI(n23476), .I0(bit_ctr[23]), .I1(GND_net), .CO(n23477));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n31942), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n23475), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_22 (.CI(n23473), .I0(bit_ctr[20]), .I1(GND_net), .CO(n23474));
    SB_CARRY timer_1191_add_4_19 (.CI(n23953), .I0(GND_net), .I1(timer[17]), 
            .CO(n23954));
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n31942), 
            .CO(n23860));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n23474), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n23474), .I0(bit_ctr[21]), .I1(GND_net), .CO(n23475));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n23446), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n23446), .I0(n2298), .I1(n2324), .CO(n23447));
    SB_CARRY mod_5_add_1808_11 (.CI(n24083), .I0(n2601), .I1(n2621), .CO(n24084));
    SB_LUT4 timer_1191_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n23952), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1191_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1191_add_4_18 (.CI(n23952), .I0(GND_net), .I1(timer[16]), 
            .CO(n23953));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n24214), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i26108_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31939));
    defparam i26108_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, GND_net, clk32MHz, 
            data_o, reg_B, n29458, ENCODER1_A_c_1, ENCODER1_B_c_0, 
            n16239, n15723) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder1_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output [1:0]reg_B;
    output n29458;
    input ENCODER1_A_c_1;
    input ENCODER1_B_c_0;
    input n16239;
    input n15723;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2799;
    
    wire n2784, n23695, n23696, n23694, n23693, n23692, n23691, 
        n23690, n23689, n23688, n23687, n23686, n23685, n23684, 
        n23683, n23682, n23681, n23680, n23679, n23678, n23677, 
        count_direction, n23676, count_enable, B_delayed, A_delayed, 
        n23699, n23698, n23697;
    
    SB_LUT4 add_577_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2784), 
            .I3(n23695), .O(n2799[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_21 (.CI(n23695), .I0(encoder1_position[19]), .I1(n2784), 
            .CO(n23696));
    SB_LUT4 add_577_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2784), 
            .I3(n23694), .O(n2799[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_20 (.CI(n23694), .I0(encoder1_position[18]), .I1(n2784), 
            .CO(n23695));
    SB_LUT4 add_577_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2784), 
            .I3(n23693), .O(n2799[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_19 (.CI(n23693), .I0(encoder1_position[17]), .I1(n2784), 
            .CO(n23694));
    SB_LUT4 add_577_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2784), 
            .I3(n23692), .O(n2799[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_18 (.CI(n23692), .I0(encoder1_position[16]), .I1(n2784), 
            .CO(n23693));
    SB_LUT4 add_577_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2784), 
            .I3(n23691), .O(n2799[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_17 (.CI(n23691), .I0(encoder1_position[15]), .I1(n2784), 
            .CO(n23692));
    SB_LUT4 add_577_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2784), 
            .I3(n23690), .O(n2799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_16 (.CI(n23690), .I0(encoder1_position[14]), .I1(n2784), 
            .CO(n23691));
    SB_LUT4 add_577_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2784), 
            .I3(n23689), .O(n2799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_15 (.CI(n23689), .I0(encoder1_position[13]), .I1(n2784), 
            .CO(n23690));
    SB_LUT4 add_577_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2784), 
            .I3(n23688), .O(n2799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_14 (.CI(n23688), .I0(encoder1_position[12]), .I1(n2784), 
            .CO(n23689));
    SB_LUT4 add_577_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2784), 
            .I3(n23687), .O(n2799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_13 (.CI(n23687), .I0(encoder1_position[11]), .I1(n2784), 
            .CO(n23688));
    SB_LUT4 add_577_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2784), 
            .I3(n23686), .O(n2799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_12 (.CI(n23686), .I0(encoder1_position[10]), .I1(n2784), 
            .CO(n23687));
    SB_LUT4 add_577_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2784), 
            .I3(n23685), .O(n2799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_11 (.CI(n23685), .I0(encoder1_position[9]), .I1(n2784), 
            .CO(n23686));
    SB_LUT4 add_577_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2784), 
            .I3(n23684), .O(n2799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_10 (.CI(n23684), .I0(encoder1_position[8]), .I1(n2784), 
            .CO(n23685));
    SB_LUT4 add_577_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2784), 
            .I3(n23683), .O(n2799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_9 (.CI(n23683), .I0(encoder1_position[7]), .I1(n2784), 
            .CO(n23684));
    SB_LUT4 add_577_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2784), 
            .I3(n23682), .O(n2799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_8 (.CI(n23682), .I0(encoder1_position[6]), .I1(n2784), 
            .CO(n23683));
    SB_LUT4 add_577_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2784), 
            .I3(n23681), .O(n2799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_7 (.CI(n23681), .I0(encoder1_position[5]), .I1(n2784), 
            .CO(n23682));
    SB_LUT4 add_577_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2784), 
            .I3(n23680), .O(n2799[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_6 (.CI(n23680), .I0(encoder1_position[4]), .I1(n2784), 
            .CO(n23681));
    SB_LUT4 add_577_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2784), 
            .I3(n23679), .O(n2799[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_5 (.CI(n23679), .I0(encoder1_position[3]), .I1(n2784), 
            .CO(n23680));
    SB_LUT4 add_577_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2784), 
            .I3(n23678), .O(n2799[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_4 (.CI(n23678), .I0(encoder1_position[2]), .I1(n2784), 
            .CO(n23679));
    SB_LUT4 add_577_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2784), 
            .I3(n23677), .O(n2799[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_3 (.CI(n23677), .I0(encoder1_position[1]), .I1(n2784), 
            .CO(n23678));
    SB_LUT4 add_577_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n23676), .O(n2799[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_2 (.CI(n23676), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n23677));
    SB_CARRY add_577_1 (.CI(GND_net), .I0(n2784), .I1(n2784), .CO(n23676));
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i905_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2784));   // quad.v(37[5] 40[8])
    defparam i905_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2799[23]));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_577_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2784), 
            .I3(n23699), .O(n2799[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_577_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2784), 
            .I3(n23698), .O(n2799[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_24 (.CI(n23698), .I0(encoder1_position[22]), .I1(n2784), 
            .CO(n23699));
    SB_LUT4 add_577_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2784), 
            .I3(n23697), .O(n2799[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_23 (.CI(n23697), .I0(encoder1_position[21]), .I1(n2784), 
            .CO(n23698));
    SB_LUT4 add_577_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2784), 
            .I3(n23696), .O(n2799[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_22 (.CI(n23696), .I0(encoder1_position[20]), .I1(n2784), 
            .CO(n23697));
    \grp_debouncer(2,5)  debounce (.reg_B({reg_B}), .GND_net(GND_net), .n29458(n29458), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n16239(n16239), .data_o({data_o}), .n15723(n15723));   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (reg_B, GND_net, n29458, ENCODER1_A_c_1, 
            clk32MHz, ENCODER1_B_c_0, n16239, data_o, n15723);
    output [1:0]reg_B;
    input GND_net;
    output n29458;
    input ENCODER1_A_c_1;
    input clk32MHz;
    input ENCODER1_B_c_0;
    input n16239;
    output [1:0]data_o;
    input n15723;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3732;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n29458), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i18636_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i18636_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18645_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i18645_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i18638_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i18638_2_lut.LUT_INIT = 16'h6666;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1199__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n16239));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i2_3_lut_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n29458));
    defparam i2_3_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n15723));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1199__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1199__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3732));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (setpoint, GND_net, \Kp[12] , \Kp[13] , \Kp[14] , 
            \Kp[15] , \Ki[13] , \Kp[1] , \Kp[0] , \Kp[2] , \Kp[3] , 
            \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Ki[14] , \Ki[15] , \Ki[1] , \Ki[0] , 
            \Ki[2] , \Ki[3] , \Ki[4] , motor_state, \Ki[5] , \Ki[6] , 
            \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , VCC_net, \Ki[11] , 
            \Ki[12] , PWMLimit, IntegralLimit, duty, clk32MHz, n25, 
            n31935) /* synthesis syn_module_defined=1 */ ;
    input [23:0]setpoint;
    input GND_net;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Ki[13] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input [23:0]motor_state;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input VCC_net;
    input \Ki[11] ;
    input \Ki[12] ;
    input [23:0]PWMLimit;
    input [23:0]IntegralLimit;
    output [23:0]duty;
    input clk32MHz;
    input n25;
    output n31935;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(21[23:26])
    
    wire n898, n971, n1044, n1117;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n956, n98, n29, n171, n244, n317, n390, n463, n536, 
        n609, n682, n755, n828, n901, n1029, n83, n1102, n14, 
        n159, n974, n24280;
    wire [19:0]n7395;
    
    wire n24281, n1047, n1120, n156;
    wire [20:0]n7372;
    
    wire n24279, n101, n83_adj_4179, n14_adj_4180, n156_adj_4181, 
        n32, n229, n302, n174, n229_adj_4182;
    wire [23:0]\PID_CONTROLLER.err_23__N_3552 ;
    
    wire n23657, n23656, n23655, n23654, n23653, n375, n23652, 
        n23651, n23650, n448, n521, n247, n23649, n23648, n320, 
        n23647, n23646, n24351;
    wire [15:0]n7477;
    
    wire n1041, n24352, n594, n23645, n23644, n667;
    wire [23:0]n28;
    
    wire n24007, n23643, n23642, n24006, n23641, n23640, n23639, 
        n740, n23638, n232, n393, n24005, n23637, n466, n23636, 
        n539, n23635, n305, n813, n24004, n886;
    wire [23:0]duty_23__N_3651;
    wire [23:0]n2901;
    wire [23:0]n2926;
    
    wire n23634, n23633, n378, n959, n1032, n612, n1105, n23632, 
        n302_adj_4184, n375_adj_4185, n822, n895, n968, n1041_adj_4186, 
        n1114, n448_adj_4187, n86, n521_adj_4188, n95, n23631, n17_adj_4189, 
        n77, n26, n8_adj_4190, n168, n23630, n159_adj_4191;
    wire [16:0]n7458;
    
    wire n968_adj_4192, n24350, n685, n23629, n600, n1102_adj_4193, 
        n24278, n241, n314, n594_adj_4194, n387, n24003, n460, 
        n533, n606, n679, n758, n752, n825, n898_adj_4195, n971_adj_4196, 
        n451, n232_adj_4197, n305_adj_4198, n524, n378_adj_4199, n451_adj_4200, 
        n524_adj_4201, n150, n597, n670, n667_adj_4202, n743, n816, 
        n889, n597_adj_4203, n962, n74, n5_adj_4204, n1035, duty_23__N_3675;
    wire [23:0]duty_23__N_3528;
    
    wire n831, n904, n977, n1050, n223, n670_adj_4205, n147, n1044_adj_4206, 
        n1108, n1117_adj_4207, n743_adj_4208, n98_adj_4209, n29_adj_4210, 
        n296, n104_adj_4211, n816_adj_4212, n171_adj_4213, n244_adj_4214, 
        n889_adj_4215, n35, n317_adj_4216, n390_adj_4217, n177, n962_adj_4218, 
        n463_adj_4219, n536_adj_4220, n220, n250, n609_adj_4221, n673, 
        n682_adj_4222, n1035_adj_4223, n755_adj_4224, n828_adj_4225, 
        n89, n901_adj_4226, n974_adj_4227, n1047_adj_4228, n323, n1120_adj_4229, 
        n396, n469, n101_adj_4230, n32_adj_4231, n542, n615, n20_adj_4232, 
        n162, n174_adj_4233, n247_adj_4234, n688, n235, n320_adj_4235, 
        n17_adj_4236, n9_adj_4237, n11_adj_4238, n31327, n31324, n740_adj_4239, 
        n32765, n31671, n308, n31562, n32747, n31560, n381, n454, 
        n527, n813_adj_4240, n369, n31558, n600_adj_4241, n673_adj_4242, 
        n32741, n27, n15_adj_4243, n13_adj_4244, n11_adj_4245, n31267, 
        n1108_adj_4246, n746, n21_adj_4247, n19_adj_4248, n17_adj_4249, 
        n9_adj_4250, n31273, n43, n16_adj_4251, n31251, n8_adj_4252, 
        n45, n24_adj_4253, n7_adj_4254, n5_adj_4255, n31287, n31534, 
        n31530, n25_adj_4256, n23_adj_4257, n31770, n31, n29_adj_4258, 
        n31647, n37, n35_adj_4259, n33, n31794, n31564, n32734, 
        n31552, n32729, n12_adj_4260, n819, n31299, n32752, n10_adj_4261, 
        n30, n31721, n892, n965, n31307, n32732, n1038, n31665, 
        n32758, n1111, n31774, n32723, n31816, n293, n89_adj_4262, 
        n32720, n20_adj_4263, n366, n16_adj_4264, n31289, n439, 
        n24_adj_4265, n6_adj_4266, n31691, n31692, n31291, n8_adj_4267, 
        n32718, n31625, n31467;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3627 ;
    
    wire n3_adj_4268, n4_adj_4269, n31681, n31682, n12_adj_4270, n31261, 
        n10_adj_4271, n30_adj_4272, n31263, n31784, n31479, n162_adj_4273, 
        n235_adj_4274, n512, n92, n31824, n31825, n39, n31805, 
        n6_adj_4275, n31683, n23_adj_4276, n31684, n31253, n165, 
        n23628, n238, n31627, n31477, n311, n41, n31255, n31750, 
        n31485, n384, n31792, n4_adj_4277, n31689, n31690, n457, 
        n31301, n585, n31782, n31469, n658, n31822, n31823, n530, 
        n31807, n31293, n603, n31748, n31475, \PID_CONTROLLER.integral_23__N_3626 , 
        n31790, n24002, \PID_CONTROLLER.integral_23__N_3624 , n23627, 
        n23626, n676, n308_adj_4278, n731, n381_adj_4279, n804, 
        n877, n454_adj_4280, n950, n1023, n527_adj_4281, n1096, 
        n749, n393_adj_4282, n466_adj_4283, n539_adj_4284, n612_adj_4285, 
        n685_adj_4286, n758_adj_4287;
    wire [23:0]n1_adj_4607;
    
    wire n831_adj_4289, n746_adj_4290, n819_adj_4291, n904_adj_4292, 
        n892_adj_4293, n977_adj_4294, n1050_adj_4295, n965_adj_4296, 
        n104_adj_4297, n35_adj_4298, n1038_adj_4299, n256, n19402, 
        n80, n11_adj_4300, n1111_adj_4301, n153, n177_adj_4302, n226, 
        n250_adj_4303, n299, n372, n445, n518, n92_adj_4306, n23_adj_4307, 
        n165_adj_4309, n591, n323_adj_4310, n396_adj_4311, n469_adj_4312, 
        n542_adj_4313, n615_adj_4314, n688_adj_4315, n761, n834, n907, 
        n980, n107_adj_4316, n38, n238_adj_4317, n311_adj_4318, n384_adj_4319, 
        n664, n457_adj_4320, n530_adj_4321, n180, n603_adj_4322, n676_adj_4323, 
        n749_adj_4324, n253, n737, n326, n399, n472, n545, n618, 
        n691, n764, n837, n910, n110, n41_adj_4326, n183, n256_adj_4327, 
        n329, n402, n475, n548;
    wire [23:0]n257;
    
    wire n33_adj_4328, n12_adj_4329, n621, n694, n767, n840, n113, 
        n44, n186, n259, n332, n405, n478, n822_adj_4333, n551, 
        n624, n697, n770, n116, n47, n189, n262, n335, n408, 
        n481, n554, n627;
    wire [23:0]n1_adj_4608;
    
    wire n700, n119, n50, n192, n265_adj_4353, n338, n442, n886_adj_4355, 
        n761_adj_4356, n23625, n959_adj_4357, n515, n834_adj_4358, 
        n1032_adj_4359, n24001, n23624, n1105_adj_4360, n588, n23623, 
        n661, n907_adj_4362, n484, n980_adj_4363, n107_adj_4365, n38_adj_4366, 
        n180_adj_4367, n24000, n253_adj_4368, n326_adj_4369, n399_adj_4370, 
        n472_adj_4371, n545_adj_4372, n23622, n557, n618_adj_4374, 
        n691_adj_4375, n764_adj_4376, n13_adj_4377, n10_adj_4378, n630, 
        n734, n35_adj_4379, n30_adj_4380, n837_adj_4381, n910_adj_4382, 
        n11_adj_4383, n9_adj_4384, n31210, n31446, n19_adj_4385, n17_adj_4386, 
        n15_adj_4387, n31442, n110_adj_4388, n25_adj_4389, n23_adj_4390, 
        n21_adj_4391, n31738, n41_adj_4392, n183_adj_4393, n256_adj_4394, 
        n329_adj_4395, n402_adj_4396, n122, n31_adj_4397, n29_adj_4398, 
        n27_adj_4399, n31607, n475_adj_4400, n548_adj_4401, n621_adj_4402, 
        n694_adj_4403, n767_adj_4404, n840_adj_4405, n807, n113_adj_4406, 
        n44_adj_4407, n186_adj_4408, n880, n23621, n53, n259_adj_4409, 
        n37_adj_4410, n31786, n1029_adj_4411, n24277, n23620, n332_adj_4412, 
        n23619, n405_adj_4413, n23999, n23618, n23617, n23616, n23615, 
        n478_adj_4415, n23998, n23614, n47_adj_4416, n23768, n23613, 
        n551_adj_4418, n43_adj_4420, n16_adj_4421, n895_adj_4422, n24349, 
        n624_adj_4423, n697_adj_4424, n770_adj_4425, n6_adj_4426, n31728, 
        n31729, n116_adj_4427, n47_adj_4428, n8_adj_4429, n23767, 
        n23612, n956_adj_4432, n24276, n45_adj_4433, n24_adj_4434, 
        n883, n24275, n23997, n23766, n23996, n23765, n189_adj_4438, 
        n31200, n31180, n23764, n262_adj_4441, n31178, n31631, n195, 
        n31702, n268, n341, n31081, n4_adj_4444, n31726, n414, 
        n487, n23763, n31727, n953, n810, n560, n125, n56, n198, 
        n31194, n31190, n23762, n271_adj_4450, n23761, n344, n23995, 
        n4_adj_4454;
    wire [3:0]n7924;
    
    wire n6_adj_4455, n417, n23760, n23994;
    wire [5:0]n7909;
    
    wire n29321, n490, n24707;
    wire [4:0]n7917;
    
    wire n24706, n24705, n23759, n24704, n24703, n23758, n204, 
        n23757;
    wire [6:0]n7900;
    
    wire n24702, n24274;
    wire [1:0]n7935;
    
    wire n24701, n31188, n31800, n24700, n24699, n24698, n23756, 
        n24697, n131, n62, n31704, n23755, n23993, n23754, n23305, 
        n4_adj_4458;
    wire [2:0]n7930;
    
    wire n12_adj_4459;
    wire [7:0]n7890;
    
    wire n24696, n23753, n24695, n8_adj_4460, n23752, n24694, n23751, 
        n11_adj_4461, n411, n24693, n6_adj_4462, n23750, n23992, 
        n23749, n23748, n23407, n24692, n18_adj_4464, n23991, n24691, 
        n23747, n13_adj_4465, n23746, n31836, n4_adj_4466, n31837, 
        n24690;
    wire [8:0]n7879;
    
    wire n24689, n24688, n39_adj_4468, n31819, n23745, n24687, n24686, 
        n24685, n23990, n41_adj_4470, n31182, n23744, n23743, n31760, 
        n23742, n23989, n23741, n23740, n23739, n23382, n23738, 
        n24684, n40, n23988, n24683, n23737, n24682, n23736, n23735, 
        n23734, n23987, n23733, n23732;
    wire [9:0]n7867;
    
    wire n24681, n23731, n24680, n24679, n23730, n31762, n24678, 
        n24348, n24677, n24676, n23986, n23729, n23728, n24675, 
        n24674, n24673, n23985, n23727;
    wire [10:0]n7854;
    
    wire n24672, n24671, n24670, n24669, n24668;
    wire [47:0]n155;
    
    wire n24667, n24666, n24665, n24664, n31114;
    wire [0:0]n5790;
    
    wire n24663;
    wire [11:0]n7840;
    
    wire n24662, n24661, n24660, n24659, n24658, n23726, n24657, 
        n24656, n24655, n24654, n41_adj_4476, n24273, n24653, n39_adj_4477, 
        n24347, n45_adj_4478, n43_adj_4479, n37_adj_4480, n29_adj_4481, 
        n31_adj_4482, n23_adj_4483, n25_adj_4484, n35_adj_4485, n33_adj_4486, 
        n11_adj_4487, n13_adj_4488, n24346, n24345, n15_adj_4489, 
        n27_adj_4490, n9_adj_4491, n17_adj_4492, n24652, n24344, n24343, 
        n24272, n24342, n24341, n24340;
    wire [12:0]n7825;
    
    wire n24651, n24650, n24649, n24648, n24647, n24646, n24645, 
        n24644, n24643, n24642, n19_adj_4493, n24271, n24339, n21_adj_4494, 
        n23725, n23724, n31239, n31230, n24270, n24269, n24268, 
        n24267;
    wire [17:0]n7438;
    
    wire n24338, n23723, n24641, n24337, n24266, n12_adj_4495, n30_adj_4496, 
        n24640, n24336, n31249, n31500, n24265, n24335, n31496, 
        n31764, n31623;
    wire [21:0]n7348;
    
    wire n24264, n31788, n24263, n24334, n24262, n6_adj_4497, n31675, 
        n31676, n24333, n16_adj_4498, n24_adj_4499;
    wire [13:0]n7809;
    
    wire n24639, n24638, n24261, n24332, n24637, n24331, n24330, 
        n24636, n31214, n24635, n24634, n24633, n24632, n8_adj_4500, 
        n31212, n31629, n24631, n24630, n31487, n24629, n24628, 
        n4_adj_4501, n31742, n23250;
    wire [1:0]n7638;
    
    wire n4_adj_4502, n24627;
    wire [2:0]n7633;
    wire [14:0]n7792;
    
    wire n24626, n31743, n31225, n24625, n10_adj_4503, n31223, n31798, 
        n31698, n31834, n24260, n24624, n31835, n31821, n31216, 
        n31754, n40_adj_4504, n31756, n24623, n24622, n24259, n24621, 
        n23216, n4_adj_4505;
    wire [3:0]n7627;
    
    wire n24620, n24329, n24619, n4_adj_4506, n6_adj_4507;
    wire [4:0]n7620;
    
    wire n23173, n24258, n24618, n24617, n24616, n24615, n24614, 
        n24613;
    wire [15:0]n7774;
    
    wire n24612, n24611, n24610, n24609, n24608, n24607, n24606, 
        n24605, n24604, n24603, n24602, n24601, n24600, n24599, 
        n24328, n24598;
    wire [16:0]n7755;
    
    wire n24597, n24596, n24595, n24594, n24593, n24592, n24591, 
        n24590, n24257, n24256, n24327, n24255, n24254, n24326, 
        n24253, n24252, n24325, n24251, n24324, n24589, n24588, 
        n24587, n24250, n24249, n24586, n24585, n24584, n24583, 
        n24582;
    wire [17:0]n7735;
    
    wire n24581, n24580, n24579, n24248, n24323, n24322, n24247, 
        n24246, n24245;
    wire [18:0]n7417;
    
    wire n24321, n24578, n24577, n24320, n24576, n24575, n24574, 
        n24319, n335_adj_4511, n24573, n24318, n24317, n24572, n24571, 
        n24570, n24569, n24568, n24567, n24566, n24565, n24316;
    wire [18:0]n7714;
    
    wire n24564, n24563, n408_adj_4512, n24562, n24244, n24561, 
        n24315, n24314, n24313, n24312, n24560, n24243, n24311, 
        n24559, n24558, n24310, n24557, n481_adj_4513, n24556, n24555, 
        n24554, n24553, n24552, n24551, n24242, n24550, n24309, 
        n24549, n24548, n24308, n24547;
    wire [19:0]n7692;
    
    wire n24546, n24545, n24544, n24241, n24543, n24542, n554_adj_4514, 
        n24240, n24541, n24540, n24539, n24307, n24239, n24538, 
        n24537, n24306, n24305, n24536, n24535, n24534, n24533, 
        n24532, n24531, n24530, n24529, n24528;
    wire [20:0]n7669;
    
    wire n24527, n24526, n24525, n627_adj_4515, n700_adj_4516, n119_adj_4517, 
        n50_adj_4518, n192_adj_4519, n24524, n24523, n24238, n24304, 
        n24522, n24521, n24520, n24519, n883_adj_4520, n24518, n810_adj_4521, 
        n24517, n737_adj_4522, n24516, n664_adj_4523, n24515, n591_adj_4524, 
        n24514, n518_adj_4525, n24513, n445_adj_4526, n24512, n24237, 
        n372_adj_4527, n24511, n299_adj_4528, n24510, n226_adj_4529, 
        n24509, n153_adj_4530, n24508, n11_adj_4531, n80_adj_4532, 
        n24236, n1099, n24235, n17_adj_4533, n86_adj_4534, n1026, 
        n24234;
    wire [21:0]n7645;
    
    wire n24507, n24506, n24505, n24504, n24503, n24502, n24501, 
        n24500, n265_adj_4535, n1096_adj_4536, n24499, n1023_adj_4537, 
        n24498, n950_adj_4538, n24497, n338_adj_4539, n877_adj_4540, 
        n24496, n804_adj_4541, n24495, n731_adj_4542, n24494, n658_adj_4543, 
        n24493, n585_adj_4544, n24492, n512_adj_4545, n24491, n439_adj_4546, 
        n24490, n366_adj_4547, n24489, n293_adj_4548, n24488, n220_adj_4549, 
        n24487, n147_adj_4550, n24486, n5_adj_4551, n74_adj_4552, 
        n24485, n24484, n24483, n24482, n24481, n24480, n24479, 
        n1099_adj_4553, n24478, n1026_adj_4554, n24477, n953_adj_4555, 
        n24476, n880_adj_4556, n24475, n807_adj_4557, n24474, n734_adj_4558, 
        n24473, n661_adj_4559, n24472, n588_adj_4560, n24471, n515_adj_4561, 
        n24470, n442_adj_4562, n24469, n369_adj_4563, n24468, n296_adj_4564, 
        n24467, n223_adj_4565, n24466, n150_adj_4566, n24465, n8_adj_4567, 
        n77_adj_4568;
    wire [5:0]n7612;
    
    wire n29930, n490_adj_4569, n24464, n417_adj_4570, n24463, n344_adj_4571, 
        n24462, n271_adj_4572, n24461, n198_adj_4573, n24460, n56_adj_4574, 
        n125_adj_4575;
    wire [6:0]n7603;
    
    wire n560_adj_4576, n24459, n487_adj_4577, n24458, n414_adj_4578, 
        n24457, n341_adj_4579, n24456, n268_adj_4580, n24455, n195_adj_4581, 
        n24454, n53_adj_4582, n122_adj_4583;
    wire [7:0]n7593;
    
    wire n630_adj_4584, n24453, n557_adj_4585, n24452, n484_adj_4586, 
        n24451, n411_adj_4587, n24450, n24449, n24448, n24447;
    wire [8:0]n7582;
    
    wire n24446, n24445, n24444, n24443, n24442, n24441, n24233, 
        n24440, n24439;
    wire [9:0]n7570;
    
    wire n24438, n24437, n24303, n24436, n24435, n24434, n24433, 
        n24432, n24302, n24431, n24232, n24430, n24231;
    wire [10:0]n7557;
    
    wire n24429, n24428, n24427, n24426, n24425, n24424, n24423, 
        n24422, n24421, n24420, n24301;
    wire [11:0]n7543;
    
    wire n24419, n24418, n24230, n24300, n24417, n24416, n24415, 
        n24414, n24413, n24412, n24411, n24410, n24409;
    wire [12:0]n7528;
    
    wire n24408, n24407, n24229, n24228, n24299, n24298, n24297, 
        n24406, n24227, n24296, n24405, n24295, n24226, n24225, 
        n24294, n24293, n24404, n24403, n24402, n24401, n24400, 
        n24399, n24398, n24397, n24224, n24223, n12_adj_4588;
    wire [13:0]n7512;
    
    wire n24396, n8_adj_4589, n11_adj_4590, n6_adj_4591, n24395, n24394, 
        n24393, n23275, n18_adj_4592, n24292, n13_adj_4593, n24222, 
        n24392, n24291, n24391, n24290, n24289, n24288, n24287, 
        n24390, n24389, n24388, n24387, n24386, n24385, n24286, 
        n24384, n24285;
    wire [14:0]n7495;
    
    wire n24383, n24382, n24381, n24380, n24284, n24379, n24283, 
        n24378, n24377, n24376, n24375, n24374, n24373, n24372, 
        n24371, n24282, n24370, n24369, n24368, n24367, n24366, 
        n24365, n825_adj_4594, n24364, n752_adj_4595, n24363, n679_adj_4596, 
        n24362, n606_adj_4597, n24361, n533_adj_4598, n24360, n460_adj_4599, 
        n24359, n387_adj_4600, n24358, n314_adj_4601, n24357, n241_adj_4602, 
        n24356, n168_adj_4603, n24355, n26_adj_4604, n95_adj_4605, 
        n24354, n24353, n1114_adj_4606;
    
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3441_18 (.CI(n24280), .I0(n7395[15]), .I1(GND_net), .CO(n24281));
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3441_17_lut (.I0(GND_net), .I1(n7395[14]), .I2(GND_net), 
            .I3(n24279), .O(n7372[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4179));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4180));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4181));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4182));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1[23]), .I3(n23657), .O(\PID_CONTROLLER.err_23__N_3552 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1[22]), .I3(n23656), .O(\PID_CONTROLLER.err_23__N_3552 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n23656), .I0(motor_state[22]), 
            .I1(n1[22]), .CO(n23657));
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1[21]), .I3(n23655), .O(\PID_CONTROLLER.err_23__N_3552 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n23655), .I0(motor_state[21]), 
            .I1(n1[21]), .CO(n23656));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1[20]), .I3(n23654), .O(\PID_CONTROLLER.err_23__N_3552 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n23654), .I0(motor_state[20]), 
            .I1(n1[20]), .CO(n23655));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1[19]), .I3(n23653), .O(\PID_CONTROLLER.err_23__N_3552 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n23653), .I0(motor_state[19]), 
            .I1(n1[19]), .CO(n23654));
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1[18]), .I3(n23652), .O(\PID_CONTROLLER.err_23__N_3552 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n23652), .I0(motor_state[18]), 
            .I1(n1[18]), .CO(n23653));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1[17]), .I3(n23651), .O(\PID_CONTROLLER.err_23__N_3552 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n23651), .I0(motor_state[17]), 
            .I1(n1[17]), .CO(n23652));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1[16]), .I3(n23650), .O(\PID_CONTROLLER.err_23__N_3552 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n23650), .I0(motor_state[16]), 
            .I1(n1[16]), .CO(n23651));
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1[15]), .I3(n23649), .O(\PID_CONTROLLER.err_23__N_3552 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n23649), .I0(motor_state[15]), 
            .I1(n1[15]), .CO(n23650));
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1[14]), .I3(n23648), .O(\PID_CONTROLLER.err_23__N_3552 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n23648), .I0(motor_state[14]), 
            .I1(n1[14]), .CO(n23649));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1[13]), .I3(n23647), .O(\PID_CONTROLLER.err_23__N_3552 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n23647), .I0(motor_state[13]), 
            .I1(n1[13]), .CO(n23648));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1[12]), .I3(n23646), .O(\PID_CONTROLLER.err_23__N_3552 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n23646), .I0(motor_state[12]), 
            .I1(n1[12]), .CO(n23647));
    SB_CARRY add_3445_15 (.CI(n24351), .I0(n7477[12]), .I1(n1041), .CO(n24352));
    SB_CARRY add_3441_17 (.CI(n24279), .I0(n7395[14]), .I1(GND_net), .CO(n24280));
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1[11]), .I3(n23645), .O(\PID_CONTROLLER.err_23__N_3552 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n23645), .I0(motor_state[11]), 
            .I1(n1[11]), .CO(n23646));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1[10]), .I3(n23644), .O(\PID_CONTROLLER.err_23__N_3552 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n23644), .I0(motor_state[10]), 
            .I1(n1[10]), .CO(n23645));
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n24007), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1[9]), .I3(n23643), .O(\PID_CONTROLLER.err_23__N_3552 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n23643), .I0(motor_state[9]), .I1(n1[9]), 
            .CO(n23644));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1[8]), .I3(n23642), .O(\PID_CONTROLLER.err_23__N_3552 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n23642), .I0(motor_state[8]), .I1(n1[8]), 
            .CO(n23643));
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n24006), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1[7]), .I3(n23641), .O(\PID_CONTROLLER.err_23__N_3552 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_9 (.CI(n23641), .I0(motor_state[7]), .I1(n1[7]), 
            .CO(n23642));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1[6]), .I3(n23640), .O(\PID_CONTROLLER.err_23__N_3552 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n23640), .I0(motor_state[6]), .I1(n1[6]), 
            .CO(n23641));
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_24  (.CI(n24006), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n24007));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1[5]), .I3(n23639), .O(\PID_CONTROLLER.err_23__N_3552 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n23639), .I0(motor_state[5]), .I1(n1[5]), 
            .CO(n23640));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1[4]), .I3(n23638), .O(\PID_CONTROLLER.err_23__N_3552 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n23638), .I0(motor_state[4]), .I1(n1[4]), 
            .CO(n23639));
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n24005), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1[3]), .I3(n23637), .O(\PID_CONTROLLER.err_23__N_3552 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n23637), .I0(motor_state[3]), .I1(n1[3]), 
            .CO(n23638));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1[2]), .I3(n23636), .O(\PID_CONTROLLER.err_23__N_3552 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n23636), .I0(motor_state[2]), .I1(n1[2]), 
            .CO(n23637));
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_23  (.CI(n24005), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n24006));
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1[1]), .I3(n23635), .O(\PID_CONTROLLER.err_23__N_3552 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n23635), .I0(motor_state[1]), .I1(n1[1]), 
            .CO(n23636));
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3552 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1[0]), 
            .CO(n23635));
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n24004), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_25_lut (.I0(GND_net), .I1(n2901[23]), .I2(n2926[23]), 
            .I3(n23634), .O(duty_23__N_3651[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_609_24_lut (.I0(GND_net), .I1(n2901[22]), .I2(n2926[22]), 
            .I3(n23633), .O(duty_23__N_3651[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_24 (.CI(n23633), .I0(n2901[22]), .I1(n2926[22]), 
            .CO(n23634));
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_23_lut (.I0(GND_net), .I1(n2901[21]), .I2(n2926[21]), 
            .I3(n23632), .O(duty_23__N_3651[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_22  (.CI(n24004), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n24005));
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4184));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4185));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_23 (.CI(n23632), .I0(n2901[21]), .I1(n2926[21]), 
            .CO(n23633));
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4186));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4187));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4188));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_22_lut (.I0(GND_net), .I1(n2901[20]), .I2(n2926[20]), 
            .I3(n23631), .O(duty_23__N_3651[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_22 (.CI(n23631), .I0(n2901[20]), .I1(n2926[20]), 
            .CO(n23632));
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4189));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4190));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_21_lut (.I0(GND_net), .I1(n2901[19]), .I2(n2926[19]), 
            .I3(n23630), .O(duty_23__N_3651[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4191));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3445_14_lut (.I0(GND_net), .I1(n7477[11]), .I2(n968_adj_4192), 
            .I3(n24350), .O(n7458[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_21 (.CI(n23630), .I0(n2901[19]), .I1(n2926[19]), 
            .CO(n23631));
    SB_LUT4 add_609_20_lut (.I0(GND_net), .I1(n2901[18]), .I2(n2926[18]), 
            .I3(n23629), .O(duty_23__N_3651[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3441_16_lut (.I0(GND_net), .I1(n7395[13]), .I2(n1102_adj_4193), 
            .I3(n24278), .O(n7372[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4194));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n24003), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4195));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4196));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4197));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4198));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4199));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4200));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4201));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4202));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_20 (.CI(n23629), .I0(n2901[18]), .I1(n2926[18]), 
            .CO(n23630));
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4203));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4204));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3651[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3651[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3651[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3651[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3651[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3651[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3651[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3651[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3651[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3651[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3651[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3651[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3651[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3651[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3651[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3651[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3651[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3651[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3651[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3651[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3651[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4205));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4206));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4207));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4208));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4209));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4210));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4211));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4212));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4213));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4214));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4215));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4216));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4217));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4218));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4219));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4220));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4221));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4222));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4223));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4224));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4225));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4226));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4227));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4228));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4229));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4230));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4231));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4232));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4233));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4234));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4235));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4236));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4237));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4238));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25496_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n31327));
    defparam i25496_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i25493_3_lut (.I0(n11_adj_4238), .I1(n9_adj_4237), .I2(n31327), 
            .I3(GND_net), .O(n31324));
    defparam i25493_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4239));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_172_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n32765));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_172_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25838_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n32765), 
            .I2(IntegralLimit[7]), .I3(n31324), .O(n31671));
    defparam i25838_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25729_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4236), 
            .I2(IntegralLimit[9]), .I3(n31671), .O(n31562));
    defparam i25729_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_154_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n32747));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_154_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25727_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4236), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4237), .O(n31560));
    defparam i25727_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4240));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25725_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n32747), 
            .I2(IntegralLimit[11]), .I3(n31560), .O(n31558));
    defparam i25725_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4241));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4242));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_148_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n32741));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_148_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25436_4_lut (.I0(n27), .I1(n15_adj_4243), .I2(n13_adj_4244), 
            .I3(n11_adj_4245), .O(n31267));
    defparam i25436_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4246));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3651[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25442_4_lut (.I0(n21_adj_4247), .I1(n19_adj_4248), .I2(n17_adj_4249), 
            .I3(n9_adj_4250), .O(n31273));
    defparam i25442_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4251));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i25420_2_lut (.I0(n43), .I1(n19_adj_4248), .I2(GND_net), .I3(GND_net), 
            .O(n31251));
    defparam i25420_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4249), .I3(GND_net), 
            .O(n8_adj_4252));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4251), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4253));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i25456_2_lut (.I0(n7_adj_4254), .I1(n5_adj_4255), .I2(GND_net), 
            .I3(GND_net), .O(n31287));
    defparam i25456_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i25701_4_lut (.I0(n13_adj_4244), .I1(n11_adj_4245), .I2(n9_adj_4250), 
            .I3(n31287), .O(n31534));
    defparam i25701_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i25697_4_lut (.I0(n19_adj_4248), .I1(n17_adj_4249), .I2(n15_adj_4243), 
            .I3(n31534), .O(n31530));
    defparam i25697_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i25937_4_lut (.I0(n25_adj_4256), .I1(n23_adj_4257), .I2(n21_adj_4247), 
            .I3(n31530), .O(n31770));
    defparam i25937_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25814_4_lut (.I0(n31), .I1(n29_adj_4258), .I2(n27), .I3(n31770), 
            .O(n31647));
    defparam i25814_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i25961_4_lut (.I0(n37), .I1(n35_adj_4259), .I2(n33), .I3(n31647), 
            .O(n31794));
    defparam i25961_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25731_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n32765), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4238), .O(n31564));
    defparam i25731_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_141_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n32734));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_141_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25719_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n32734), 
            .I2(IntegralLimit[14]), .I3(n31564), .O(n31552));
    defparam i25719_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_136_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n32729));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_136_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4260));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25468_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n31299));
    defparam i25468_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_159_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n32752));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_159_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4261));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4260), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25888_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n32747), 
            .I2(IntegralLimit[11]), .I3(n31562), .O(n31721));
    defparam i25888_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25476_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n32741), 
            .I2(IntegralLimit[13]), .I3(n31721), .O(n31307));
    defparam i25476_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_139_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n32732));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_139_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25832_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n32732), 
            .I2(IntegralLimit[15]), .I3(n31307), .O(n31665));
    defparam i25832_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_165_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n32758));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_165_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25941_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n32758), 
            .I2(IntegralLimit[17]), .I3(n31665), .O(n31774));
    defparam i25941_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_130_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n32723));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_130_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25983_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n32723), 
            .I2(IntegralLimit[19]), .I3(n31774), .O(n31816));
    defparam i25983_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4262));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_127_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n32720));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_127_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4263));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4264));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25458_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n31289));
    defparam i25458_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4264), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4265));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4266));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25858_3_lut (.I0(n6_adj_4266), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n31691));   // verilog/motorControl.v(31[10:34])
    defparam i25858_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25859_3_lut (.I0(n31691), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n31692));   // verilog/motorControl.v(31[10:34])
    defparam i25859_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25460_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n32741), 
            .I2(IntegralLimit[21]), .I3(n31558), .O(n31291));
    defparam i25460_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i25792_4_lut (.I0(n24_adj_4265), .I1(n8_adj_4267), .I2(n32718), 
            .I3(n31289), .O(n31625));   // verilog/motorControl.v(31[10:34])
    defparam i25792_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i25634_3_lut (.I0(n31692), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n31467));   // verilog/motorControl.v(31[10:34])
    defparam i25634_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3627 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4268), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4269));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i25848_3_lut (.I0(n4_adj_4269), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n31681));   // verilog/motorControl.v(31[38:63])
    defparam i25848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25849_3_lut (.I0(n31681), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4258), .I3(GND_net), .O(n31682));   // verilog/motorControl.v(31[38:63])
    defparam i25849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4270));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i25430_2_lut (.I0(n33), .I1(n15_adj_4243), .I2(GND_net), .I3(GND_net), 
            .O(n31261));
    defparam i25430_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4244), .I3(GND_net), 
            .O(n10_adj_4271));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4270), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4259), .I3(GND_net), 
            .O(n30_adj_4272));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i25432_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4258), .I3(n31267), 
            .O(n31263));
    defparam i25432_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i25951_4_lut (.I0(n30_adj_4272), .I1(n10_adj_4271), .I2(n35_adj_4259), 
            .I3(n31261), .O(n31784));   // verilog/motorControl.v(31[38:63])
    defparam i25951_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i25646_3_lut (.I0(n31682), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n31479));   // verilog/motorControl.v(31[38:63])
    defparam i25646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4273));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4274));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25991_4_lut (.I0(n31479), .I1(n31784), .I2(n35_adj_4259), 
            .I3(n31263), .O(n31824));   // verilog/motorControl.v(31[38:63])
    defparam i25991_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25992_3_lut (.I0(n31824), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n31825));   // verilog/motorControl.v(31[38:63])
    defparam i25992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25972_3_lut (.I0(n31825), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n31805));   // verilog/motorControl.v(31[38:63])
    defparam i25972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4254), .I3(GND_net), 
            .O(n6_adj_4275));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i25850_3_lut (.I0(n6_adj_4275), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4247), .I3(GND_net), .O(n31683));   // verilog/motorControl.v(31[38:63])
    defparam i25850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4276));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25851_3_lut (.I0(n31683), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4257), .I3(GND_net), .O(n31684));   // verilog/motorControl.v(31[38:63])
    defparam i25851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25422_4_lut (.I0(n43), .I1(n25_adj_4256), .I2(n23_adj_4257), 
            .I3(n31273), .O(n31253));
    defparam i25422_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_19_lut (.I0(GND_net), .I1(n2901[17]), .I2(n2926[17]), 
            .I3(n23628), .O(duty_23__N_3651[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25794_4_lut (.I0(n24_adj_4253), .I1(n8_adj_4252), .I2(n45), 
            .I3(n31251), .O(n31627));   // verilog/motorControl.v(31[38:63])
    defparam i25794_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i25644_3_lut (.I0(n31684), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4256), .I3(GND_net), .O(n31477));   // verilog/motorControl.v(31[38:63])
    defparam i25644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25424_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n31794), 
            .O(n31255));
    defparam i25424_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i25917_4_lut (.I0(n31477), .I1(n31627), .I2(n45), .I3(n31253), 
            .O(n31750));   // verilog/motorControl.v(31[38:63])
    defparam i25917_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25652_3_lut (.I0(n31805), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41), .I3(GND_net), .O(n31485));   // verilog/motorControl.v(31[38:63])
    defparam i25652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_19 (.CI(n23628), .I0(n2901[17]), .I1(n2926[17]), 
            .CO(n23629));
    SB_LUT4 i25959_4_lut (.I0(n31485), .I1(n31750), .I2(n45), .I3(n31255), 
            .O(n31792));   // verilog/motorControl.v(31[38:63])
    defparam i25959_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4277));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i25856_3_lut (.I0(n4_adj_4277), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n31689));   // verilog/motorControl.v(31[10:34])
    defparam i25856_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25857_3_lut (.I0(n31689), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n31690));   // verilog/motorControl.v(31[10:34])
    defparam i25857_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25470_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n32729), 
            .I2(IntegralLimit[16]), .I3(n31552), .O(n31301));
    defparam i25470_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25949_4_lut (.I0(n30), .I1(n10_adj_4261), .I2(n32752), .I3(n31299), 
            .O(n31782));   // verilog/motorControl.v(31[10:34])
    defparam i25949_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i25636_3_lut (.I0(n31690), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n31469));   // verilog/motorControl.v(31[10:34])
    defparam i25636_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25989_4_lut (.I0(n31469), .I1(n31782), .I2(n32752), .I3(n31301), 
            .O(n31822));   // verilog/motorControl.v(31[10:34])
    defparam i25989_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25990_3_lut (.I0(n31822), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n31823));   // verilog/motorControl.v(31[10:34])
    defparam i25990_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25974_3_lut (.I0(n31823), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n31807));   // verilog/motorControl.v(31[10:34])
    defparam i25974_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25462_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n32720), 
            .I2(IntegralLimit[21]), .I3(n31816), .O(n31293));
    defparam i25462_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_125_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n32718));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_125_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_21  (.CI(n24003), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n24004));
    SB_LUT4 i25915_4_lut (.I0(n31467), .I1(n31625), .I2(n32718), .I3(n31291), 
            .O(n31748));   // verilog/motorControl.v(31[10:34])
    defparam i25915_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25642_3_lut (.I0(n31807), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n31475));   // verilog/motorControl.v(31[10:34])
    defparam i25642_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25960_3_lut (.I0(n31792), .I1(\PID_CONTROLLER.integral_23__N_3627 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3626 ));   // verilog/motorControl.v(31[38:63])
    defparam i25960_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3441_16 (.CI(n24278), .I0(n7395[13]), .I1(n1102_adj_4193), 
            .CO(n24279));
    SB_LUT4 i25957_4_lut (.I0(n31475), .I1(n31748), .I2(n32718), .I3(n31293), 
            .O(n31790));   // verilog/motorControl.v(31[10:34])
    defparam i25957_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n24002), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_838_4_lut  (.I0(n31790), .I1(\PID_CONTROLLER.integral_23__N_3626 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3624 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_838_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 add_609_18_lut (.I0(GND_net), .I1(n2901[16]), .I2(n2926[16]), 
            .I3(n23627), .O(duty_23__N_3651[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_18 (.CI(n23627), .I0(n2901[16]), .I1(n2926[16]), 
            .CO(n23628));
    SB_LUT4 add_609_17_lut (.I0(GND_net), .I1(n2901[15]), .I2(n2926[15]), 
            .I3(n23626), .O(duty_23__N_3651[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4278));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4279));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4280));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4281));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3651[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4282));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4283));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4284));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4285));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4286));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4287));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4289));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4290));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4291));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4292));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4293));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4294));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4295));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4296));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4297));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4298));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4299));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14870_1_lut (.I0(n256), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n19402));   // verilog/motorControl.v(38[19:35])
    defparam i14870_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4300));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4301));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4302));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4303));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_609_17 (.CI(n23626), .I0(n2901[15]), .I1(n2926[15]), 
            .CO(n23627));
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4306));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4307));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4309));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4310));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4311));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4312));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4313));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4314));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4315));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4316));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4317));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4318));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4319));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4320));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4321));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4322));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4323));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4324));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4326));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4327));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4328), 
            .I3(GND_net), .O(n12_adj_4329));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4333));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[0]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_20  (.CI(n24002), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n24003));
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[1]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[2]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4353));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[3]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4355));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4356));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_16_lut (.I0(GND_net), .I1(n2901[14]), .I2(n2926[14]), 
            .I3(n23625), .O(duty_23__N_3651[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4357));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4358));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4359));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n24001), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_609_16 (.CI(n23625), .I0(n2901[14]), .I1(n2926[14]), 
            .CO(n23626));
    SB_LUT4 add_609_15_lut (.I0(GND_net), .I1(n2901[13]), .I2(n2926[13]), 
            .I3(n23624), .O(duty_23__N_3651[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4360));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_15 (.CI(n23624), .I0(n2901[13]), .I1(n2926[13]), 
            .CO(n23625));
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[6]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3528[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_14_lut (.I0(GND_net), .I1(n2901[12]), .I2(n2926[12]), 
            .I3(n23623), .O(duty_23__N_3651[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4362));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4363));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[7]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_19  (.CI(n24001), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n24002));
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4365));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4366));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4367));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n24000), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_609_14 (.CI(n23623), .I0(n2901[12]), .I1(n2926[12]), 
            .CO(n23624));
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4368));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4369));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4370));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4371));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4372));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_13_lut (.I0(GND_net), .I1(n2901[11]), .I2(n2926[11]), 
            .I3(n23622), .O(duty_23__N_3651[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[8]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4374));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4375));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4376));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4377), 
            .I3(GND_net), .O(n10_adj_4378));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4329), .I1(n257[17]), .I2(n35_adj_4379), 
            .I3(GND_net), .O(n30_adj_4380));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4381));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4382));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25613_4_lut (.I0(n13_adj_4377), .I1(n11_adj_4383), .I2(n9_adj_4384), 
            .I3(n31210), .O(n31446));
    defparam i25613_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i25609_4_lut (.I0(n19_adj_4385), .I1(n17_adj_4386), .I2(n15_adj_4387), 
            .I3(n31446), .O(n31442));
    defparam i25609_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4388));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25905_4_lut (.I0(n25_adj_4389), .I1(n23_adj_4390), .I2(n21_adj_4391), 
            .I3(n31442), .O(n31738));
    defparam i25905_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4392));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4393));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4394));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_13 (.CI(n23622), .I0(n2901[11]), .I1(n2926[11]), 
            .CO(n23623));
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4395));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4396));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25774_4_lut (.I0(n31_adj_4397), .I1(n29_adj_4398), .I2(n27_adj_4399), 
            .I3(n31738), .O(n31607));
    defparam i25774_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4400));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4401));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4402));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4403));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4404));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4405));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4406));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4407));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4408));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_12_lut (.I0(GND_net), .I1(n2901[10]), .I2(n2926[10]), 
            .I3(n23621), .O(duty_23__N_3651[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4409));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_12 (.CI(n23621), .I0(n2901[10]), .I1(n2926[10]), 
            .CO(n23622));
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_18  (.CI(n24000), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n24001));
    SB_LUT4 i25953_4_lut (.I0(n37_adj_4410), .I1(n35_adj_4379), .I2(n33_adj_4328), 
            .I3(n31607), .O(n31786));
    defparam i25953_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3441_15_lut (.I0(GND_net), .I1(n7395[12]), .I2(n1029_adj_4411), 
            .I3(n24277), .O(n7372[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_609_11_lut (.I0(GND_net), .I1(n2901[9]), .I2(n2926[9]), 
            .I3(n23620), .O(duty_23__N_3651[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_11 (.CI(n23620), .I0(n2901[9]), .I1(n2926[9]), .CO(n23621));
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4412));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_609_10_lut (.I0(GND_net), .I1(n2901[8]), .I2(n2926[8]), 
            .I3(n23619), .O(duty_23__N_3651[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_14 (.CI(n24350), .I0(n7477[11]), .I1(n968_adj_4192), 
            .CO(n24351));
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4413));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_10 (.CI(n23619), .I0(n2901[8]), .I1(n2926[8]), .CO(n23620));
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n23999), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_609_9_lut (.I0(GND_net), .I1(n2901[7]), .I2(n2926[7]), 
            .I3(n23618), .O(duty_23__N_3651[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_9 (.CI(n23618), .I0(n2901[7]), .I1(n2926[7]), .CO(n23619));
    SB_LUT4 add_609_8_lut (.I0(GND_net), .I1(n2901[6]), .I2(n2926[6]), 
            .I3(n23617), .O(duty_23__N_3651[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_8 (.CI(n23617), .I0(n2901[6]), .I1(n2926[6]), .CO(n23618));
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_17  (.CI(n23999), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n24000));
    SB_LUT4 add_609_7_lut (.I0(GND_net), .I1(n2901[5]), .I2(n2926[5]), 
            .I3(n23616), .O(duty_23__N_3651[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_7 (.CI(n23616), .I0(n2901[5]), .I1(n2926[5]), .CO(n23617));
    SB_LUT4 add_609_6_lut (.I0(GND_net), .I1(n2901[4]), .I2(n2926[4]), 
            .I3(n23615), .O(duty_23__N_3651[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_6 (.CI(n23615), .I0(n2901[4]), .I1(n2926[4]), .CO(n23616));
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4415));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n23998), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_15 (.CI(n24277), .I0(n7395[12]), .I1(n1029_adj_4411), 
            .CO(n24278));
    SB_LUT4 add_609_5_lut (.I0(GND_net), .I1(n2901[3]), .I2(n2926[3]), 
            .I3(n23614), .O(duty_23__N_3651[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_609_5 (.CI(n23614), .I0(n2901[3]), .I1(n2926[3]), .CO(n23615));
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_16  (.CI(n23998), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n23999));
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1_adj_4608[23]), 
            .I3(n23768), .O(n47_adj_4416)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_609_4_lut (.I0(GND_net), .I1(n2901[2]), .I2(n2926[2]), 
            .I3(n23613), .O(duty_23__N_3651[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4418));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[9]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4420), 
            .I3(GND_net), .O(n16_adj_4421));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3445_13_lut (.I0(GND_net), .I1(n7477[10]), .I2(n895_adj_4422), 
            .I3(n24349), .O(n7458[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4423));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4424));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4425));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25895_3_lut (.I0(n6_adj_4426), .I1(n257[10]), .I2(n21_adj_4391), 
            .I3(GND_net), .O(n31728));   // verilog/motorControl.v(38[19:35])
    defparam i25895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25896_3_lut (.I0(n31728), .I1(n257[11]), .I2(n23_adj_4390), 
            .I3(GND_net), .O(n31729));   // verilog/motorControl.v(38[19:35])
    defparam i25896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4427));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4428));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_609_4 (.CI(n23613), .I0(n2901[2]), .I1(n2926[2]), .CO(n23614));
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4386), 
            .I3(GND_net), .O(n8_adj_4429));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[22]), 
            .I3(n23767), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_609_3_lut (.I0(GND_net), .I1(n2901[1]), .I2(n2926[1]), 
            .I3(n23612), .O(duty_23__N_3651[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_13 (.CI(n24349), .I0(n7477[10]), .I1(n895_adj_4422), 
            .CO(n24350));
    SB_CARRY add_609_3 (.CI(n23612), .I0(n2901[1]), .I1(n2926[1]), .CO(n23613));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n23767), .I0(GND_net), .I1(n1_adj_4608[22]), 
            .CO(n23768));
    SB_LUT4 add_609_2_lut (.I0(GND_net), .I1(n2901[0]), .I2(n2926[0]), 
            .I3(GND_net), .O(duty_23__N_3651[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_609_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_14_lut (.I0(GND_net), .I1(n7395[11]), .I2(n956_adj_4432), 
            .I3(n24276), .O(n7372[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3441_14 (.CI(n24276), .I0(n7395[11]), .I1(n956_adj_4432), 
            .CO(n24277));
    SB_CARRY add_609_2 (.CI(GND_net), .I0(n2901[0]), .I1(n2926[0]), .CO(n23612));
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4421), .I1(n257[22]), .I2(n45_adj_4433), 
            .I3(GND_net), .O(n24_adj_4434));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3441_13_lut (.I0(GND_net), .I1(n7395[10]), .I2(n883), 
            .I3(n24275), .O(n7372[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n23997), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_15  (.CI(n23997), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n23998));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[21]), 
            .I3(n23766), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n23766), .I0(GND_net), .I1(n1_adj_4608[21]), 
            .CO(n23767));
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n23996), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[20]), 
            .I3(n23765), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4438));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25349_4_lut (.I0(n43_adj_4420), .I1(n25_adj_4389), .I2(n23_adj_4390), 
            .I3(n31200), .O(n31180));
    defparam i25349_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n23765), .I0(GND_net), .I1(n1_adj_4608[20]), 
            .CO(n23766));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[19]), 
            .I3(n23764), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4441));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[10]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n23764), .I0(GND_net), .I1(n1_adj_4608[19]), 
            .CO(n23765));
    SB_LUT4 i25798_4_lut (.I0(n24_adj_4434), .I1(n8_adj_4429), .I2(n45_adj_4433), 
            .I3(n31178), .O(n31631));   // verilog/motorControl.v(38[19:35])
    defparam i25798_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[11]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25869_3_lut (.I0(n31729), .I1(n257[12]), .I2(n25_adj_4389), 
            .I3(GND_net), .O(n31702));   // verilog/motorControl.v(38[19:35])
    defparam i25869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n31081), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_4444));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25893_3_lut (.I0(n4_adj_4444), .I1(n257[13]), .I2(n27_adj_4399), 
            .I3(GND_net), .O(n31726));   // verilog/motorControl.v(38[19:35])
    defparam i25893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[18]), 
            .I3(n23763), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25894_3_lut (.I0(n31726), .I1(n257[14]), .I2(n29_adj_4398), 
            .I3(GND_net), .O(n31727));   // verilog/motorControl.v(38[19:35])
    defparam i25894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n23763), .I0(GND_net), .I1(n1_adj_4608[18]), 
            .CO(n23764));
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3441_13 (.CI(n24275), .I0(n7395[10]), .I1(n883), .CO(n24276));
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[12]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[13]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25359_4_lut (.I0(n33_adj_4328), .I1(n31_adj_4397), .I2(n29_adj_4398), 
            .I3(n31194), .O(n31190));
    defparam i25359_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_14  (.CI(n23996), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n23997));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[17]), 
            .I3(n23762), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4450));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n23762), .I0(GND_net), .I1(n1_adj_4608[17]), 
            .CO(n23763));
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[4]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[16]), 
            .I3(n23761), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[14]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n23761), .I0(GND_net), .I1(n1_adj_4608[16]), 
            .CO(n23762));
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n23995), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i18794_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_4454), .I3(n7924[1]), .O(n6_adj_4455));   // verilog/motorControl.v(34[26:37])
    defparam i18794_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_13  (.CI(n23995), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n23996));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[15]), 
            .I3(n23760), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n23994), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3478_7_lut (.I0(GND_net), .I1(n29321), .I2(n490), .I3(n24707), 
            .O(n7909[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3478_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n23760), .I0(GND_net), .I1(n1_adj_4608[15]), 
            .CO(n23761));
    SB_LUT4 add_3478_6_lut (.I0(GND_net), .I1(n7917[3]), .I2(n417), .I3(n24706), 
            .O(n7909[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3478_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3478_6 (.CI(n24706), .I0(n7917[3]), .I1(n417), .CO(n24707));
    SB_LUT4 add_3478_5_lut (.I0(GND_net), .I1(n7917[2]), .I2(n344), .I3(n24705), 
            .O(n7909[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3478_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[14]), 
            .I3(n23759), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3478_5 (.CI(n24705), .I0(n7917[2]), .I1(n344), .CO(n24706));
    SB_LUT4 i2_4_lut (.I0(n6_adj_4455), .I1(\Ki[4] ), .I2(n7924[2]), .I3(\PID_CONTROLLER.integral [18]), 
            .O(n7917[3]));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 add_3478_4_lut (.I0(GND_net), .I1(n7917[1]), .I2(n271_adj_4450), 
            .I3(n24704), .O(n7909[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3478_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3478_4 (.CI(n24704), .I0(n7917[1]), .I1(n271_adj_4450), 
            .CO(n24705));
    SB_LUT4 add_3478_3_lut (.I0(GND_net), .I1(n7917[0]), .I2(n198), .I3(n24703), 
            .O(n7909[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3478_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n23759), .I0(GND_net), .I1(n1_adj_4608[14]), 
            .CO(n23760));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[13]), 
            .I3(n23758), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n23758), .I0(GND_net), .I1(n1_adj_4608[13]), 
            .CO(n23759));
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3478_3 (.CI(n24703), .I0(n7917[0]), .I1(n198), .CO(n24704));
    SB_LUT4 add_3478_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n7909[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3478_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3478_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n24703));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[12]), 
            .I3(n23757), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3477_8_lut (.I0(GND_net), .I1(n7909[5]), .I2(n560), .I3(n24702), 
            .O(n7900[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3477_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_12  (.CI(n23994), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n23995));
    SB_LUT4 add_3441_12_lut (.I0(GND_net), .I1(n7395[9]), .I2(n810), .I3(n24274), 
            .O(n7372[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n23757), .I0(GND_net), .I1(n1_adj_4608[12]), 
            .CO(n23758));
    SB_LUT4 i18866_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n7935[0]));   // verilog/motorControl.v(34[26:37])
    defparam i18866_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_3477_7_lut (.I0(GND_net), .I1(n7909[4]), .I2(n487), .I3(n24701), 
            .O(n7900[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3477_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3477_7 (.CI(n24701), .I0(n7909[4]), .I1(n487), .CO(n24702));
    SB_LUT4 i25967_4_lut (.I0(n30_adj_4380), .I1(n10_adj_4378), .I2(n35_adj_4379), 
            .I3(n31188), .O(n31800));   // verilog/motorControl.v(38[19:35])
    defparam i25967_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3477_6_lut (.I0(GND_net), .I1(n7909[3]), .I2(n414), .I3(n24700), 
            .O(n7900[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3477_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3477_6 (.CI(n24700), .I0(n7909[3]), .I1(n414), .CO(n24701));
    SB_LUT4 add_3477_5_lut (.I0(GND_net), .I1(n7909[2]), .I2(n341), .I3(n24699), 
            .O(n7900[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3477_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3477_5 (.CI(n24699), .I0(n7909[2]), .I1(n341), .CO(n24700));
    SB_LUT4 add_3477_4_lut (.I0(GND_net), .I1(n7909[1]), .I2(n268), .I3(n24698), 
            .O(n7900[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3477_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3477_4 (.CI(n24698), .I0(n7909[1]), .I1(n268), .CO(n24699));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[11]), 
            .I3(n23756), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3477_3_lut (.I0(GND_net), .I1(n7909[0]), .I2(n195), .I3(n24697), 
            .O(n7900[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3477_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n23756), .I0(GND_net), .I1(n1_adj_4608[11]), 
            .CO(n23757));
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25871_3_lut (.I0(n31727), .I1(n257[15]), .I2(n31_adj_4397), 
            .I3(GND_net), .O(n31704));   // verilog/motorControl.v(38[19:35])
    defparam i25871_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3477_3 (.CI(n24697), .I0(n7909[0]), .I1(n195), .CO(n24698));
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n7924[1]), .I3(n4_adj_4454), .O(n7917[2]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[10]), 
            .I3(n23755), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n23993), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n23755), .I0(GND_net), .I1(n1_adj_4608[10]), 
            .CO(n23756));
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[9]), 
            .I3(n23754), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1473 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n7924[0]), .I3(n23305), .O(n7917[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1473.LUT_INIT = 16'h8778;
    SB_LUT4 i2_4_lut_adj_1474 (.I0(n4_adj_4458), .I1(\Ki[3] ), .I2(n7930[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n7924[2]));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut_adj_1474.LUT_INIT = 16'h965a;
    SB_LUT4 add_3477_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n7900[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3477_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n23754), .I0(GND_net), .I1(n1_adj_4608[9]), 
            .CO(n23755));
    SB_CARRY add_3477_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n24697));
    SB_LUT4 i2_4_lut_adj_1475 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_4459));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut_adj_1475.LUT_INIT = 16'h9c50;
    SB_LUT4 add_3476_9_lut (.I0(GND_net), .I1(n7900[6]), .I2(n630), .I3(n24696), 
            .O(n7890[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[8]), 
            .I3(n23753), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n23753), .I0(GND_net), .I1(n1_adj_4608[8]), 
            .CO(n23754));
    SB_LUT4 add_3476_8_lut (.I0(GND_net), .I1(n7900[5]), .I2(n557), .I3(n24695), 
            .O(n7890[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3476_8 (.CI(n24695), .I0(n7900[5]), .I1(n557), .CO(n24696));
    SB_LUT4 i18802_4_lut (.I0(n7924[2]), .I1(\Ki[4] ), .I2(n6_adj_4455), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_4460));   // verilog/motorControl.v(34[26:37])
    defparam i18802_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[7]), 
            .I3(n23752), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3476_7_lut (.I0(GND_net), .I1(n7900[4]), .I2(n484), .I3(n24694), 
            .O(n7890[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_11  (.CI(n23993), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n23994));
    SB_CARRY unary_minus_16_add_3_9 (.CI(n23752), .I0(GND_net), .I1(n1_adj_4608[7]), 
            .CO(n23753));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[6]), 
            .I3(n23751), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_4461));   // verilog/motorControl.v(34[26:37])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_3476_7 (.CI(n24694), .I0(n7900[4]), .I1(n484), .CO(n24695));
    SB_CARRY unary_minus_16_add_3_8 (.CI(n23751), .I0(GND_net), .I1(n1_adj_4608[6]), 
            .CO(n23752));
    SB_LUT4 add_3476_6_lut (.I0(GND_net), .I1(n7900[3]), .I2(n411), .I3(n24693), 
            .O(n7890[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18833_4_lut (.I0(n7930[1]), .I1(\Ki[3] ), .I2(n4_adj_4458), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_4462));   // verilog/motorControl.v(34[26:37])
    defparam i18833_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[5]), 
            .I3(n23750), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n23750), .I0(GND_net), .I1(n1_adj_4608[5]), 
            .CO(n23751));
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n23992), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[4]), 
            .I3(n23749), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3476_6 (.CI(n24693), .I0(n7900[3]), .I1(n411), .CO(n24694));
    SB_CARRY unary_minus_16_add_3_6 (.CI(n23749), .I0(GND_net), .I1(n1_adj_4608[4]), 
            .CO(n23750));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[3]), 
            .I3(n23748), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_10  (.CI(n23992), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n23993));
    SB_LUT4 i18868_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n23407));   // verilog/motorControl.v(34[26:37])
    defparam i18868_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n23748), .I0(GND_net), .I1(n1_adj_4608[3]), 
            .CO(n23749));
    SB_LUT4 add_3476_5_lut (.I0(GND_net), .I1(n7900[2]), .I2(n338), .I3(n24692), 
            .O(n7890[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3476_5 (.CI(n24692), .I0(n7900[2]), .I1(n338), .CO(n24693));
    SB_LUT4 i8_4_lut (.I0(n6_adj_4462), .I1(n11_adj_4461), .I2(n8_adj_4460), 
            .I3(n12_adj_4459), .O(n18_adj_4464));   // verilog/motorControl.v(34[26:37])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n23991), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3476_4_lut (.I0(GND_net), .I1(n7900[1]), .I2(n265_adj_4353), 
            .I3(n24691), .O(n7890[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[2]), 
            .I3(n23747), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18786_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n23305), .I3(n7924[0]), .O(n4_adj_4454));   // verilog/motorControl.v(34[26:37])
    defparam i18786_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_4465));   // verilog/motorControl.v(34[26:37])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n23747), .I0(GND_net), .I1(n1_adj_4608[2]), 
            .CO(n23748));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4608[1]), 
            .I3(n23746), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26003_4_lut (.I0(n31704), .I1(n31800), .I2(n35_adj_4379), 
            .I3(n31190), .O(n31836));   // verilog/motorControl.v(38[19:35])
    defparam i26003_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4465), .I1(n18_adj_4464), .I2(n23407), 
            .I3(n4_adj_4466), .O(n29321));   // verilog/motorControl.v(34[26:37])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18773_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n7917[0]));   // verilog/motorControl.v(34[26:37])
    defparam i18773_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i26004_3_lut (.I0(n31836), .I1(n257[18]), .I2(n37_adj_4410), 
            .I3(GND_net), .O(n31837));   // verilog/motorControl.v(38[19:35])
    defparam i26004_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3476_4 (.CI(n24691), .I0(n7900[1]), .I1(n265_adj_4353), 
            .CO(n24692));
    SB_LUT4 i18775_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n23305));   // verilog/motorControl.v(34[26:37])
    defparam i18775_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3476_3_lut (.I0(GND_net), .I1(n7900[0]), .I2(n192), .I3(n24690), 
            .O(n7890[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n23746), .I0(GND_net), .I1(n1_adj_4608[1]), 
            .CO(n23747));
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_9  (.CI(n23991), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n23992));
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[15]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3476_3 (.CI(n24690), .I0(n7900[0]), .I1(n192), .CO(n24691));
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[16]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3476_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n7890[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3476_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3476_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n24690));
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[17]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3475_10_lut (.I0(GND_net), .I1(n7890[7]), .I2(n700), .I3(n24689), 
            .O(n7879[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1_adj_4608[0]), 
            .I3(VCC_net), .O(n31081)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3475_9_lut (.I0(GND_net), .I1(n7890[6]), .I2(n627), .I3(n24688), 
            .O(n7879[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25986_3_lut (.I0(n31837), .I1(n257[19]), .I2(n39_adj_4468), 
            .I3(GND_net), .O(n31819));   // verilog/motorControl.v(38[19:35])
    defparam i25986_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4608[0]), 
            .CO(n23746));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[23]), 
            .I3(n23745), .O(\PID_CONTROLLER.integral_23__N_3627 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3475_9 (.CI(n24688), .I0(n7890[6]), .I1(n627), .CO(n24689));
    SB_LUT4 add_3475_8_lut (.I0(GND_net), .I1(n7890[5]), .I2(n554), .I3(n24687), 
            .O(n7879[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3475_8 (.CI(n24687), .I0(n7890[5]), .I1(n554), .CO(n24688));
    SB_LUT4 add_3475_7_lut (.I0(GND_net), .I1(n7890[4]), .I2(n481), .I3(n24686), 
            .O(n7879[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3475_7 (.CI(n24686), .I0(n7890[4]), .I1(n481), .CO(n24687));
    SB_LUT4 add_3475_6_lut (.I0(GND_net), .I1(n7890[3]), .I2(n408), .I3(n24685), 
            .O(n7879[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n23990), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i25351_4_lut (.I0(n43_adj_4420), .I1(n41_adj_4470), .I2(n39_adj_4468), 
            .I3(n31786), .O(n31182));
    defparam i25351_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3475_6 (.CI(n24685), .I0(n7890[3]), .I1(n408), .CO(n24686));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4607[22]), .I3(n23744), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_8  (.CI(n23990), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n23991));
    SB_CARRY unary_minus_5_add_3_24 (.CI(n23744), .I0(GND_net), .I1(n1_adj_4607[22]), 
            .CO(n23745));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4607[21]), .I3(n23743), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n23743), .I0(GND_net), .I1(n1_adj_4607[21]), 
            .CO(n23744));
    SB_LUT4 i25927_4_lut (.I0(n31702), .I1(n31631), .I2(n45_adj_4433), 
            .I3(n31180), .O(n31760));   // verilog/motorControl.v(38[19:35])
    defparam i25927_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4607[20]), .I3(n23742), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n23989), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n23742), .I0(GND_net), .I1(n1_adj_4607[20]), 
            .CO(n23743));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4607[19]), .I3(n23741), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n23741), .I0(GND_net), .I1(n1_adj_4607[19]), 
            .CO(n23742));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4607[18]), .I3(n23740), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_7  (.CI(n23989), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n23990));
    SB_CARRY unary_minus_5_add_3_20 (.CI(n23740), .I0(GND_net), .I1(n1_adj_4607[18]), 
            .CO(n23741));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4607[17]), .I3(n23739), .O(n35_adj_4259)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18856_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n23382), .I3(n7935[0]), .O(n4_adj_4466));   // verilog/motorControl.v(34[26:37])
    defparam i18856_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n23739), .I0(GND_net), .I1(n1_adj_4607[17]), 
            .CO(n23740));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4607[16]), .I3(n23738), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3475_5_lut (.I0(GND_net), .I1(n7890[2]), .I2(n335), .I3(n24684), 
            .O(n7879[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25980_3_lut (.I0(n31819), .I1(n257[20]), .I2(n41_adj_4470), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(38[19:35])
    defparam i25980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1476 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n7935[0]), .I3(n23382), .O(n7930[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1476.LUT_INIT = 16'h8778;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n23988), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n23738), .I0(GND_net), .I1(n1_adj_4607[16]), 
            .CO(n23739));
    SB_CARRY add_3475_5 (.CI(n24684), .I0(n7890[2]), .I1(n335), .CO(n24685));
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[18]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[5]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3475_4_lut (.I0(GND_net), .I1(n7890[1]), .I2(n262), .I3(n24683), 
            .O(n7879[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4607[15]), .I3(n23737), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3475_4 (.CI(n24683), .I0(n7890[1]), .I1(n262), .CO(n24684));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n23737), .I0(GND_net), .I1(n1_adj_4607[15]), 
            .CO(n23738));
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[19]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3475_3_lut (.I0(GND_net), .I1(n7890[0]), .I2(n189), .I3(n24682), 
            .O(n7879[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3475_3 (.CI(n24682), .I0(n7890[0]), .I1(n189), .CO(n24683));
    SB_LUT4 add_3475_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n7879[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3475_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4607[14]), .I3(n23736), .O(n29_adj_4258)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_6  (.CI(n23988), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n23989));
    SB_CARRY unary_minus_5_add_3_16 (.CI(n23736), .I0(GND_net), .I1(n1_adj_4607[14]), 
            .CO(n23737));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4607[13]), .I3(n23735), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n23735), .I0(GND_net), .I1(n1_adj_4607[13]), 
            .CO(n23736));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4607[12]), .I3(n23734), .O(n25_adj_4256)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26104_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31935));   // verilog/motorControl.v(29[14] 48[8])
    defparam i26104_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n23987), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n23734), .I0(GND_net), .I1(n1_adj_4607[12]), 
            .CO(n23735));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4607[11]), .I3(n23733), .O(n23_adj_4257)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3475_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n24682));
    SB_CARRY unary_minus_5_add_3_13 (.CI(n23733), .I0(GND_net), .I1(n1_adj_4607[11]), 
            .CO(n23734));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4607[10]), .I3(n23732), .O(n21_adj_4247)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_5  (.CI(n23987), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n23988));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n23732), .I0(GND_net), .I1(n1_adj_4607[10]), 
            .CO(n23733));
    SB_LUT4 i2_3_lut_4_lut_adj_1477 (.I0(n62), .I1(n131), .I2(n7930[0]), 
            .I3(n204), .O(n7924[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1477.LUT_INIT = 16'h8778;
    SB_LUT4 add_3474_11_lut (.I0(GND_net), .I1(n7879[8]), .I2(n770), .I3(n24681), 
            .O(n7867[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4607[9]), .I3(n23731), .O(n19_adj_4248)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3474_10_lut (.I0(GND_net), .I1(n7879[7]), .I2(n697), .I3(n24680), 
            .O(n7867[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n23731), .I0(GND_net), .I1(n1_adj_4607[9]), 
            .CO(n23732));
    SB_CARRY add_3474_10 (.CI(n24680), .I0(n7879[7]), .I1(n697), .CO(n24681));
    SB_LUT4 add_3474_9_lut (.I0(GND_net), .I1(n7879[6]), .I2(n624), .I3(n24679), 
            .O(n7867[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18825_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n7930[0]), 
            .O(n4_adj_4458));   // verilog/motorControl.v(34[26:37])
    defparam i18825_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4607[8]), .I3(n23730), .O(n17_adj_4249)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25929_4_lut (.I0(n40), .I1(n31760), .I2(n45_adj_4433), .I3(n31182), 
            .O(n31762));   // verilog/motorControl.v(38[19:35])
    defparam i25929_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3474_9 (.CI(n24679), .I0(n7879[6]), .I1(n624), .CO(n24680));
    SB_LUT4 add_3474_8_lut (.I0(GND_net), .I1(n7879[5]), .I2(n551), .I3(n24678), 
            .O(n7867[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3474_8 (.CI(n24678), .I0(n7879[5]), .I1(n551), .CO(n24679));
    SB_LUT4 add_3445_12_lut (.I0(GND_net), .I1(n7477[9]), .I2(n822_adj_4333), 
            .I3(n24348), .O(n7458[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3474_7_lut (.I0(GND_net), .I1(n7879[4]), .I2(n478), .I3(n24677), 
            .O(n7867[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[20]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3441_12 (.CI(n24274), .I0(n7395[9]), .I1(n810), .CO(n24275));
    SB_LUT4 i18845_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n23382));   // verilog/motorControl.v(34[26:37])
    defparam i18845_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_3474_7 (.CI(n24677), .I0(n7879[4]), .I1(n478), .CO(n24678));
    SB_LUT4 i25930_3_lut (.I0(n31762), .I1(duty[23]), .I2(n47_adj_4416), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(38[19:35])
    defparam i25930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3474_6_lut (.I0(GND_net), .I1(n7879[3]), .I2(n405), .I3(n24676), 
            .O(n7867[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[21]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n23730), .I0(GND_net), .I1(n1_adj_4607[8]), 
            .CO(n23731));
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n23986), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4607[7]), .I3(n23729), .O(n15_adj_4243)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n23729), .I0(GND_net), .I1(n1_adj_4607[7]), 
            .CO(n23730));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4607[6]), .I3(n23728), .O(n13_adj_4244)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3474_6 (.CI(n24676), .I0(n7879[3]), .I1(n405), .CO(n24677));
    SB_LUT4 i18843_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n7930[0]));   // verilog/motorControl.v(34[26:37])
    defparam i18843_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_3474_5_lut (.I0(GND_net), .I1(n7879[2]), .I2(n332), .I3(n24675), 
            .O(n7867[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n23728), .I0(GND_net), .I1(n1_adj_4607[6]), 
            .CO(n23729));
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_4  (.CI(n23986), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n23987));
    SB_CARRY add_3474_5 (.CI(n24675), .I0(n7879[2]), .I1(n332), .CO(n24676));
    SB_LUT4 add_3474_4_lut (.I0(GND_net), .I1(n7879[1]), .I2(n259), .I3(n24674), 
            .O(n7867[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4432));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_607_i1_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256), .I3(\Ki[0] ), .O(n2926[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_CARRY add_3474_4 (.CI(n24674), .I0(n7879[1]), .I1(n259), .CO(n24675));
    SB_LUT4 add_3474_3_lut (.I0(GND_net), .I1(n7879[0]), .I2(n186), .I3(n24673), 
            .O(n7867[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n23985), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4607[5]), .I3(n23727), .O(n11_adj_4245)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_3  (.CI(n23985), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n23986));
    SB_CARRY add_3474_3 (.CI(n24673), .I0(n7879[0]), .I1(n186), .CO(n24674));
    SB_LUT4 add_3474_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n7867[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3474_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3474_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n24673));
    SB_LUT4 add_3473_12_lut (.I0(GND_net), .I1(n7867[9]), .I2(n840), .I3(n24672), 
            .O(n7854[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3473_11_lut (.I0(GND_net), .I1(n7867[8]), .I2(n767), .I3(n24671), 
            .O(n7854[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_11 (.CI(n24671), .I0(n7867[8]), .I1(n767), .CO(n24672));
    SB_LUT4 add_3473_10_lut (.I0(GND_net), .I1(n7867[7]), .I2(n694), .I3(n24670), 
            .O(n7854[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_10 (.CI(n24670), .I0(n7867[7]), .I1(n694), .CO(n24671));
    SB_LUT4 add_3473_9_lut (.I0(GND_net), .I1(n7867[6]), .I2(n621), .I3(n24669), 
            .O(n7854[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_9 (.CI(n24669), .I0(n7867[6]), .I1(n621), .CO(n24670));
    SB_LUT4 add_3473_8_lut (.I0(GND_net), .I1(n7867[5]), .I2(n548), .I3(n24668), 
            .O(n7854[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_8 (.CI(n24668), .I0(n7867[5]), .I1(n548), .CO(n24669));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n23727), .I0(GND_net), .I1(n1_adj_4607[5]), 
            .CO(n23728));
    SB_LUT4 i14665_3_lut (.I0(\Kp[0] ), .I1(n256), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n2901[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam i14665_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mux_607_i2_3_lut (.I0(n155[1]), .I1(PWMLimit[1]), .I2(n256), 
            .I3(GND_net), .O(n2926[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3473_7_lut (.I0(GND_net), .I1(n7867[4]), .I2(n475), .I3(n24667), 
            .O(n7854[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_12 (.CI(n24348), .I0(n7477[9]), .I1(n822_adj_4333), 
            .CO(n24349));
    SB_LUT4 \PID_CONTROLLER.integral_1193_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1193_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_7 (.CI(n24667), .I0(n7867[4]), .I1(n475), .CO(n24668));
    SB_LUT4 add_3473_6_lut (.I0(GND_net), .I1(n7867[3]), .I2(n402), .I3(n24666), 
            .O(n7854[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1193_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n23985));
    SB_CARRY add_3473_6 (.CI(n24666), .I0(n7867[3]), .I1(n402), .CO(n24667));
    SB_LUT4 add_3473_5_lut (.I0(GND_net), .I1(n7867[2]), .I2(n329), .I3(n24665), 
            .O(n7854[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_5 (.CI(n24665), .I0(n7867[2]), .I1(n329), .CO(n24666));
    SB_LUT4 add_3473_4_lut (.I0(GND_net), .I1(n7867[1]), .I2(n256_adj_4327), 
            .I3(n24664), .O(n7854[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_607_i24_3_lut (.I0(n31114), .I1(PWMLimit[23]), .I2(n256), 
            .I3(GND_net), .O(n2926[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3473_4 (.CI(n24664), .I0(n7867[1]), .I1(n256_adj_4327), 
            .CO(n24665));
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[22]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14893_2_lut (.I0(n5790[0]), .I1(n256), .I2(GND_net), .I3(GND_net), 
            .O(n2901[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam i14893_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4422));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_607_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256), 
            .I3(GND_net), .O(n2926[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4608[23]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_607_i4_3_lut (.I0(n155[3]), .I1(PWMLimit[3]), .I2(n256), 
            .I3(GND_net), .O(n2926[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i4_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_607_i5_3_lut (.I0(n155[4]), .I1(PWMLimit[4]), .I2(n256), 
            .I3(GND_net), .O(n2926[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i5_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_607_i6_3_lut (.I0(n155[5]), .I1(PWMLimit[5]), .I2(n256), 
            .I3(GND_net), .O(n2926[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i6_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_607_i7_3_lut (.I0(n155[6]), .I1(PWMLimit[6]), .I2(n256), 
            .I3(GND_net), .O(n2926[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_607_i8_3_lut (.I0(n155[7]), .I1(PWMLimit[7]), .I2(n256), 
            .I3(GND_net), .O(n2926[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_607_i9_3_lut (.I0(n155[8]), .I1(PWMLimit[8]), .I2(n256), 
            .I3(GND_net), .O(n2926[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_607_i10_3_lut (.I0(n155[9]), .I1(PWMLimit[9]), .I2(n256), 
            .I3(GND_net), .O(n2926[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4411));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_607_i11_3_lut (.I0(n155[10]), .I1(PWMLimit[10]), .I2(n256), 
            .I3(GND_net), .O(n2926[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3473_3_lut (.I0(GND_net), .I1(n7867[0]), .I2(n183), .I3(n24663), 
            .O(n7854[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_3 (.CI(n24663), .I0(n7867[0]), .I1(n183), .CO(n24664));
    SB_LUT4 add_3473_2_lut (.I0(GND_net), .I1(n41_adj_4326), .I2(n110), 
            .I3(GND_net), .O(n7854[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_2 (.CI(GND_net), .I0(n41_adj_4326), .I1(n110), .CO(n24663));
    SB_LUT4 add_3472_13_lut (.I0(GND_net), .I1(n7854[10]), .I2(n910), 
            .I3(n24662), .O(n7840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3472_12_lut (.I0(GND_net), .I1(n7854[9]), .I2(n837), .I3(n24661), 
            .O(n7840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_12 (.CI(n24661), .I0(n7854[9]), .I1(n837), .CO(n24662));
    SB_LUT4 add_3472_11_lut (.I0(GND_net), .I1(n7854[8]), .I2(n764), .I3(n24660), 
            .O(n7840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_11 (.CI(n24660), .I0(n7854[8]), .I1(n764), .CO(n24661));
    SB_LUT4 add_3472_10_lut (.I0(GND_net), .I1(n7854[7]), .I2(n691), .I3(n24659), 
            .O(n7840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_10 (.CI(n24659), .I0(n7854[7]), .I1(n691), .CO(n24660));
    SB_LUT4 add_3472_9_lut (.I0(GND_net), .I1(n7854[6]), .I2(n618), .I3(n24658), 
            .O(n7840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4607[4]), .I3(n23726), .O(n9_adj_4250)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3472_9 (.CI(n24658), .I0(n7854[6]), .I1(n618), .CO(n24659));
    SB_LUT4 mux_607_i12_3_lut (.I0(n155[11]), .I1(PWMLimit[11]), .I2(n256), 
            .I3(GND_net), .O(n2926[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3472_8_lut (.I0(GND_net), .I1(n7854[5]), .I2(n545), .I3(n24657), 
            .O(n7840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_8 (.CI(n24657), .I0(n7854[5]), .I1(n545), .CO(n24658));
    SB_LUT4 mux_607_i13_3_lut (.I0(n155[12]), .I1(PWMLimit[12]), .I2(n256), 
            .I3(GND_net), .O(n2926[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3472_7_lut (.I0(GND_net), .I1(n7854[4]), .I2(n472), .I3(n24656), 
            .O(n7840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_7 (.CI(n24656), .I0(n7854[4]), .I1(n472), .CO(n24657));
    SB_LUT4 add_3472_6_lut (.I0(GND_net), .I1(n7854[3]), .I2(n399), .I3(n24655), 
            .O(n7840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_6 (.CI(n24655), .I0(n7854[3]), .I1(n399), .CO(n24656));
    SB_LUT4 add_3472_5_lut (.I0(GND_net), .I1(n7854[2]), .I2(n326), .I3(n24654), 
            .O(n7840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_5 (.CI(n24654), .I0(n7854[2]), .I1(n326), .CO(n24655));
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4476));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3441_11_lut (.I0(GND_net), .I1(n7395[8]), .I2(n737), .I3(n24273), 
            .O(n7372[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_11 (.CI(n24273), .I0(n7395[8]), .I1(n737), .CO(n24274));
    SB_LUT4 add_3472_4_lut (.I0(GND_net), .I1(n7854[1]), .I2(n253), .I3(n24653), 
            .O(n7840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_4 (.CI(n24653), .I0(n7854[1]), .I1(n253), .CO(n24654));
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4477));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3445_11_lut (.I0(GND_net), .I1(n7477[8]), .I2(n749_adj_4324), 
            .I3(n24347), .O(n7458[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4478));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4479));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4480));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4481));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4482));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4483));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4484));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4485));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4486));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4487));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4488));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3445_11 (.CI(n24347), .I0(n7477[8]), .I1(n749_adj_4324), 
            .CO(n24348));
    SB_LUT4 add_3445_10_lut (.I0(GND_net), .I1(n7477[7]), .I2(n676_adj_4323), 
            .I3(n24346), .O(n7458[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_10 (.CI(n24346), .I0(n7477[7]), .I1(n676_adj_4323), 
            .CO(n24347));
    SB_LUT4 add_3445_9_lut (.I0(GND_net), .I1(n7477[6]), .I2(n603_adj_4322), 
            .I3(n24345), .O(n7458[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_9 (.CI(n24345), .I0(n7477[6]), .I1(n603_adj_4322), 
            .CO(n24346));
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4489));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4490));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4491));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4492));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3472_3_lut (.I0(GND_net), .I1(n7854[0]), .I2(n180), .I3(n24652), 
            .O(n7840[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3445_8_lut (.I0(GND_net), .I1(n7477[5]), .I2(n530_adj_4321), 
            .I3(n24344), .O(n7458[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_8 (.CI(n24344), .I0(n7477[5]), .I1(n530_adj_4321), 
            .CO(n24345));
    SB_LUT4 add_3445_7_lut (.I0(GND_net), .I1(n7477[4]), .I2(n457_adj_4320), 
            .I3(n24343), .O(n7458[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_10_lut (.I0(GND_net), .I1(n7395[7]), .I2(n664), .I3(n24272), 
            .O(n7372[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_10 (.CI(n24272), .I0(n7395[7]), .I1(n664), .CO(n24273));
    SB_CARRY add_3445_7 (.CI(n24343), .I0(n7477[4]), .I1(n457_adj_4320), 
            .CO(n24344));
    SB_LUT4 add_3445_6_lut (.I0(GND_net), .I1(n7477[3]), .I2(n384_adj_4319), 
            .I3(n24342), .O(n7458[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_6 (.CI(n24342), .I0(n7477[3]), .I1(n384_adj_4319), 
            .CO(n24343));
    SB_LUT4 add_3445_5_lut (.I0(GND_net), .I1(n7477[2]), .I2(n311_adj_4318), 
            .I3(n24341), .O(n7458[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_5 (.CI(n24341), .I0(n7477[2]), .I1(n311_adj_4318), 
            .CO(n24342));
    SB_LUT4 add_3445_4_lut (.I0(GND_net), .I1(n7477[1]), .I2(n238_adj_4317), 
            .I3(n24340), .O(n7458[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n23726), .I0(GND_net), .I1(n1_adj_4607[4]), 
            .CO(n23727));
    SB_CARRY add_3472_3 (.CI(n24652), .I0(n7854[0]), .I1(n180), .CO(n24653));
    SB_LUT4 add_3472_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_4316), 
            .I3(GND_net), .O(n7840[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3472_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3472_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_4316), .CO(n24652));
    SB_LUT4 add_3471_14_lut (.I0(GND_net), .I1(n7840[11]), .I2(n980), 
            .I3(n24651), .O(n7825[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_13_lut (.I0(GND_net), .I1(n7840[10]), .I2(n907), 
            .I3(n24650), .O(n7825[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_13 (.CI(n24650), .I0(n7840[10]), .I1(n907), .CO(n24651));
    SB_LUT4 add_3471_12_lut (.I0(GND_net), .I1(n7840[9]), .I2(n834), .I3(n24649), 
            .O(n7825[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_12 (.CI(n24649), .I0(n7840[9]), .I1(n834), .CO(n24650));
    SB_LUT4 add_3471_11_lut (.I0(GND_net), .I1(n7840[8]), .I2(n761), .I3(n24648), 
            .O(n7825[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_11 (.CI(n24648), .I0(n7840[8]), .I1(n761), .CO(n24649));
    SB_LUT4 add_3471_10_lut (.I0(GND_net), .I1(n7840[7]), .I2(n688_adj_4315), 
            .I3(n24647), .O(n7825[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_10 (.CI(n24647), .I0(n7840[7]), .I1(n688_adj_4315), 
            .CO(n24648));
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3471_9_lut (.I0(GND_net), .I1(n7840[6]), .I2(n615_adj_4314), 
            .I3(n24646), .O(n7825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_9 (.CI(n24646), .I0(n7840[6]), .I1(n615_adj_4314), 
            .CO(n24647));
    SB_LUT4 add_3471_8_lut (.I0(GND_net), .I1(n7840[5]), .I2(n542_adj_4313), 
            .I3(n24645), .O(n7825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_8 (.CI(n24645), .I0(n7840[5]), .I1(n542_adj_4313), 
            .CO(n24646));
    SB_LUT4 add_3471_7_lut (.I0(GND_net), .I1(n7840[4]), .I2(n469_adj_4312), 
            .I3(n24644), .O(n7825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_7 (.CI(n24644), .I0(n7840[4]), .I1(n469_adj_4312), 
            .CO(n24645));
    SB_LUT4 add_3471_6_lut (.I0(GND_net), .I1(n7840[3]), .I2(n396_adj_4311), 
            .I3(n24643), .O(n7825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_6 (.CI(n24643), .I0(n7840[3]), .I1(n396_adj_4311), 
            .CO(n24644));
    SB_LUT4 add_3471_5_lut (.I0(GND_net), .I1(n7840[2]), .I2(n323_adj_4310), 
            .I3(n24642), .O(n7825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4493));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3441_9_lut (.I0(GND_net), .I1(n7395[6]), .I2(n591), .I3(n24271), 
            .O(n7372[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_4 (.CI(n24340), .I0(n7477[1]), .I1(n238_adj_4317), 
            .CO(n24341));
    SB_CARRY add_3441_9 (.CI(n24271), .I0(n7395[6]), .I1(n591), .CO(n24272));
    SB_LUT4 add_3445_3_lut (.I0(GND_net), .I1(n7477[0]), .I2(n165_adj_4309), 
            .I3(n24339), .O(n7458[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4494));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3445_3 (.CI(n24339), .I0(n7477[0]), .I1(n165_adj_4309), 
            .CO(n24340));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4607[3]), .I3(n23725), .O(n7_adj_4254)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n23725), .I0(GND_net), .I1(n1_adj_4607[3]), 
            .CO(n23726));
    SB_LUT4 add_3445_2_lut (.I0(GND_net), .I1(n23_adj_4307), .I2(n92_adj_4306), 
            .I3(GND_net), .O(n7458[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4607[2]), .I3(n23724), .O(n5_adj_4255)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25408_4_lut (.I0(n21_adj_4494), .I1(n19_adj_4493), .I2(n17_adj_4492), 
            .I3(n9_adj_4491), .O(n31239));
    defparam i25408_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3471_5 (.CI(n24642), .I0(n7840[2]), .I1(n323_adj_4310), 
            .CO(n24643));
    SB_LUT4 i25399_4_lut (.I0(n27_adj_4490), .I1(n15_adj_4489), .I2(n13_adj_4488), 
            .I3(n11_adj_4487), .O(n31230));
    defparam i25399_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3441_8_lut (.I0(GND_net), .I1(n7395[5]), .I2(n518), .I3(n24270), 
            .O(n7372[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_8 (.CI(n24270), .I0(n7395[5]), .I1(n518), .CO(n24271));
    SB_LUT4 add_3441_7_lut (.I0(GND_net), .I1(n7395[4]), .I2(n445), .I3(n24269), 
            .O(n7372[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_7 (.CI(n24269), .I0(n7395[4]), .I1(n445), .CO(n24270));
    SB_LUT4 add_3441_6_lut (.I0(GND_net), .I1(n7395[3]), .I2(n372), .I3(n24268), 
            .O(n7372[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_6 (.CI(n24268), .I0(n7395[3]), .I1(n372), .CO(n24269));
    SB_CARRY add_3445_2 (.CI(GND_net), .I0(n23_adj_4307), .I1(n92_adj_4306), 
            .CO(n24339));
    SB_LUT4 add_3441_5_lut (.I0(GND_net), .I1(n7395[2]), .I2(n299), .I3(n24267), 
            .O(n7372[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n23724), .I0(GND_net), .I1(n1_adj_4607[2]), 
            .CO(n23725));
    SB_LUT4 add_3444_19_lut (.I0(GND_net), .I1(n7458[16]), .I2(GND_net), 
            .I3(n24338), .O(n7438[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4607[1]), .I3(n23723), .O(n3_adj_4268)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3441_5 (.CI(n24267), .I0(n7395[2]), .I1(n299), .CO(n24268));
    SB_LUT4 add_3471_4_lut (.I0(GND_net), .I1(n7840[1]), .I2(n250_adj_4303), 
            .I3(n24641), .O(n7825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n23723), .I0(GND_net), .I1(n1_adj_4607[1]), 
            .CO(n23724));
    SB_LUT4 add_3444_18_lut (.I0(GND_net), .I1(n7458[15]), .I2(GND_net), 
            .I3(n24337), .O(n7438[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_4 (.CI(n24641), .I0(n7840[1]), .I1(n250_adj_4303), 
            .CO(n24642));
    SB_CARRY add_3444_18 (.CI(n24337), .I0(n7458[15]), .I1(GND_net), .CO(n24338));
    SB_LUT4 add_3441_4_lut (.I0(GND_net), .I1(n7395[1]), .I2(n226), .I3(n24266), 
            .O(n7372[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12_adj_4495), .I1(duty[17]), .I2(n35_adj_4485), 
            .I3(GND_net), .O(n30_adj_4496));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3471_3_lut (.I0(GND_net), .I1(n7840[0]), .I2(n177_adj_4302), 
            .I3(n24640), .O(n7825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_3 (.CI(n24640), .I0(n7840[0]), .I1(n177_adj_4302), 
            .CO(n24641));
    SB_LUT4 add_3444_17_lut (.I0(GND_net), .I1(n7458[14]), .I2(GND_net), 
            .I3(n24336), .O(n7438[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25667_4_lut (.I0(n13_adj_4488), .I1(n11_adj_4487), .I2(n9_adj_4491), 
            .I3(n31249), .O(n31500));
    defparam i25667_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_3441_4 (.CI(n24266), .I0(n7395[1]), .I1(n226), .CO(n24267));
    SB_LUT4 add_3441_3_lut (.I0(GND_net), .I1(n7395[0]), .I2(n153), .I3(n24265), 
            .O(n7372[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3444_17 (.CI(n24336), .I0(n7458[14]), .I1(GND_net), .CO(n24337));
    SB_LUT4 add_3444_16_lut (.I0(GND_net), .I1(n7458[13]), .I2(n1111_adj_4301), 
            .I3(n24335), .O(n7438[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_3 (.CI(n24265), .I0(n7395[0]), .I1(n153), .CO(n24266));
    SB_LUT4 i25663_4_lut (.I0(n19_adj_4493), .I1(n17_adj_4492), .I2(n15_adj_4489), 
            .I3(n31500), .O(n31496));
    defparam i25663_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_3441_2_lut (.I0(GND_net), .I1(n11_adj_4300), .I2(n80), 
            .I3(GND_net), .O(n7372[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_2 (.CI(GND_net), .I0(n11_adj_4300), .I1(n80), .CO(n24265));
    SB_LUT4 i25931_4_lut (.I0(n25_adj_4484), .I1(n23_adj_4483), .I2(n21_adj_4494), 
            .I3(n31496), .O(n31764));
    defparam i25931_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25790_4_lut (.I0(n31_adj_4482), .I1(n29_adj_4481), .I2(n27_adj_4490), 
            .I3(n31764), .O(n31623));
    defparam i25790_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n7348[21]), 
            .I2(GND_net), .I3(n24264), .O(n5790[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3444_16 (.CI(n24335), .I0(n7458[13]), .I1(n1111_adj_4301), 
            .CO(n24336));
    SB_LUT4 i25955_4_lut (.I0(n37_adj_4480), .I1(n35_adj_4485), .I2(n33_adj_4486), 
            .I3(n31623), .O(n31788));
    defparam i25955_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n19402), .I1(n7348[20]), .I2(GND_net), 
            .I3(n24263), .O(n2901[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_23 (.CI(n24263), .I0(n7348[20]), .I1(GND_net), 
            .CO(n24264));
    SB_LUT4 add_3444_15_lut (.I0(GND_net), .I1(n7458[12]), .I2(n1038_adj_4299), 
            .I3(n24334), .O(n7438[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3444_15 (.CI(n24334), .I0(n7458[12]), .I1(n1038_adj_4299), 
            .CO(n24335));
    SB_LUT4 add_3471_2_lut (.I0(GND_net), .I1(n35_adj_4298), .I2(n104_adj_4297), 
            .I3(GND_net), .O(n7825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n19402), .I1(n7348[19]), .I2(GND_net), 
            .I3(n24262), .O(n2901[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i25842_3_lut (.I0(n6_adj_4497), .I1(duty[10]), .I2(n21_adj_4494), 
            .I3(GND_net), .O(n31675));   // verilog/motorControl.v(36[10:25])
    defparam i25842_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3471_2 (.CI(GND_net), .I0(n35_adj_4298), .I1(n104_adj_4297), 
            .CO(n24640));
    SB_LUT4 i25843_3_lut (.I0(n31675), .I1(duty[11]), .I2(n23_adj_4483), 
            .I3(GND_net), .O(n31676));   // verilog/motorControl.v(36[10:25])
    defparam i25843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3444_14_lut (.I0(GND_net), .I1(n7458[11]), .I2(n965_adj_4296), 
            .I3(n24333), .O(n7438[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16_adj_4498), .I1(duty[22]), .I2(n45_adj_4478), 
            .I3(GND_net), .O(n24_adj_4499));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_10_add_1225_22 (.CI(n24262), .I0(n7348[19]), .I1(GND_net), 
            .CO(n24263));
    SB_CARRY add_3444_14 (.CI(n24333), .I0(n7458[11]), .I1(n965_adj_4296), 
            .CO(n24334));
    SB_LUT4 add_3470_15_lut (.I0(GND_net), .I1(n7825[12]), .I2(n1050_adj_4295), 
            .I3(n24639), .O(n7809[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3470_14_lut (.I0(GND_net), .I1(n7825[11]), .I2(n977_adj_4294), 
            .I3(n24638), .O(n7809[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_14 (.CI(n24638), .I0(n7825[11]), .I1(n977_adj_4294), 
            .CO(n24639));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n19402), .I1(n7348[18]), .I2(GND_net), 
            .I3(n24261), .O(n2901[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3444_13_lut (.I0(GND_net), .I1(n7458[10]), .I2(n892_adj_4293), 
            .I3(n24332), .O(n7438[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3444_13 (.CI(n24332), .I0(n7458[10]), .I1(n892_adj_4293), 
            .CO(n24333));
    SB_LUT4 add_3470_13_lut (.I0(GND_net), .I1(n7825[10]), .I2(n904_adj_4292), 
            .I3(n24637), .O(n7809[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3444_12_lut (.I0(GND_net), .I1(n7458[9]), .I2(n819_adj_4291), 
            .I3(n24331), .O(n7438[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3444_12 (.CI(n24331), .I0(n7458[9]), .I1(n819_adj_4291), 
            .CO(n24332));
    SB_CARRY add_3470_13 (.CI(n24637), .I0(n7825[10]), .I1(n904_adj_4292), 
            .CO(n24638));
    SB_LUT4 add_3444_11_lut (.I0(GND_net), .I1(n7458[8]), .I2(n746_adj_4290), 
            .I3(n24330), .O(n7438[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3470_12_lut (.I0(GND_net), .I1(n7825[9]), .I2(n831_adj_4289), 
            .I3(n24636), .O(n7809[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3627 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25383_4_lut (.I0(n43_adj_4479), .I1(n25_adj_4484), .I2(n23_adj_4483), 
            .I3(n31239), .O(n31214));
    defparam i25383_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3470_12 (.CI(n24636), .I0(n7825[9]), .I1(n831_adj_4289), 
            .CO(n24637));
    SB_LUT4 add_3470_11_lut (.I0(GND_net), .I1(n7825[8]), .I2(n758_adj_4287), 
            .I3(n24635), .O(n7809[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_11 (.CI(n24635), .I0(n7825[8]), .I1(n758_adj_4287), 
            .CO(n24636));
    SB_LUT4 add_3470_10_lut (.I0(GND_net), .I1(n7825[7]), .I2(n685_adj_4286), 
            .I3(n24634), .O(n7809[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_10 (.CI(n24634), .I0(n7825[7]), .I1(n685_adj_4286), 
            .CO(n24635));
    SB_LUT4 add_3470_9_lut (.I0(GND_net), .I1(n7825[6]), .I2(n612_adj_4285), 
            .I3(n24633), .O(n7809[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_9 (.CI(n24633), .I0(n7825[6]), .I1(n612_adj_4285), 
            .CO(n24634));
    SB_LUT4 add_3470_8_lut (.I0(GND_net), .I1(n7825[5]), .I2(n539_adj_4284), 
            .I3(n24632), .O(n7809[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25796_4_lut (.I0(n24_adj_4499), .I1(n8_adj_4500), .I2(n45_adj_4478), 
            .I3(n31212), .O(n31629));   // verilog/motorControl.v(36[10:25])
    defparam i25796_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3470_8 (.CI(n24632), .I0(n7825[5]), .I1(n539_adj_4284), 
            .CO(n24633));
    SB_LUT4 add_3470_7_lut (.I0(GND_net), .I1(n7825[4]), .I2(n466_adj_4283), 
            .I3(n24631), .O(n7809[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_7 (.CI(n24631), .I0(n7825[4]), .I1(n466_adj_4283), 
            .CO(n24632));
    SB_LUT4 add_3470_6_lut (.I0(GND_net), .I1(n7825[3]), .I2(n393_adj_4282), 
            .I3(n24630), .O(n7809[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_6 (.CI(n24630), .I0(n7825[3]), .I1(n393_adj_4282), 
            .CO(n24631));
    SB_DFFE \PID_CONTROLLER.integral_1193__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[0]));   // verilog/motorControl.v(32[21:33])
    SB_LUT4 i25654_3_lut (.I0(n31676), .I1(duty[12]), .I2(n25_adj_4484), 
            .I3(GND_net), .O(n31487));   // verilog/motorControl.v(36[10:25])
    defparam i25654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3470_5_lut (.I0(GND_net), .I1(n7825[2]), .I2(n320_adj_4235), 
            .I3(n24629), .O(n7809[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_5 (.CI(n24629), .I0(n7825[2]), .I1(n320_adj_4235), 
            .CO(n24630));
    SB_LUT4 add_3470_4_lut (.I0(GND_net), .I1(n7825[1]), .I2(n247_adj_4234), 
            .I3(n24628), .O(n7809[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_4501));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i25909_3_lut (.I0(n4_adj_4501), .I1(duty[13]), .I2(n27_adj_4490), 
            .I3(GND_net), .O(n31742));   // verilog/motorControl.v(36[10:25])
    defparam i25909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18734_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n23250), .I3(n7638[0]), .O(n4_adj_4502));   // verilog/motorControl.v(34[17:23])
    defparam i18734_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_3470_4 (.CI(n24628), .I0(n7825[1]), .I1(n247_adj_4234), 
            .CO(n24629));
    SB_LUT4 add_3470_3_lut (.I0(GND_net), .I1(n7825[0]), .I2(n174_adj_4233), 
            .I3(n24627), .O(n7809[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_3 (.CI(n24627), .I0(n7825[0]), .I1(n174_adj_4233), 
            .CO(n24628));
    SB_LUT4 add_3470_2_lut (.I0(GND_net), .I1(n32_adj_4231), .I2(n101_adj_4230), 
            .I3(GND_net), .O(n7809[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3470_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3470_2 (.CI(GND_net), .I0(n32_adj_4231), .I1(n101_adj_4230), 
            .CO(n24627));
    SB_LUT4 i2_3_lut_4_lut_adj_1478 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n7638[0]), .I3(n23250), .O(n7633[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1478.LUT_INIT = 16'h8778;
    SB_LUT4 add_3469_16_lut (.I0(GND_net), .I1(n7809[13]), .I2(n1120_adj_4229), 
            .I3(n24626), .O(n7792[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25910_3_lut (.I0(n31742), .I1(duty[14]), .I2(n29_adj_4481), 
            .I3(GND_net), .O(n31743));   // verilog/motorControl.v(36[10:25])
    defparam i25910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25394_4_lut (.I0(n33_adj_4486), .I1(n31_adj_4482), .I2(n29_adj_4481), 
            .I3(n31230), .O(n31225));
    defparam i25394_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3469_15_lut (.I0(GND_net), .I1(n7809[12]), .I2(n1047_adj_4228), 
            .I3(n24625), .O(n7792[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18723_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n23250));   // verilog/motorControl.v(34[17:23])
    defparam i18723_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i25965_4_lut (.I0(n30_adj_4496), .I1(n10_adj_4503), .I2(n35_adj_4485), 
            .I3(n31223), .O(n31798));   // verilog/motorControl.v(36[10:25])
    defparam i25965_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY mult_10_add_1225_21 (.CI(n24261), .I0(n7348[18]), .I1(GND_net), 
            .CO(n24262));
    SB_LUT4 i25865_3_lut (.I0(n31743), .I1(duty[15]), .I2(n31_adj_4482), 
            .I3(GND_net), .O(n31698));   // verilog/motorControl.v(36[10:25])
    defparam i25865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26001_4_lut (.I0(n31698), .I1(n31798), .I2(n35_adj_4485), 
            .I3(n31225), .O(n31834));   // verilog/motorControl.v(36[10:25])
    defparam i26001_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n19402), .I1(n7348[17]), .I2(GND_net), 
            .I3(n24260), .O(n2901[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3469_15 (.CI(n24625), .I0(n7809[12]), .I1(n1047_adj_4228), 
            .CO(n24626));
    SB_LUT4 add_3469_14_lut (.I0(GND_net), .I1(n7809[11]), .I2(n974_adj_4227), 
            .I3(n24624), .O(n7792[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26002_3_lut (.I0(n31834), .I1(duty[18]), .I2(n37_adj_4480), 
            .I3(GND_net), .O(n31835));   // verilog/motorControl.v(36[10:25])
    defparam i26002_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3469_14 (.CI(n24624), .I0(n7809[11]), .I1(n974_adj_4227), 
            .CO(n24625));
    SB_LUT4 i25988_3_lut (.I0(n31835), .I1(duty[19]), .I2(n39_adj_4477), 
            .I3(GND_net), .O(n31821));   // verilog/motorControl.v(36[10:25])
    defparam i25988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25385_4_lut (.I0(n43_adj_4479), .I1(n41_adj_4476), .I2(n39_adj_4477), 
            .I3(n31788), .O(n31216));
    defparam i25385_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i18721_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n7633[0]));   // verilog/motorControl.v(34[17:23])
    defparam i18721_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25921_4_lut (.I0(n31487), .I1(n31629), .I2(n45_adj_4478), 
            .I3(n31214), .O(n31754));   // verilog/motorControl.v(36[10:25])
    defparam i25921_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25978_3_lut (.I0(n31821), .I1(duty[20]), .I2(n41_adj_4476), 
            .I3(GND_net), .O(n40_adj_4504));   // verilog/motorControl.v(36[10:25])
    defparam i25978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25923_4_lut (.I0(n40_adj_4504), .I1(n31754), .I2(n45_adj_4478), 
            .I3(n31216), .O(n31756));   // verilog/motorControl.v(36[10:25])
    defparam i25923_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3444_11 (.CI(n24330), .I0(n7458[8]), .I1(n746_adj_4290), 
            .CO(n24331));
    SB_LUT4 add_3469_13_lut (.I0(GND_net), .I1(n7809[10]), .I2(n901_adj_4226), 
            .I3(n24623), .O(n7792[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n24260), .I0(n7348[17]), .I1(GND_net), 
            .CO(n24261));
    SB_CARRY add_3469_13 (.CI(n24623), .I0(n7809[10]), .I1(n901_adj_4226), 
            .CO(n24624));
    SB_LUT4 add_3469_12_lut (.I0(GND_net), .I1(n7809[9]), .I2(n828_adj_4225), 
            .I3(n24622), .O(n7792[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n19402), .I1(n7348[16]), .I2(GND_net), 
            .I3(n24259), .O(n2901[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3469_12 (.CI(n24622), .I0(n7809[9]), .I1(n828_adj_4225), 
            .CO(n24623));
    SB_LUT4 i25924_3_lut (.I0(n31756), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3675));   // verilog/motorControl.v(36[10:25])
    defparam i25924_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3469_11_lut (.I0(GND_net), .I1(n7809[8]), .I2(n755_adj_4224), 
            .I3(n24621), .O(n7792[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18703_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n23216), .I3(n7633[0]), .O(n4_adj_4505));   // verilog/motorControl.v(34[17:23])
    defparam i18703_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1479 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n7633[0]), .I3(n23216), .O(n7627[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1479.LUT_INIT = 16'h8778;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3651[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3675), .I3(GND_net), .O(duty_23__N_3528[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18690_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n7627[0]));   // verilog/motorControl.v(34[17:23])
    defparam i18690_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_3469_11 (.CI(n24621), .I0(n7809[8]), .I1(n755_adj_4224), 
            .CO(n24622));
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4607[0]), 
            .CO(n23723));
    SB_LUT4 add_3469_10_lut (.I0(GND_net), .I1(n7809[7]), .I2(n682_adj_4222), 
            .I3(n24620), .O(n7792[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18692_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n23216));   // verilog/motorControl.v(34[17:23])
    defparam i18692_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_3469_10 (.CI(n24620), .I0(n7809[7]), .I1(n682_adj_4222), 
            .CO(n24621));
    SB_LUT4 add_3444_10_lut (.I0(GND_net), .I1(n7458[7]), .I2(n673), .I3(n24329), 
            .O(n7438[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n24259), .I0(n7348[16]), .I1(GND_net), 
            .CO(n24260));
    SB_LUT4 add_3469_9_lut (.I0(GND_net), .I1(n7809[6]), .I2(n609_adj_4221), 
            .I3(n24619), .O(n7792[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18672_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_4506), .I3(n7627[1]), .O(n6_adj_4507));   // verilog/motorControl.v(34[17:23])
    defparam i18672_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1480 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n7627[1]), .I3(n4_adj_4506), .O(n7620[2]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1480.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n7627[0]), .I3(n23173), .O(n7620[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h8778;
    SB_LUT4 mux_607_i14_3_lut (.I0(n155[13]), .I1(PWMLimit[13]), .I2(n256), 
            .I3(GND_net), .O(n2926[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i14_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n19402), .I1(n7348[15]), .I2(GND_net), 
            .I3(n24258), .O(n2901[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3469_9 (.CI(n24619), .I0(n7809[6]), .I1(n609_adj_4221), 
            .CO(n24620));
    SB_LUT4 add_3469_8_lut (.I0(GND_net), .I1(n7809[5]), .I2(n536_adj_4220), 
            .I3(n24618), .O(n7792[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3469_8 (.CI(n24618), .I0(n7809[5]), .I1(n536_adj_4220), 
            .CO(n24619));
    SB_LUT4 add_3469_7_lut (.I0(GND_net), .I1(n7809[4]), .I2(n463_adj_4219), 
            .I3(n24617), .O(n7792[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18664_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n23173), .I3(n7627[0]), .O(n4_adj_4506));   // verilog/motorControl.v(34[17:23])
    defparam i18664_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY mult_10_add_1225_18 (.CI(n24258), .I0(n7348[15]), .I1(GND_net), 
            .CO(n24259));
    SB_CARRY add_3469_7 (.CI(n24617), .I0(n7809[4]), .I1(n463_adj_4219), 
            .CO(n24618));
    SB_LUT4 add_3469_6_lut (.I0(GND_net), .I1(n7809[3]), .I2(n390_adj_4217), 
            .I3(n24616), .O(n7792[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3469_6 (.CI(n24616), .I0(n7809[3]), .I1(n390_adj_4217), 
            .CO(n24617));
    SB_LUT4 add_3469_5_lut (.I0(GND_net), .I1(n7809[2]), .I2(n317_adj_4216), 
            .I3(n24615), .O(n7792[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18653_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n23173));   // verilog/motorControl.v(34[17:23])
    defparam i18653_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i18651_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n7620[0]));   // verilog/motorControl.v(34[17:23])
    defparam i18651_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_607_i15_3_lut (.I0(n155[14]), .I1(PWMLimit[14]), .I2(n256), 
            .I3(GND_net), .O(n2926[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_607_i16_3_lut (.I0(n155[15]), .I1(PWMLimit[15]), .I2(n256), 
            .I3(GND_net), .O(n2926[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3469_5 (.CI(n24615), .I0(n7809[2]), .I1(n317_adj_4216), 
            .CO(n24616));
    SB_LUT4 add_3469_4_lut (.I0(GND_net), .I1(n7809[1]), .I2(n244_adj_4214), 
            .I3(n24614), .O(n7792[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3469_4 (.CI(n24614), .I0(n7809[1]), .I1(n244_adj_4214), 
            .CO(n24615));
    SB_LUT4 add_3469_3_lut (.I0(GND_net), .I1(n7809[0]), .I2(n171_adj_4213), 
            .I3(n24613), .O(n7792[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3469_3 (.CI(n24613), .I0(n7809[0]), .I1(n171_adj_4213), 
            .CO(n24614));
    SB_LUT4 add_3469_2_lut (.I0(GND_net), .I1(n29_adj_4210), .I2(n98_adj_4209), 
            .I3(GND_net), .O(n7792[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3469_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3469_2 (.CI(GND_net), .I0(n29_adj_4210), .I1(n98_adj_4209), 
            .CO(n24613));
    SB_LUT4 add_3468_17_lut (.I0(GND_net), .I1(n7792[14]), .I2(GND_net), 
            .I3(n24612), .O(n7774[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3468_16_lut (.I0(GND_net), .I1(n7792[13]), .I2(n1117_adj_4207), 
            .I3(n24611), .O(n7774[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_16 (.CI(n24611), .I0(n7792[13]), .I1(n1117_adj_4207), 
            .CO(n24612));
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_607_i17_3_lut (.I0(n155[16]), .I1(PWMLimit[16]), .I2(n256), 
            .I3(GND_net), .O(n2926[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_607_i18_3_lut (.I0(n155[17]), .I1(PWMLimit[17]), .I2(n256), 
            .I3(GND_net), .O(n2926[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i18_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4193));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_607_i19_3_lut (.I0(n155[18]), .I1(PWMLimit[18]), .I2(n256), 
            .I3(GND_net), .O(n2926[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4192));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3444_10 (.CI(n24329), .I0(n7458[7]), .I1(n673), .CO(n24330));
    SB_LUT4 mux_607_i20_3_lut (.I0(n155[19]), .I1(PWMLimit[19]), .I2(n256), 
            .I3(GND_net), .O(n2926[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3468_15_lut (.I0(GND_net), .I1(n7792[12]), .I2(n1044_adj_4206), 
            .I3(n24610), .O(n7774[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_15 (.CI(n24610), .I0(n7792[12]), .I1(n1044_adj_4206), 
            .CO(n24611));
    SB_LUT4 mux_607_i21_3_lut (.I0(n155[20]), .I1(PWMLimit[20]), .I2(n256), 
            .I3(GND_net), .O(n2926[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25379_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n31210));   // verilog/motorControl.v(38[19:35])
    defparam i25379_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_607_i22_3_lut (.I0(n155[21]), .I1(PWMLimit[21]), .I2(n256), 
            .I3(GND_net), .O(n2926[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_4426));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mux_607_i23_3_lut (.I0(n155[22]), .I1(PWMLimit[22]), .I2(n256), 
            .I3(GND_net), .O(n2926[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_607_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4470));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4468));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4433));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4398));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4397));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4420));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4410));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4379));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4390));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4389));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3468_14_lut (.I0(GND_net), .I1(n7792[11]), .I2(n971_adj_4196), 
            .I3(n24609), .O(n7774[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_14 (.CI(n24609), .I0(n7792[11]), .I1(n971_adj_4196), 
            .CO(n24610));
    SB_LUT4 add_3468_13_lut (.I0(GND_net), .I1(n7792[10]), .I2(n898_adj_4195), 
            .I3(n24608), .O(n7774[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_13 (.CI(n24608), .I0(n7792[10]), .I1(n898_adj_4195), 
            .CO(n24609));
    SB_LUT4 add_3468_12_lut (.I0(GND_net), .I1(n7792[9]), .I2(n825), .I3(n24607), 
            .O(n7774[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_12 (.CI(n24607), .I0(n7792[9]), .I1(n825), .CO(n24608));
    SB_LUT4 add_3468_11_lut (.I0(GND_net), .I1(n7792[8]), .I2(n752), .I3(n24606), 
            .O(n7774[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_11 (.CI(n24606), .I0(n7792[8]), .I1(n752), .CO(n24607));
    SB_LUT4 add_3468_10_lut (.I0(GND_net), .I1(n7792[7]), .I2(n679), .I3(n24605), 
            .O(n7774[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_10 (.CI(n24605), .I0(n7792[7]), .I1(n679), .CO(n24606));
    SB_LUT4 add_3468_9_lut (.I0(GND_net), .I1(n7792[6]), .I2(n606), .I3(n24604), 
            .O(n7774[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_9 (.CI(n24604), .I0(n7792[6]), .I1(n606), .CO(n24605));
    SB_LUT4 add_3468_8_lut (.I0(GND_net), .I1(n7792[5]), .I2(n533), .I3(n24603), 
            .O(n7774[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_8 (.CI(n24603), .I0(n7792[5]), .I1(n533), .CO(n24604));
    SB_LUT4 add_3468_7_lut (.I0(GND_net), .I1(n7792[4]), .I2(n460), .I3(n24602), 
            .O(n7774[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_7 (.CI(n24602), .I0(n7792[4]), .I1(n460), .CO(n24603));
    SB_LUT4 add_3468_6_lut (.I0(GND_net), .I1(n7792[3]), .I2(n387), .I3(n24601), 
            .O(n7774[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_6 (.CI(n24601), .I0(n7792[3]), .I1(n387), .CO(n24602));
    SB_LUT4 add_3468_5_lut (.I0(GND_net), .I1(n7792[2]), .I2(n314), .I3(n24600), 
            .O(n7774[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_5 (.CI(n24600), .I0(n7792[2]), .I1(n314), .CO(n24601));
    SB_LUT4 add_3468_4_lut (.I0(GND_net), .I1(n7792[1]), .I2(n241), .I3(n24599), 
            .O(n7774[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3444_9_lut (.I0(GND_net), .I1(n7458[6]), .I2(n600), .I3(n24328), 
            .O(n7438[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_4 (.CI(n24599), .I0(n7792[1]), .I1(n241), .CO(n24600));
    SB_LUT4 add_3468_3_lut (.I0(GND_net), .I1(n7792[0]), .I2(n168), .I3(n24598), 
            .O(n7774[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_3 (.CI(n24598), .I0(n7792[0]), .I1(n168), .CO(n24599));
    SB_LUT4 add_3468_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n7774[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3468_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3468_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n24598));
    SB_LUT4 add_3467_18_lut (.I0(GND_net), .I1(n7774[15]), .I2(GND_net), 
            .I3(n24597), .O(n7755[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3467_17_lut (.I0(GND_net), .I1(n7774[14]), .I2(GND_net), 
            .I3(n24596), .O(n7755[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_17 (.CI(n24596), .I0(n7774[14]), .I1(GND_net), .CO(n24597));
    SB_CARRY add_3444_9 (.CI(n24328), .I0(n7458[6]), .I1(n600), .CO(n24329));
    SB_LUT4 add_3467_16_lut (.I0(GND_net), .I1(n7774[13]), .I2(n1114), 
            .I3(n24595), .O(n7755[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_16 (.CI(n24595), .I0(n7774[13]), .I1(n1114), .CO(n24596));
    SB_LUT4 add_3467_15_lut (.I0(GND_net), .I1(n7774[12]), .I2(n1041_adj_4186), 
            .I3(n24594), .O(n7755[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_15 (.CI(n24594), .I0(n7774[12]), .I1(n1041_adj_4186), 
            .CO(n24595));
    SB_LUT4 add_3467_14_lut (.I0(GND_net), .I1(n7774[11]), .I2(n968), 
            .I3(n24593), .O(n7755[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_14 (.CI(n24593), .I0(n7774[11]), .I1(n968), .CO(n24594));
    SB_LUT4 add_3467_13_lut (.I0(GND_net), .I1(n7774[10]), .I2(n895), 
            .I3(n24592), .O(n7755[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_13 (.CI(n24592), .I0(n7774[10]), .I1(n895), .CO(n24593));
    SB_LUT4 add_3467_12_lut (.I0(GND_net), .I1(n7774[9]), .I2(n822), .I3(n24591), 
            .O(n7755[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_4500));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25381_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n31212));
    defparam i25381_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16_adj_4498));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_4503));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25392_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n31223));
    defparam i25392_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12_adj_4495));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3467_12 (.CI(n24591), .I0(n7774[9]), .I1(n822), .CO(n24592));
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3528[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_3467_11_lut (.I0(GND_net), .I1(n7774[8]), .I2(n749), .I3(n24590), 
            .O(n7755[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_11 (.CI(n24590), .I0(n7774[8]), .I1(n749), .CO(n24591));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n19402), .I1(n7348[14]), .I2(GND_net), 
            .I3(n24257), .O(n2901[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_17 (.CI(n24257), .I0(n7348[14]), .I1(GND_net), 
            .CO(n24258));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n19402), .I1(n7348[13]), .I2(n1096), 
            .I3(n24256), .O(n2901[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_16 (.CI(n24256), .I0(n7348[13]), .I1(n1096), 
            .CO(n24257));
    SB_LUT4 add_3444_8_lut (.I0(GND_net), .I1(n7458[5]), .I2(n527_adj_4281), 
            .I3(n24327), .O(n7438[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n19402), .I1(n7348[12]), .I2(n1023), 
            .I3(n24255), .O(n2901[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_15 (.CI(n24255), .I0(n7348[12]), .I1(n1023), 
            .CO(n24256));
    SB_CARRY add_3444_8 (.CI(n24327), .I0(n7458[5]), .I1(n527_adj_4281), 
            .CO(n24328));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n19402), .I1(n7348[11]), .I2(n950), 
            .I3(n24254), .O(n2901[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_14 (.CI(n24254), .I0(n7348[11]), .I1(n950), 
            .CO(n24255));
    SB_LUT4 add_3444_7_lut (.I0(GND_net), .I1(n7458[4]), .I2(n454_adj_4280), 
            .I3(n24326), .O(n7438[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n19402), .I1(n7348[10]), .I2(n877), 
            .I3(n24253), .O(n2901[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_13 (.CI(n24253), .I0(n7348[10]), .I1(n877), 
            .CO(n24254));
    SB_CARRY add_3444_7 (.CI(n24326), .I0(n7458[4]), .I1(n454_adj_4280), 
            .CO(n24327));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n19402), .I1(n7348[9]), .I2(n804), 
            .I3(n24252), .O(n2901[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_12 (.CI(n24252), .I0(n7348[9]), .I1(n804), 
            .CO(n24253));
    SB_LUT4 add_3444_6_lut (.I0(GND_net), .I1(n7458[3]), .I2(n381_adj_4279), 
            .I3(n24325), .O(n7438[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n19402), .I1(n7348[8]), .I2(n731), 
            .I3(n24251), .O(n2901[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_11 (.CI(n24251), .I0(n7348[8]), .I1(n731), 
            .CO(n24252));
    SB_CARRY add_3444_6 (.CI(n24325), .I0(n7458[3]), .I1(n381_adj_4279), 
            .CO(n24326));
    SB_LUT4 add_3444_5_lut (.I0(GND_net), .I1(n7458[2]), .I2(n308_adj_4278), 
            .I3(n24324), .O(n7438[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3467_10_lut (.I0(GND_net), .I1(n7774[7]), .I2(n676), .I3(n24589), 
            .O(n7755[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_10 (.CI(n24589), .I0(n7774[7]), .I1(n676), .CO(n24590));
    SB_LUT4 add_3467_9_lut (.I0(GND_net), .I1(n7774[6]), .I2(n603), .I3(n24588), 
            .O(n7755[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_9 (.CI(n24588), .I0(n7774[6]), .I1(n603), .CO(n24589));
    SB_LUT4 add_3467_8_lut (.I0(GND_net), .I1(n7774[5]), .I2(n530), .I3(n24587), 
            .O(n7755[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_8 (.CI(n24587), .I0(n7774[5]), .I1(n530), .CO(n24588));
    SB_CARRY add_3444_5 (.CI(n24324), .I0(n7458[2]), .I1(n308_adj_4278), 
            .CO(n24325));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n19402), .I1(n7348[7]), .I2(n658), 
            .I3(n24250), .O(n2901[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_10 (.CI(n24250), .I0(n7348[7]), .I1(n658), 
            .CO(n24251));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n19402), .I1(n7348[6]), .I2(n585), 
            .I3(n24249), .O(n2901[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3467_7_lut (.I0(GND_net), .I1(n7774[4]), .I2(n457), .I3(n24586), 
            .O(n7755[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_7 (.CI(n24586), .I0(n7774[4]), .I1(n457), .CO(n24587));
    SB_LUT4 add_3467_6_lut (.I0(GND_net), .I1(n7774[3]), .I2(n384), .I3(n24585), 
            .O(n7755[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n24249), .I0(n7348[6]), .I1(n585), 
            .CO(n24250));
    SB_CARRY add_3467_6 (.CI(n24585), .I0(n7774[3]), .I1(n384), .CO(n24586));
    SB_LUT4 add_3467_5_lut (.I0(GND_net), .I1(n7774[2]), .I2(n311), .I3(n24584), 
            .O(n7755[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_5 (.CI(n24584), .I0(n7774[2]), .I1(n311), .CO(n24585));
    SB_LUT4 add_3467_4_lut (.I0(GND_net), .I1(n7774[1]), .I2(n238), .I3(n24583), 
            .O(n7755[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_4 (.CI(n24583), .I0(n7774[1]), .I1(n238), .CO(n24584));
    SB_LUT4 add_3467_3_lut (.I0(GND_net), .I1(n7774[0]), .I2(n165), .I3(n24582), 
            .O(n7755[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_3 (.CI(n24582), .I0(n7774[0]), .I1(n165), .CO(n24583));
    SB_LUT4 add_3467_2_lut (.I0(GND_net), .I1(n23_adj_4276), .I2(n92), 
            .I3(GND_net), .O(n7755[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3467_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3467_2 (.CI(GND_net), .I0(n23_adj_4276), .I1(n92), .CO(n24582));
    SB_LUT4 add_3466_19_lut (.I0(GND_net), .I1(n7755[16]), .I2(GND_net), 
            .I3(n24581), .O(n7735[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3466_18_lut (.I0(GND_net), .I1(n7755[15]), .I2(GND_net), 
            .I3(n24580), .O(n7735[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_18 (.CI(n24580), .I0(n7755[15]), .I1(GND_net), .CO(n24581));
    SB_LUT4 add_3466_17_lut (.I0(GND_net), .I1(n7755[14]), .I2(GND_net), 
            .I3(n24579), .O(n7735[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n19402), .I1(n7348[5]), .I2(n512), 
            .I3(n24248), .O(n2901[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3444_4_lut (.I0(GND_net), .I1(n7458[1]), .I2(n235_adj_4274), 
            .I3(n24323), .O(n7438[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3444_4 (.CI(n24323), .I0(n7458[1]), .I1(n235_adj_4274), 
            .CO(n24324));
    SB_CARRY add_3466_17 (.CI(n24579), .I0(n7755[14]), .I1(GND_net), .CO(n24580));
    SB_LUT4 add_3444_3_lut (.I0(GND_net), .I1(n7458[0]), .I2(n162_adj_4273), 
            .I3(n24322), .O(n7438[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_8 (.CI(n24248), .I0(n7348[5]), .I1(n512), 
            .CO(n24249));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n19402), .I1(n7348[4]), .I2(n439), 
            .I3(n24247), .O(n2901[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_7 (.CI(n24247), .I0(n7348[4]), .I1(n439), 
            .CO(n24248));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n19402), .I1(n7348[3]), .I2(n366), 
            .I3(n24246), .O(n2901[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3444_3 (.CI(n24322), .I0(n7458[0]), .I1(n162_adj_4273), 
            .CO(n24323));
    SB_CARRY mult_10_add_1225_6 (.CI(n24246), .I0(n7348[3]), .I1(n366), 
            .CO(n24247));
    SB_LUT4 add_3444_2_lut (.I0(GND_net), .I1(n20_adj_4263), .I2(n89_adj_4262), 
            .I3(GND_net), .O(n7438[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3444_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n19402), .I1(n7348[2]), .I2(n293), 
            .I3(n24245), .O(n2901[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3444_2 (.CI(GND_net), .I0(n20_adj_4263), .I1(n89_adj_4262), 
            .CO(n24322));
    SB_LUT4 add_3443_20_lut (.I0(GND_net), .I1(n7438[17]), .I2(GND_net), 
            .I3(n24321), .O(n7417[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3466_16_lut (.I0(GND_net), .I1(n7755[13]), .I2(n1111), 
            .I3(n24578), .O(n7735[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_16 (.CI(n24578), .I0(n7755[13]), .I1(n1111), .CO(n24579));
    SB_LUT4 add_3466_15_lut (.I0(GND_net), .I1(n7755[12]), .I2(n1038), 
            .I3(n24577), .O(n7735[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_19_lut (.I0(GND_net), .I1(n7438[16]), .I2(GND_net), 
            .I3(n24320), .O(n7417[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_15 (.CI(n24577), .I0(n7755[12]), .I1(n1038), .CO(n24578));
    SB_LUT4 add_3466_14_lut (.I0(GND_net), .I1(n7755[11]), .I2(n965), 
            .I3(n24576), .O(n7735[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_14 (.CI(n24576), .I0(n7755[11]), .I1(n965), .CO(n24577));
    SB_LUT4 add_3466_13_lut (.I0(GND_net), .I1(n7755[10]), .I2(n892), 
            .I3(n24575), .O(n7735[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_13 (.CI(n24575), .I0(n7755[10]), .I1(n892), .CO(n24576));
    SB_LUT4 add_3466_12_lut (.I0(GND_net), .I1(n7755[9]), .I2(n819), .I3(n24574), 
            .O(n7735[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_19 (.CI(n24320), .I0(n7438[16]), .I1(GND_net), .CO(n24321));
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3528[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_3443_18_lut (.I0(GND_net), .I1(n7438[15]), .I2(GND_net), 
            .I3(n24319), .O(n7417[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_12 (.CI(n24574), .I0(n7755[9]), .I1(n819), .CO(n24575));
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4511));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3466_11_lut (.I0(GND_net), .I1(n7755[8]), .I2(n746), .I3(n24573), 
            .O(n7735[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_18 (.CI(n24319), .I0(n7438[15]), .I1(GND_net), .CO(n24320));
    SB_CARRY mult_10_add_1225_5 (.CI(n24245), .I0(n7348[2]), .I1(n293), 
            .CO(n24246));
    SB_LUT4 add_3443_17_lut (.I0(GND_net), .I1(n7438[14]), .I2(GND_net), 
            .I3(n24318), .O(n7417[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_17 (.CI(n24318), .I0(n7438[14]), .I1(GND_net), .CO(n24319));
    SB_LUT4 add_3443_16_lut (.I0(GND_net), .I1(n7438[13]), .I2(n1108_adj_4246), 
            .I3(n24317), .O(n7417[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_16 (.CI(n24317), .I0(n7438[13]), .I1(n1108_adj_4246), 
            .CO(n24318));
    SB_CARRY add_3466_11 (.CI(n24573), .I0(n7755[8]), .I1(n746), .CO(n24574));
    SB_LUT4 add_3466_10_lut (.I0(GND_net), .I1(n7755[7]), .I2(n673_adj_4242), 
            .I3(n24572), .O(n7735[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_10 (.CI(n24572), .I0(n7755[7]), .I1(n673_adj_4242), 
            .CO(n24573));
    SB_LUT4 add_3466_9_lut (.I0(GND_net), .I1(n7755[6]), .I2(n600_adj_4241), 
            .I3(n24571), .O(n7735[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_9 (.CI(n24571), .I0(n7755[6]), .I1(n600_adj_4241), 
            .CO(n24572));
    SB_LUT4 add_3466_8_lut (.I0(GND_net), .I1(n7755[5]), .I2(n527), .I3(n24570), 
            .O(n7735[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_8 (.CI(n24570), .I0(n7755[5]), .I1(n527), .CO(n24571));
    SB_LUT4 add_3466_7_lut (.I0(GND_net), .I1(n7755[4]), .I2(n454), .I3(n24569), 
            .O(n7735[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_7 (.CI(n24569), .I0(n7755[4]), .I1(n454), .CO(n24570));
    SB_LUT4 add_3466_6_lut (.I0(GND_net), .I1(n7755[3]), .I2(n381), .I3(n24568), 
            .O(n7735[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_6 (.CI(n24568), .I0(n7755[3]), .I1(n381), .CO(n24569));
    SB_LUT4 add_3466_5_lut (.I0(GND_net), .I1(n7755[2]), .I2(n308), .I3(n24567), 
            .O(n7735[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_5 (.CI(n24567), .I0(n7755[2]), .I1(n308), .CO(n24568));
    SB_LUT4 add_3466_4_lut (.I0(GND_net), .I1(n7755[1]), .I2(n235), .I3(n24566), 
            .O(n7735[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_4 (.CI(n24566), .I0(n7755[1]), .I1(n235), .CO(n24567));
    SB_LUT4 add_3466_3_lut (.I0(GND_net), .I1(n7755[0]), .I2(n162), .I3(n24565), 
            .O(n7735[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_3 (.CI(n24565), .I0(n7755[0]), .I1(n162), .CO(n24566));
    SB_LUT4 add_3466_2_lut (.I0(GND_net), .I1(n20_adj_4232), .I2(n89), 
            .I3(GND_net), .O(n7735[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3466_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3466_2 (.CI(GND_net), .I0(n20_adj_4232), .I1(n89), .CO(n24565));
    SB_LUT4 add_3443_15_lut (.I0(GND_net), .I1(n7438[12]), .I2(n1035_adj_4223), 
            .I3(n24316), .O(n7417[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3465_20_lut (.I0(GND_net), .I1(n7735[17]), .I2(GND_net), 
            .I3(n24564), .O(n7714[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3465_19_lut (.I0(GND_net), .I1(n7735[16]), .I2(GND_net), 
            .I3(n24563), .O(n7714[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_19 (.CI(n24563), .I0(n7735[16]), .I1(GND_net), .CO(n24564));
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4512));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3465_18_lut (.I0(GND_net), .I1(n7735[15]), .I2(GND_net), 
            .I3(n24562), .O(n7714[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_15 (.CI(n24316), .I0(n7438[12]), .I1(n1035_adj_4223), 
            .CO(n24317));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n19402), .I1(n7348[1]), .I2(n220), 
            .I3(n24244), .O(n2901[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3465_18 (.CI(n24562), .I0(n7735[15]), .I1(GND_net), .CO(n24563));
    SB_LUT4 add_3465_17_lut (.I0(GND_net), .I1(n7735[14]), .I2(GND_net), 
            .I3(n24561), .O(n7714[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_14_lut (.I0(GND_net), .I1(n7438[11]), .I2(n962_adj_4218), 
            .I3(n24315), .O(n7417[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_14 (.CI(n24315), .I0(n7438[11]), .I1(n962_adj_4218), 
            .CO(n24316));
    SB_LUT4 add_3443_13_lut (.I0(GND_net), .I1(n7438[10]), .I2(n889_adj_4215), 
            .I3(n24314), .O(n7417[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_13 (.CI(n24314), .I0(n7438[10]), .I1(n889_adj_4215), 
            .CO(n24315));
    SB_CARRY add_3465_17 (.CI(n24561), .I0(n7735[14]), .I1(GND_net), .CO(n24562));
    SB_LUT4 add_3443_12_lut (.I0(GND_net), .I1(n7438[9]), .I2(n816_adj_4212), 
            .I3(n24313), .O(n7417[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_12 (.CI(n24313), .I0(n7438[9]), .I1(n816_adj_4212), 
            .CO(n24314));
    SB_CARRY mult_10_add_1225_4 (.CI(n24244), .I0(n7348[1]), .I1(n220), 
            .CO(n24245));
    SB_LUT4 add_3443_11_lut (.I0(GND_net), .I1(n7438[8]), .I2(n743_adj_4208), 
            .I3(n24312), .O(n7417[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_11 (.CI(n24312), .I0(n7438[8]), .I1(n743_adj_4208), 
            .CO(n24313));
    SB_LUT4 add_3465_16_lut (.I0(GND_net), .I1(n7735[13]), .I2(n1108), 
            .I3(n24560), .O(n7714[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n19402), .I1(n7348[0]), .I2(n147), 
            .I3(n24243), .O(n2901[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i18812_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral [19]), .O(n7924[0]));   // verilog/motorControl.v(34[26:37])
    defparam i18812_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY mult_10_add_1225_3 (.CI(n24243), .I0(n7348[0]), .I1(n147), 
            .CO(n24244));
    SB_LUT4 add_3443_10_lut (.I0(GND_net), .I1(n7438[7]), .I2(n670_adj_4205), 
            .I3(n24311), .O(n7417[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_16 (.CI(n24560), .I0(n7735[13]), .I1(n1108), .CO(n24561));
    SB_CARRY add_3443_10 (.CI(n24311), .I0(n7438[7]), .I1(n670_adj_4205), 
            .CO(n24312));
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3528[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3528[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3528[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3528[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3528[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3528[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3528[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3528[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3528[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3528[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3528[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3528[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3528[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3528[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3528[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3528[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3528[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3528[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3528[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3528[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3528[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3552 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_3465_15_lut (.I0(GND_net), .I1(n7735[12]), .I2(n1035), 
            .I3(n24559), .O(n7714[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n19402), .I1(n5_adj_4204), .I2(n74), 
            .I3(GND_net), .O(n2901[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3465_15 (.CI(n24559), .I0(n7735[12]), .I1(n1035), .CO(n24560));
    SB_LUT4 add_3465_14_lut (.I0(GND_net), .I1(n7735[11]), .I2(n962), 
            .I3(n24558), .O(n7714[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_9_lut (.I0(GND_net), .I1(n7438[6]), .I2(n597_adj_4203), 
            .I3(n24310), .O(n7417[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4204), .I1(n74), 
            .CO(n24243));
    SB_CARRY add_3465_14 (.CI(n24558), .I0(n7735[11]), .I1(n962), .CO(n24559));
    SB_LUT4 add_3465_13_lut (.I0(GND_net), .I1(n7735[10]), .I2(n889), 
            .I3(n24557), .O(n7714[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4513));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3465_13 (.CI(n24557), .I0(n7735[10]), .I1(n889), .CO(n24558));
    SB_LUT4 add_3465_12_lut (.I0(GND_net), .I1(n7735[9]), .I2(n816), .I3(n24556), 
            .O(n7714[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_9 (.CI(n24310), .I0(n7438[6]), .I1(n597_adj_4203), 
            .CO(n24311));
    SB_CARRY add_3465_12 (.CI(n24556), .I0(n7735[9]), .I1(n816), .CO(n24557));
    SB_LUT4 add_3465_11_lut (.I0(GND_net), .I1(n7735[8]), .I2(n743), .I3(n24555), 
            .O(n7714[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_11 (.CI(n24555), .I0(n7735[8]), .I1(n743), .CO(n24556));
    SB_LUT4 add_3465_10_lut (.I0(GND_net), .I1(n7735[7]), .I2(n670), .I3(n24554), 
            .O(n7714[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_10 (.CI(n24554), .I0(n7735[7]), .I1(n670), .CO(n24555));
    SB_LUT4 add_3465_9_lut (.I0(GND_net), .I1(n7735[6]), .I2(n597), .I3(n24553), 
            .O(n7714[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_9 (.CI(n24553), .I0(n7735[6]), .I1(n597), .CO(n24554));
    SB_LUT4 add_3465_8_lut (.I0(GND_net), .I1(n7735[5]), .I2(n524_adj_4201), 
            .I3(n24552), .O(n7714[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_8 (.CI(n24552), .I0(n7735[5]), .I1(n524_adj_4201), 
            .CO(n24553));
    SB_LUT4 add_3465_7_lut (.I0(GND_net), .I1(n7735[4]), .I2(n451_adj_4200), 
            .I3(n24551), .O(n7714[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_7 (.CI(n24551), .I0(n7735[4]), .I1(n451_adj_4200), 
            .CO(n24552));
    SB_LUT4 add_3440_23_lut (.I0(GND_net), .I1(n7372[20]), .I2(GND_net), 
            .I3(n24242), .O(n7348[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3465_6_lut (.I0(GND_net), .I1(n7735[3]), .I2(n378_adj_4199), 
            .I3(n24550), .O(n7714[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_6 (.CI(n24550), .I0(n7735[3]), .I1(n378_adj_4199), 
            .CO(n24551));
    SB_LUT4 add_3443_8_lut (.I0(GND_net), .I1(n7438[5]), .I2(n524), .I3(n24309), 
            .O(n7417[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3465_5_lut (.I0(GND_net), .I1(n7735[2]), .I2(n305_adj_4198), 
            .I3(n24549), .O(n7714[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_5 (.CI(n24549), .I0(n7735[2]), .I1(n305_adj_4198), 
            .CO(n24550));
    SB_LUT4 add_3465_4_lut (.I0(GND_net), .I1(n7735[1]), .I2(n232_adj_4197), 
            .I3(n24548), .O(n7714[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_8 (.CI(n24309), .I0(n7438[5]), .I1(n524), .CO(n24310));
    SB_LUT4 add_3443_7_lut (.I0(GND_net), .I1(n7438[4]), .I2(n451), .I3(n24308), 
            .O(n7417[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_4 (.CI(n24548), .I0(n7735[1]), .I1(n232_adj_4197), 
            .CO(n24549));
    SB_LUT4 add_3465_3_lut (.I0(GND_net), .I1(n7735[0]), .I2(n159_adj_4191), 
            .I3(n24547), .O(n7714[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_3 (.CI(n24547), .I0(n7735[0]), .I1(n159_adj_4191), 
            .CO(n24548));
    SB_LUT4 add_3465_2_lut (.I0(GND_net), .I1(n17_adj_4189), .I2(n86), 
            .I3(GND_net), .O(n7714[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3465_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3465_2 (.CI(GND_net), .I0(n17_adj_4189), .I1(n86), .CO(n24547));
    SB_LUT4 add_3464_21_lut (.I0(GND_net), .I1(n7714[18]), .I2(GND_net), 
            .I3(n24546), .O(n7692[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_20_lut (.I0(GND_net), .I1(n7714[17]), .I2(GND_net), 
            .I3(n24545), .O(n7692[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_20 (.CI(n24545), .I0(n7714[17]), .I1(GND_net), .CO(n24546));
    SB_LUT4 add_3464_19_lut (.I0(GND_net), .I1(n7714[16]), .I2(GND_net), 
            .I3(n24544), .O(n7692[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_19 (.CI(n24544), .I0(n7714[16]), .I1(GND_net), .CO(n24545));
    SB_LUT4 add_3440_22_lut (.I0(GND_net), .I1(n7372[19]), .I2(GND_net), 
            .I3(n24241), .O(n7348[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_18_lut (.I0(GND_net), .I1(n7714[15]), .I2(GND_net), 
            .I3(n24543), .O(n7692[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_18 (.CI(n24543), .I0(n7714[15]), .I1(GND_net), .CO(n24544));
    SB_LUT4 add_3464_17_lut (.I0(GND_net), .I1(n7714[14]), .I2(GND_net), 
            .I3(n24542), .O(n7692[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4514));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3464_17 (.CI(n24542), .I0(n7714[14]), .I1(GND_net), .CO(n24543));
    SB_CARRY add_3440_22 (.CI(n24241), .I0(n7372[19]), .I1(GND_net), .CO(n24242));
    SB_LUT4 add_3440_21_lut (.I0(GND_net), .I1(n7372[18]), .I2(GND_net), 
            .I3(n24240), .O(n7348[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_16_lut (.I0(GND_net), .I1(n7714[13]), .I2(n1105), 
            .I3(n24541), .O(n7692[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_16 (.CI(n24541), .I0(n7714[13]), .I1(n1105), .CO(n24542));
    SB_LUT4 add_3464_15_lut (.I0(GND_net), .I1(n7714[12]), .I2(n1032), 
            .I3(n24540), .O(n7692[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_15 (.CI(n24540), .I0(n7714[12]), .I1(n1032), .CO(n24541));
    SB_CARRY add_3440_21 (.CI(n24240), .I0(n7372[18]), .I1(GND_net), .CO(n24241));
    SB_CARRY add_3443_7 (.CI(n24308), .I0(n7438[4]), .I1(n451), .CO(n24309));
    SB_LUT4 add_3464_14_lut (.I0(GND_net), .I1(n7714[11]), .I2(n959), 
            .I3(n24539), .O(n7692[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_6_lut (.I0(GND_net), .I1(n7438[3]), .I2(n378), .I3(n24307), 
            .O(n7417[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_14 (.CI(n24539), .I0(n7714[11]), .I1(n959), .CO(n24540));
    SB_LUT4 add_3440_20_lut (.I0(GND_net), .I1(n7372[17]), .I2(GND_net), 
            .I3(n24239), .O(n7348[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_13_lut (.I0(GND_net), .I1(n7714[10]), .I2(n886), 
            .I3(n24538), .O(n7692[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_20 (.CI(n24239), .I0(n7372[17]), .I1(GND_net), .CO(n24240));
    SB_CARRY add_3464_13 (.CI(n24538), .I0(n7714[10]), .I1(n886), .CO(n24539));
    SB_LUT4 add_3464_12_lut (.I0(GND_net), .I1(n7714[9]), .I2(n813), .I3(n24537), 
            .O(n7692[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_12 (.CI(n24537), .I0(n7714[9]), .I1(n813), .CO(n24538));
    SB_CARRY add_3443_6 (.CI(n24307), .I0(n7438[3]), .I1(n378), .CO(n24308));
    SB_LUT4 add_3443_5_lut (.I0(GND_net), .I1(n7438[2]), .I2(n305), .I3(n24306), 
            .O(n7417[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_5 (.CI(n24306), .I0(n7438[2]), .I1(n305), .CO(n24307));
    SB_LUT4 add_3443_4_lut (.I0(GND_net), .I1(n7438[1]), .I2(n232), .I3(n24305), 
            .O(n7417[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_11_lut (.I0(GND_net), .I1(n7714[8]), .I2(n740), .I3(n24536), 
            .O(n7692[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_11 (.CI(n24536), .I0(n7714[8]), .I1(n740), .CO(n24537));
    SB_LUT4 add_3464_10_lut (.I0(GND_net), .I1(n7714[7]), .I2(n667), .I3(n24535), 
            .O(n7692[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_10 (.CI(n24535), .I0(n7714[7]), .I1(n667), .CO(n24536));
    SB_LUT4 add_3464_9_lut (.I0(GND_net), .I1(n7714[6]), .I2(n594), .I3(n24534), 
            .O(n7692[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_9 (.CI(n24534), .I0(n7714[6]), .I1(n594), .CO(n24535));
    SB_LUT4 add_3464_8_lut (.I0(GND_net), .I1(n7714[5]), .I2(n521), .I3(n24533), 
            .O(n7692[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_4 (.CI(n24305), .I0(n7438[1]), .I1(n232), .CO(n24306));
    SB_CARRY add_3464_8 (.CI(n24533), .I0(n7714[5]), .I1(n521), .CO(n24534));
    SB_LUT4 add_3464_7_lut (.I0(GND_net), .I1(n7714[4]), .I2(n448), .I3(n24532), 
            .O(n7692[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_7 (.CI(n24532), .I0(n7714[4]), .I1(n448), .CO(n24533));
    SB_LUT4 add_3464_6_lut (.I0(GND_net), .I1(n7714[3]), .I2(n375), .I3(n24531), 
            .O(n7692[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_6 (.CI(n24531), .I0(n7714[3]), .I1(n375), .CO(n24532));
    SB_LUT4 add_3464_5_lut (.I0(GND_net), .I1(n7714[2]), .I2(n302), .I3(n24530), 
            .O(n7692[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_5 (.CI(n24530), .I0(n7714[2]), .I1(n302), .CO(n24531));
    SB_LUT4 add_3464_4_lut (.I0(GND_net), .I1(n7714[1]), .I2(n229), .I3(n24529), 
            .O(n7692[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_4 (.CI(n24529), .I0(n7714[1]), .I1(n229), .CO(n24530));
    SB_LUT4 add_3464_3_lut (.I0(GND_net), .I1(n7714[0]), .I2(n156_adj_4181), 
            .I3(n24528), .O(n7692[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_3 (.CI(n24528), .I0(n7714[0]), .I1(n156_adj_4181), 
            .CO(n24529));
    SB_LUT4 add_3464_2_lut (.I0(GND_net), .I1(n14_adj_4180), .I2(n83_adj_4179), 
            .I3(GND_net), .O(n7692[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_2 (.CI(GND_net), .I0(n14_adj_4180), .I1(n83_adj_4179), 
            .CO(n24528));
    SB_LUT4 add_3463_22_lut (.I0(GND_net), .I1(n7692[19]), .I2(GND_net), 
            .I3(n24527), .O(n7669[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3463_21_lut (.I0(GND_net), .I1(n7692[18]), .I2(GND_net), 
            .I3(n24526), .O(n7669[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_21 (.CI(n24526), .I0(n7692[18]), .I1(GND_net), .CO(n24527));
    SB_LUT4 add_3463_20_lut (.I0(GND_net), .I1(n7692[17]), .I2(GND_net), 
            .I3(n24525), .O(n7669[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25347_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n31178));
    defparam i25347_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_3463_20 (.CI(n24525), .I0(n7692[17]), .I1(GND_net), .CO(n24526));
    SB_LUT4 i25357_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n31188));
    defparam i25357_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4515));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4516));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4517));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4518));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4328));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4519));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3463_19_lut (.I0(GND_net), .I1(n7692[16]), .I2(GND_net), 
            .I3(n24524), .O(n7669[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_19 (.CI(n24524), .I0(n7692[16]), .I1(GND_net), .CO(n24525));
    SB_LUT4 add_3463_18_lut (.I0(GND_net), .I1(n7692[15]), .I2(GND_net), 
            .I3(n24523), .O(n7669[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3440_19_lut (.I0(GND_net), .I1(n7372[16]), .I2(GND_net), 
            .I3(n24238), .O(n7348[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_3_lut (.I0(GND_net), .I1(n7438[0]), .I2(n159), .I3(n24304), 
            .O(n7417[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_18 (.CI(n24523), .I0(n7692[15]), .I1(GND_net), .CO(n24524));
    SB_CARRY add_3440_19 (.CI(n24238), .I0(n7372[16]), .I1(GND_net), .CO(n24239));
    SB_LUT4 add_3463_17_lut (.I0(GND_net), .I1(n7692[14]), .I2(GND_net), 
            .I3(n24522), .O(n7669[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_17 (.CI(n24522), .I0(n7692[14]), .I1(GND_net), .CO(n24523));
    SB_LUT4 add_3463_16_lut (.I0(GND_net), .I1(n7692[13]), .I2(n1102), 
            .I3(n24521), .O(n7669[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_16 (.CI(n24521), .I0(n7692[13]), .I1(n1102), .CO(n24522));
    SB_LUT4 add_3463_15_lut (.I0(GND_net), .I1(n7692[12]), .I2(n1029), 
            .I3(n24520), .O(n7669[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_15 (.CI(n24520), .I0(n7692[12]), .I1(n1029), .CO(n24521));
    SB_LUT4 add_3463_14_lut (.I0(GND_net), .I1(n7692[11]), .I2(n956), 
            .I3(n24519), .O(n7669[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_14 (.CI(n24519), .I0(n7692[11]), .I1(n956), .CO(n24520));
    SB_LUT4 add_3463_13_lut (.I0(GND_net), .I1(n7692[10]), .I2(n883_adj_4520), 
            .I3(n24518), .O(n7669[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_13 (.CI(n24518), .I0(n7692[10]), .I1(n883_adj_4520), 
            .CO(n24519));
    SB_LUT4 add_3463_12_lut (.I0(GND_net), .I1(n7692[9]), .I2(n810_adj_4521), 
            .I3(n24517), .O(n7669[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_12 (.CI(n24517), .I0(n7692[9]), .I1(n810_adj_4521), 
            .CO(n24518));
    SB_LUT4 add_3463_11_lut (.I0(GND_net), .I1(n7692[8]), .I2(n737_adj_4522), 
            .I3(n24516), .O(n7669[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_11 (.CI(n24516), .I0(n7692[8]), .I1(n737_adj_4522), 
            .CO(n24517));
    SB_LUT4 add_3463_10_lut (.I0(GND_net), .I1(n7692[7]), .I2(n664_adj_4523), 
            .I3(n24515), .O(n7669[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_10 (.CI(n24515), .I0(n7692[7]), .I1(n664_adj_4523), 
            .CO(n24516));
    SB_LUT4 add_3463_9_lut (.I0(GND_net), .I1(n7692[6]), .I2(n591_adj_4524), 
            .I3(n24514), .O(n7669[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_9 (.CI(n24514), .I0(n7692[6]), .I1(n591_adj_4524), 
            .CO(n24515));
    SB_LUT4 add_3463_8_lut (.I0(GND_net), .I1(n7692[5]), .I2(n518_adj_4525), 
            .I3(n24513), .O(n7669[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_8 (.CI(n24513), .I0(n7692[5]), .I1(n518_adj_4525), 
            .CO(n24514));
    SB_LUT4 add_3463_7_lut (.I0(GND_net), .I1(n7692[4]), .I2(n445_adj_4526), 
            .I3(n24512), .O(n7669[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3440_18_lut (.I0(GND_net), .I1(n7372[15]), .I2(GND_net), 
            .I3(n24237), .O(n7348[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_7 (.CI(n24512), .I0(n7692[4]), .I1(n445_adj_4526), 
            .CO(n24513));
    SB_LUT4 add_3463_6_lut (.I0(GND_net), .I1(n7692[3]), .I2(n372_adj_4527), 
            .I3(n24511), .O(n7669[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_6 (.CI(n24511), .I0(n7692[3]), .I1(n372_adj_4527), 
            .CO(n24512));
    SB_LUT4 add_3463_5_lut (.I0(GND_net), .I1(n7692[2]), .I2(n299_adj_4528), 
            .I3(n24510), .O(n7669[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_5 (.CI(n24510), .I0(n7692[2]), .I1(n299_adj_4528), 
            .CO(n24511));
    SB_CARRY add_3440_18 (.CI(n24237), .I0(n7372[15]), .I1(GND_net), .CO(n24238));
    SB_LUT4 add_3463_4_lut (.I0(GND_net), .I1(n7692[1]), .I2(n226_adj_4529), 
            .I3(n24509), .O(n7669[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_4 (.CI(n24509), .I0(n7692[1]), .I1(n226_adj_4529), 
            .CO(n24510));
    SB_LUT4 add_3463_3_lut (.I0(GND_net), .I1(n7692[0]), .I2(n153_adj_4530), 
            .I3(n24508), .O(n7669[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_3 (.CI(n24508), .I0(n7692[0]), .I1(n153_adj_4530), 
            .CO(n24509));
    SB_LUT4 add_3463_2_lut (.I0(GND_net), .I1(n11_adj_4531), .I2(n80_adj_4532), 
            .I3(GND_net), .O(n7669[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3463_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3440_17_lut (.I0(GND_net), .I1(n7372[14]), .I2(GND_net), 
            .I3(n24236), .O(n7348[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_17 (.CI(n24236), .I0(n7372[14]), .I1(GND_net), .CO(n24237));
    SB_LUT4 add_3440_16_lut (.I0(GND_net), .I1(n7372[13]), .I2(n1099), 
            .I3(n24235), .O(n7348[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_3 (.CI(n24304), .I0(n7438[0]), .I1(n159), .CO(n24305));
    SB_LUT4 add_3443_2_lut (.I0(GND_net), .I1(n17_adj_4533), .I2(n86_adj_4534), 
            .I3(GND_net), .O(n7417[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_16 (.CI(n24235), .I0(n7372[13]), .I1(n1099), .CO(n24236));
    SB_LUT4 add_3440_15_lut (.I0(GND_net), .I1(n7372[12]), .I2(n1026), 
            .I3(n24234), .O(n7348[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3463_2 (.CI(GND_net), .I0(n11_adj_4531), .I1(n80_adj_4532), 
            .CO(n24508));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n7645[21]), 
            .I2(GND_net), .I3(n24507), .O(n31114)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n7645[20]), .I2(GND_net), 
            .I3(n24506), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n24506), .I0(n7645[20]), .I1(GND_net), 
            .CO(n24507));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n7645[19]), .I2(GND_net), 
            .I3(n24505), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n24505), .I0(n7645[19]), .I1(GND_net), 
            .CO(n24506));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n7645[18]), .I2(GND_net), 
            .I3(n24504), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n24504), .I0(n7645[18]), .I1(GND_net), 
            .CO(n24505));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n7645[17]), .I2(GND_net), 
            .I3(n24503), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n24503), .I0(n7645[17]), .I1(GND_net), 
            .CO(n24504));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n7645[16]), .I2(GND_net), 
            .I3(n24502), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n24502), .I0(n7645[16]), .I1(GND_net), 
            .CO(n24503));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n7645[15]), .I2(GND_net), 
            .I3(n24501), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n24501), .I0(n7645[15]), .I1(GND_net), 
            .CO(n24502));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n7645[14]), .I2(GND_net), 
            .I3(n24500), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n24500), .I0(n7645[14]), .I1(GND_net), 
            .CO(n24501));
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4535));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4383));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n7645[13]), .I2(n1096_adj_4536), 
            .I3(n24499), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n24499), .I0(n7645[13]), .I1(n1096_adj_4536), 
            .CO(n24500));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n7645[12]), .I2(n1023_adj_4537), 
            .I3(n24498), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n24498), .I0(n7645[12]), .I1(n1023_adj_4537), 
            .CO(n24499));
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4377));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4387));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n7645[11]), .I2(n950_adj_4538), 
            .I3(n24497), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n24497), .I0(n7645[11]), .I1(n950_adj_4538), 
            .CO(n24498));
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4539));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n7645[10]), .I2(n877_adj_4540), 
            .I3(n24496), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n24496), .I0(n7645[10]), .I1(n877_adj_4540), 
            .CO(n24497));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n7645[9]), .I2(n804_adj_4541), 
            .I3(n24495), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n24495), .I0(n7645[9]), .I1(n804_adj_4541), 
            .CO(n24496));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n7645[8]), .I2(n731_adj_4542), 
            .I3(n24494), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n24494), .I0(n7645[8]), .I1(n731_adj_4542), 
            .CO(n24495));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n7645[7]), .I2(n658_adj_4543), 
            .I3(n24493), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n24493), .I0(n7645[7]), .I1(n658_adj_4543), 
            .CO(n24494));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n7645[6]), .I2(n585_adj_4544), 
            .I3(n24492), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n24492), .I0(n7645[6]), .I1(n585_adj_4544), 
            .CO(n24493));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n7645[5]), .I2(n512_adj_4545), 
            .I3(n24491), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n24491), .I0(n7645[5]), .I1(n512_adj_4545), 
            .CO(n24492));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n7645[4]), .I2(n439_adj_4546), 
            .I3(n24490), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n24490), .I0(n7645[4]), .I1(n439_adj_4546), 
            .CO(n24491));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n7645[3]), .I2(n366_adj_4547), 
            .I3(n24489), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n24489), .I0(n7645[3]), .I1(n366_adj_4547), 
            .CO(n24490));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n7645[2]), .I2(n293_adj_4548), 
            .I3(n24488), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4399));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_11_add_1225_5 (.CI(n24488), .I0(n7645[2]), .I1(n293_adj_4548), 
            .CO(n24489));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n7645[1]), .I2(n220_adj_4549), 
            .I3(n24487), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n24487), .I0(n7645[1]), .I1(n220_adj_4549), 
            .CO(n24488));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n7645[0]), .I2(n147_adj_4550), 
            .I3(n24486), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n24486), .I0(n7645[0]), .I1(n147_adj_4550), 
            .CO(n24487));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4551), .I2(n74_adj_4552), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4551), .I1(n74_adj_4552), 
            .CO(n24486));
    SB_LUT4 add_3462_23_lut (.I0(GND_net), .I1(n7669[20]), .I2(GND_net), 
            .I3(n24485), .O(n7645[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3462_22_lut (.I0(GND_net), .I1(n7669[19]), .I2(GND_net), 
            .I3(n24484), .O(n7645[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_22 (.CI(n24484), .I0(n7669[19]), .I1(GND_net), .CO(n24485));
    SB_LUT4 add_3462_21_lut (.I0(GND_net), .I1(n7669[18]), .I2(GND_net), 
            .I3(n24483), .O(n7645[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_21 (.CI(n24483), .I0(n7669[18]), .I1(GND_net), .CO(n24484));
    SB_LUT4 add_3462_20_lut (.I0(GND_net), .I1(n7669[17]), .I2(GND_net), 
            .I3(n24482), .O(n7645[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_20 (.CI(n24482), .I0(n7669[17]), .I1(GND_net), .CO(n24483));
    SB_LUT4 add_3462_19_lut (.I0(GND_net), .I1(n7669[16]), .I2(GND_net), 
            .I3(n24481), .O(n7645[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_19 (.CI(n24481), .I0(n7669[16]), .I1(GND_net), .CO(n24482));
    SB_LUT4 add_3462_18_lut (.I0(GND_net), .I1(n7669[15]), .I2(GND_net), 
            .I3(n24480), .O(n7645[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_18 (.CI(n24480), .I0(n7669[15]), .I1(GND_net), .CO(n24481));
    SB_LUT4 add_3462_17_lut (.I0(GND_net), .I1(n7669[14]), .I2(GND_net), 
            .I3(n24479), .O(n7645[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_17 (.CI(n24479), .I0(n7669[14]), .I1(GND_net), .CO(n24480));
    SB_LUT4 add_3462_16_lut (.I0(GND_net), .I1(n7669[13]), .I2(n1099_adj_4553), 
            .I3(n24478), .O(n7645[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_16 (.CI(n24478), .I0(n7669[13]), .I1(n1099_adj_4553), 
            .CO(n24479));
    SB_LUT4 add_3462_15_lut (.I0(GND_net), .I1(n7669[12]), .I2(n1026_adj_4554), 
            .I3(n24477), .O(n7645[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_15 (.CI(n24477), .I0(n7669[12]), .I1(n1026_adj_4554), 
            .CO(n24478));
    SB_LUT4 add_3462_14_lut (.I0(GND_net), .I1(n7669[11]), .I2(n953_adj_4555), 
            .I3(n24476), .O(n7645[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_14 (.CI(n24476), .I0(n7669[11]), .I1(n953_adj_4555), 
            .CO(n24477));
    SB_LUT4 add_3462_13_lut (.I0(GND_net), .I1(n7669[10]), .I2(n880_adj_4556), 
            .I3(n24475), .O(n7645[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_13 (.CI(n24475), .I0(n7669[10]), .I1(n880_adj_4556), 
            .CO(n24476));
    SB_LUT4 add_3462_12_lut (.I0(GND_net), .I1(n7669[9]), .I2(n807_adj_4557), 
            .I3(n24474), .O(n7645[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_12 (.CI(n24474), .I0(n7669[9]), .I1(n807_adj_4557), 
            .CO(n24475));
    SB_LUT4 add_3462_11_lut (.I0(GND_net), .I1(n7669[8]), .I2(n734_adj_4558), 
            .I3(n24473), .O(n7645[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_11 (.CI(n24473), .I0(n7669[8]), .I1(n734_adj_4558), 
            .CO(n24474));
    SB_LUT4 add_3462_10_lut (.I0(GND_net), .I1(n7669[7]), .I2(n661_adj_4559), 
            .I3(n24472), .O(n7645[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_10 (.CI(n24472), .I0(n7669[7]), .I1(n661_adj_4559), 
            .CO(n24473));
    SB_LUT4 add_3462_9_lut (.I0(GND_net), .I1(n7669[6]), .I2(n588_adj_4560), 
            .I3(n24471), .O(n7645[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_9 (.CI(n24471), .I0(n7669[6]), .I1(n588_adj_4560), 
            .CO(n24472));
    SB_LUT4 add_3462_8_lut (.I0(GND_net), .I1(n7669[5]), .I2(n515_adj_4561), 
            .I3(n24470), .O(n7645[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_8 (.CI(n24470), .I0(n7669[5]), .I1(n515_adj_4561), 
            .CO(n24471));
    SB_LUT4 add_3462_7_lut (.I0(GND_net), .I1(n7669[4]), .I2(n442_adj_4562), 
            .I3(n24469), .O(n7645[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_7 (.CI(n24469), .I0(n7669[4]), .I1(n442_adj_4562), 
            .CO(n24470));
    SB_LUT4 add_3462_6_lut (.I0(GND_net), .I1(n7669[3]), .I2(n369_adj_4563), 
            .I3(n24468), .O(n7645[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_6 (.CI(n24468), .I0(n7669[3]), .I1(n369_adj_4563), 
            .CO(n24469));
    SB_LUT4 add_3462_5_lut (.I0(GND_net), .I1(n7669[2]), .I2(n296_adj_4564), 
            .I3(n24467), .O(n7645[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_5 (.CI(n24467), .I0(n7669[2]), .I1(n296_adj_4564), 
            .CO(n24468));
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4384));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3462_4_lut (.I0(GND_net), .I1(n7669[1]), .I2(n223_adj_4565), 
            .I3(n24466), .O(n7645[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_4 (.CI(n24466), .I0(n7669[1]), .I1(n223_adj_4565), 
            .CO(n24467));
    SB_LUT4 add_3462_3_lut (.I0(GND_net), .I1(n7669[0]), .I2(n150_adj_4566), 
            .I3(n24465), .O(n7645[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_3 (.CI(n24465), .I0(n7669[0]), .I1(n150_adj_4566), 
            .CO(n24466));
    SB_LUT4 add_3462_2_lut (.I0(GND_net), .I1(n8_adj_4567), .I2(n77_adj_4568), 
            .I3(GND_net), .O(n7645[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_2 (.CI(GND_net), .I0(n8_adj_4567), .I1(n77_adj_4568), 
            .CO(n24465));
    SB_LUT4 add_3456_7_lut (.I0(GND_net), .I1(n29930), .I2(n490_adj_4569), 
            .I3(n24464), .O(n7612[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3456_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3456_6_lut (.I0(GND_net), .I1(n7620[3]), .I2(n417_adj_4570), 
            .I3(n24463), .O(n7612[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3456_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3456_6 (.CI(n24463), .I0(n7620[3]), .I1(n417_adj_4570), 
            .CO(n24464));
    SB_LUT4 add_3456_5_lut (.I0(GND_net), .I1(n7620[2]), .I2(n344_adj_4571), 
            .I3(n24462), .O(n7612[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3456_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3456_5 (.CI(n24462), .I0(n7620[2]), .I1(n344_adj_4571), 
            .CO(n24463));
    SB_LUT4 add_3456_4_lut (.I0(GND_net), .I1(n7620[1]), .I2(n271_adj_4572), 
            .I3(n24461), .O(n7612[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3456_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3456_4 (.CI(n24461), .I0(n7620[1]), .I1(n271_adj_4572), 
            .CO(n24462));
    SB_LUT4 add_3456_3_lut (.I0(GND_net), .I1(n7620[0]), .I2(n198_adj_4573), 
            .I3(n24460), .O(n7612[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3456_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3456_3 (.CI(n24460), .I0(n7620[0]), .I1(n198_adj_4573), 
            .CO(n24461));
    SB_LUT4 add_3456_2_lut (.I0(GND_net), .I1(n56_adj_4574), .I2(n125_adj_4575), 
            .I3(GND_net), .O(n7612[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3456_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3456_2 (.CI(GND_net), .I0(n56_adj_4574), .I1(n125_adj_4575), 
            .CO(n24460));
    SB_LUT4 add_3455_8_lut (.I0(GND_net), .I1(n7612[5]), .I2(n560_adj_4576), 
            .I3(n24459), .O(n7603[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3455_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3455_7_lut (.I0(GND_net), .I1(n7612[4]), .I2(n487_adj_4577), 
            .I3(n24458), .O(n7603[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3455_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3455_7 (.CI(n24458), .I0(n7612[4]), .I1(n487_adj_4577), 
            .CO(n24459));
    SB_LUT4 add_3455_6_lut (.I0(GND_net), .I1(n7612[3]), .I2(n414_adj_4578), 
            .I3(n24457), .O(n7603[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3455_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3455_6 (.CI(n24457), .I0(n7612[3]), .I1(n414_adj_4578), 
            .CO(n24458));
    SB_LUT4 add_3455_5_lut (.I0(GND_net), .I1(n7612[2]), .I2(n341_adj_4579), 
            .I3(n24456), .O(n7603[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3455_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3455_5 (.CI(n24456), .I0(n7612[2]), .I1(n341_adj_4579), 
            .CO(n24457));
    SB_LUT4 add_3455_4_lut (.I0(GND_net), .I1(n7612[1]), .I2(n268_adj_4580), 
            .I3(n24455), .O(n7603[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3455_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3455_4 (.CI(n24455), .I0(n7612[1]), .I1(n268_adj_4580), 
            .CO(n24456));
    SB_LUT4 add_3455_3_lut (.I0(GND_net), .I1(n7612[0]), .I2(n195_adj_4581), 
            .I3(n24454), .O(n7603[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3455_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4386));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3455_3 (.CI(n24454), .I0(n7612[0]), .I1(n195_adj_4581), 
            .CO(n24455));
    SB_LUT4 add_3455_2_lut (.I0(GND_net), .I1(n53_adj_4582), .I2(n122_adj_4583), 
            .I3(GND_net), .O(n7603[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3455_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3455_2 (.CI(GND_net), .I0(n53_adj_4582), .I1(n122_adj_4583), 
            .CO(n24454));
    SB_LUT4 add_3454_9_lut (.I0(GND_net), .I1(n7603[6]), .I2(n630_adj_4584), 
            .I3(n24453), .O(n7593[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3454_8_lut (.I0(GND_net), .I1(n7603[5]), .I2(n557_adj_4585), 
            .I3(n24452), .O(n7593[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_8 (.CI(n24452), .I0(n7603[5]), .I1(n557_adj_4585), 
            .CO(n24453));
    SB_CARRY add_3443_2 (.CI(GND_net), .I0(n17_adj_4533), .I1(n86_adj_4534), 
            .CO(n24304));
    SB_LUT4 add_3454_7_lut (.I0(GND_net), .I1(n7603[4]), .I2(n484_adj_4586), 
            .I3(n24451), .O(n7593[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_7 (.CI(n24451), .I0(n7603[4]), .I1(n484_adj_4586), 
            .CO(n24452));
    SB_LUT4 add_3454_6_lut (.I0(GND_net), .I1(n7603[3]), .I2(n411_adj_4587), 
            .I3(n24450), .O(n7593[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_6 (.CI(n24450), .I0(n7603[3]), .I1(n411_adj_4587), 
            .CO(n24451));
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4587));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3454_5_lut (.I0(GND_net), .I1(n7603[2]), .I2(n338_adj_4539), 
            .I3(n24449), .O(n7593[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_5 (.CI(n24449), .I0(n7603[2]), .I1(n338_adj_4539), 
            .CO(n24450));
    SB_LUT4 add_3454_4_lut (.I0(GND_net), .I1(n7603[1]), .I2(n265_adj_4535), 
            .I3(n24448), .O(n7593[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4586));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3454_4 (.CI(n24448), .I0(n7603[1]), .I1(n265_adj_4535), 
            .CO(n24449));
    SB_LUT4 add_3454_3_lut (.I0(GND_net), .I1(n7603[0]), .I2(n192_adj_4519), 
            .I3(n24447), .O(n7593[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_3 (.CI(n24447), .I0(n7603[0]), .I1(n192_adj_4519), 
            .CO(n24448));
    SB_LUT4 add_3454_2_lut (.I0(GND_net), .I1(n50_adj_4518), .I2(n119_adj_4517), 
            .I3(GND_net), .O(n7593[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_2 (.CI(GND_net), .I0(n50_adj_4518), .I1(n119_adj_4517), 
            .CO(n24447));
    SB_LUT4 add_3453_10_lut (.I0(GND_net), .I1(n7593[7]), .I2(n700_adj_4516), 
            .I3(n24446), .O(n7582[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3453_9_lut (.I0(GND_net), .I1(n7593[6]), .I2(n627_adj_4515), 
            .I3(n24445), .O(n7582[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_15 (.CI(n24234), .I0(n7372[12]), .I1(n1026), .CO(n24235));
    SB_CARRY add_3453_9 (.CI(n24445), .I0(n7593[6]), .I1(n627_adj_4515), 
            .CO(n24446));
    SB_LUT4 add_3453_8_lut (.I0(GND_net), .I1(n7593[5]), .I2(n554_adj_4514), 
            .I3(n24444), .O(n7582[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3453_8 (.CI(n24444), .I0(n7593[5]), .I1(n554_adj_4514), 
            .CO(n24445));
    SB_LUT4 add_3453_7_lut (.I0(GND_net), .I1(n7593[4]), .I2(n481_adj_4513), 
            .I3(n24443), .O(n7582[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3453_7 (.CI(n24443), .I0(n7593[4]), .I1(n481_adj_4513), 
            .CO(n24444));
    SB_LUT4 add_3453_6_lut (.I0(GND_net), .I1(n7593[3]), .I2(n408_adj_4512), 
            .I3(n24442), .O(n7582[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3453_6 (.CI(n24442), .I0(n7593[3]), .I1(n408_adj_4512), 
            .CO(n24443));
    SB_LUT4 add_3453_5_lut (.I0(GND_net), .I1(n7593[2]), .I2(n335_adj_4511), 
            .I3(n24441), .O(n7582[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3453_5 (.CI(n24441), .I0(n7593[2]), .I1(n335_adj_4511), 
            .CO(n24442));
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4585));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4584));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4583));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4582));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3440_14_lut (.I0(GND_net), .I1(n7372[11]), .I2(n953), 
            .I3(n24233), .O(n7348[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3453_4_lut (.I0(GND_net), .I1(n7593[1]), .I2(n262_adj_4441), 
            .I3(n24440), .O(n7582[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_14 (.CI(n24233), .I0(n7372[11]), .I1(n953), .CO(n24234));
    SB_CARRY add_3453_4 (.CI(n24440), .I0(n7593[1]), .I1(n262_adj_4441), 
            .CO(n24441));
    SB_LUT4 add_3453_3_lut (.I0(GND_net), .I1(n7593[0]), .I2(n189_adj_4438), 
            .I3(n24439), .O(n7582[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3453_3 (.CI(n24439), .I0(n7593[0]), .I1(n189_adj_4438), 
            .CO(n24440));
    SB_LUT4 add_3453_2_lut (.I0(GND_net), .I1(n47_adj_4428), .I2(n116_adj_4427), 
            .I3(GND_net), .O(n7582[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3453_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3453_2 (.CI(GND_net), .I0(n47_adj_4428), .I1(n116_adj_4427), 
            .CO(n24439));
    SB_LUT4 add_3452_11_lut (.I0(GND_net), .I1(n7582[8]), .I2(n770_adj_4425), 
            .I3(n24438), .O(n7570[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3452_10_lut (.I0(GND_net), .I1(n7582[7]), .I2(n697_adj_4424), 
            .I3(n24437), .O(n7570[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3442_21_lut (.I0(GND_net), .I1(n7417[18]), .I2(GND_net), 
            .I3(n24303), .O(n7395[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_10 (.CI(n24437), .I0(n7582[7]), .I1(n697_adj_4424), 
            .CO(n24438));
    SB_LUT4 add_3452_9_lut (.I0(GND_net), .I1(n7582[6]), .I2(n624_adj_4423), 
            .I3(n24436), .O(n7570[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_9 (.CI(n24436), .I0(n7582[6]), .I1(n624_adj_4423), 
            .CO(n24437));
    SB_LUT4 add_3452_8_lut (.I0(GND_net), .I1(n7582[5]), .I2(n551_adj_4418), 
            .I3(n24435), .O(n7570[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_8 (.CI(n24435), .I0(n7582[5]), .I1(n551_adj_4418), 
            .CO(n24436));
    SB_LUT4 add_3452_7_lut (.I0(GND_net), .I1(n7582[4]), .I2(n478_adj_4415), 
            .I3(n24434), .O(n7570[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_7 (.CI(n24434), .I0(n7582[4]), .I1(n478_adj_4415), 
            .CO(n24435));
    SB_LUT4 add_3452_6_lut (.I0(GND_net), .I1(n7582[3]), .I2(n405_adj_4413), 
            .I3(n24433), .O(n7570[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_6 (.CI(n24433), .I0(n7582[3]), .I1(n405_adj_4413), 
            .CO(n24434));
    SB_LUT4 add_3452_5_lut (.I0(GND_net), .I1(n7582[2]), .I2(n332_adj_4412), 
            .I3(n24432), .O(n7570[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3442_20_lut (.I0(GND_net), .I1(n7417[17]), .I2(GND_net), 
            .I3(n24302), .O(n7395[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_5 (.CI(n24432), .I0(n7582[2]), .I1(n332_adj_4412), 
            .CO(n24433));
    SB_LUT4 add_3452_4_lut (.I0(GND_net), .I1(n7582[1]), .I2(n259_adj_4409), 
            .I3(n24431), .O(n7570[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3440_13_lut (.I0(GND_net), .I1(n7372[10]), .I2(n880), 
            .I3(n24232), .O(n7348[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_13 (.CI(n24232), .I0(n7372[10]), .I1(n880), .CO(n24233));
    SB_CARRY add_3452_4 (.CI(n24431), .I0(n7582[1]), .I1(n259_adj_4409), 
            .CO(n24432));
    SB_LUT4 add_3452_3_lut (.I0(GND_net), .I1(n7582[0]), .I2(n186_adj_4408), 
            .I3(n24430), .O(n7570[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_3 (.CI(n24430), .I0(n7582[0]), .I1(n186_adj_4408), 
            .CO(n24431));
    SB_LUT4 add_3452_2_lut (.I0(GND_net), .I1(n44_adj_4407), .I2(n113_adj_4406), 
            .I3(GND_net), .O(n7570[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_2 (.CI(GND_net), .I0(n44_adj_4407), .I1(n113_adj_4406), 
            .CO(n24430));
    SB_LUT4 add_3440_12_lut (.I0(GND_net), .I1(n7372[9]), .I2(n807), .I3(n24231), 
            .O(n7348[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3451_12_lut (.I0(GND_net), .I1(n7570[9]), .I2(n840_adj_4405), 
            .I3(n24429), .O(n7557[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3451_11_lut (.I0(GND_net), .I1(n7570[8]), .I2(n767_adj_4404), 
            .I3(n24428), .O(n7557[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_11 (.CI(n24428), .I0(n7570[8]), .I1(n767_adj_4404), 
            .CO(n24429));
    SB_LUT4 add_3451_10_lut (.I0(GND_net), .I1(n7570[7]), .I2(n694_adj_4403), 
            .I3(n24427), .O(n7557[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_10 (.CI(n24427), .I0(n7570[7]), .I1(n694_adj_4403), 
            .CO(n24428));
    SB_LUT4 add_3451_9_lut (.I0(GND_net), .I1(n7570[6]), .I2(n621_adj_4402), 
            .I3(n24426), .O(n7557[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_9 (.CI(n24426), .I0(n7570[6]), .I1(n621_adj_4402), 
            .CO(n24427));
    SB_LUT4 add_3451_8_lut (.I0(GND_net), .I1(n7570[5]), .I2(n548_adj_4401), 
            .I3(n24425), .O(n7557[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_20 (.CI(n24302), .I0(n7417[17]), .I1(GND_net), .CO(n24303));
    SB_CARRY add_3451_8 (.CI(n24425), .I0(n7570[5]), .I1(n548_adj_4401), 
            .CO(n24426));
    SB_LUT4 add_3451_7_lut (.I0(GND_net), .I1(n7570[4]), .I2(n475_adj_4400), 
            .I3(n24424), .O(n7557[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_7 (.CI(n24424), .I0(n7570[4]), .I1(n475_adj_4400), 
            .CO(n24425));
    SB_LUT4 add_3451_6_lut (.I0(GND_net), .I1(n7570[3]), .I2(n402_adj_4396), 
            .I3(n24423), .O(n7557[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_6 (.CI(n24423), .I0(n7570[3]), .I1(n402_adj_4396), 
            .CO(n24424));
    SB_LUT4 add_3451_5_lut (.I0(GND_net), .I1(n7570[2]), .I2(n329_adj_4395), 
            .I3(n24422), .O(n7557[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_5 (.CI(n24422), .I0(n7570[2]), .I1(n329_adj_4395), 
            .CO(n24423));
    SB_LUT4 add_3451_4_lut (.I0(GND_net), .I1(n7570[1]), .I2(n256_adj_4394), 
            .I3(n24421), .O(n7557[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_4 (.CI(n24421), .I0(n7570[1]), .I1(n256_adj_4394), 
            .CO(n24422));
    SB_LUT4 add_3451_3_lut (.I0(GND_net), .I1(n7570[0]), .I2(n183_adj_4393), 
            .I3(n24420), .O(n7557[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3451_3 (.CI(n24420), .I0(n7570[0]), .I1(n183_adj_4393), 
            .CO(n24421));
    SB_LUT4 add_3451_2_lut (.I0(GND_net), .I1(n41_adj_4392), .I2(n110_adj_4388), 
            .I3(GND_net), .O(n7557[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3451_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3442_19_lut (.I0(GND_net), .I1(n7417[16]), .I2(GND_net), 
            .I3(n24301), .O(n7395[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_12 (.CI(n24231), .I0(n7372[9]), .I1(n807), .CO(n24232));
    SB_CARRY add_3451_2 (.CI(GND_net), .I0(n41_adj_4392), .I1(n110_adj_4388), 
            .CO(n24420));
    SB_LUT4 add_3450_13_lut (.I0(GND_net), .I1(n7557[10]), .I2(n910_adj_4382), 
            .I3(n24419), .O(n7543[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3450_12_lut (.I0(GND_net), .I1(n7557[9]), .I2(n837_adj_4381), 
            .I3(n24418), .O(n7543[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_19 (.CI(n24301), .I0(n7417[16]), .I1(GND_net), .CO(n24302));
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4385));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4581));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4580));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4391));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3440_11_lut (.I0(GND_net), .I1(n7372[8]), .I2(n734), .I3(n24230), 
            .O(n7348[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_12 (.CI(n24418), .I0(n7557[9]), .I1(n837_adj_4381), 
            .CO(n24419));
    SB_CARRY add_3440_11 (.CI(n24230), .I0(n7372[8]), .I1(n734), .CO(n24231));
    SB_LUT4 add_3442_18_lut (.I0(GND_net), .I1(n7417[15]), .I2(GND_net), 
            .I3(n24300), .O(n7395[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3450_11_lut (.I0(GND_net), .I1(n7557[8]), .I2(n764_adj_4376), 
            .I3(n24417), .O(n7543[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_18 (.CI(n24300), .I0(n7417[15]), .I1(GND_net), .CO(n24301));
    SB_CARRY add_3450_11 (.CI(n24417), .I0(n7557[8]), .I1(n764_adj_4376), 
            .CO(n24418));
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4579));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4578));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4577));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4576));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4575));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4574));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4573));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4572));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3450_10_lut (.I0(GND_net), .I1(n7557[7]), .I2(n691_adj_4375), 
            .I3(n24416), .O(n7543[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_10 (.CI(n24416), .I0(n7557[7]), .I1(n691_adj_4375), 
            .CO(n24417));
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4571));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4570));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1482 (.I0(n6_adj_4507), .I1(\Kp[4] ), .I2(n7627[2]), 
            .I3(\PID_CONTROLLER.err [18]), .O(n7620[3]));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1482.LUT_INIT = 16'h965a;
    SB_LUT4 add_3450_9_lut (.I0(GND_net), .I1(n7557[6]), .I2(n618_adj_4374), 
            .I3(n24415), .O(n7543[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_9 (.CI(n24415), .I0(n7557[6]), .I1(n618_adj_4374), 
            .CO(n24416));
    SB_LUT4 add_3450_8_lut (.I0(GND_net), .I1(n7557[5]), .I2(n545_adj_4372), 
            .I3(n24414), .O(n7543[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_8 (.CI(n24414), .I0(n7557[5]), .I1(n545_adj_4372), 
            .CO(n24415));
    SB_LUT4 add_3450_7_lut (.I0(GND_net), .I1(n7557[4]), .I2(n472_adj_4371), 
            .I3(n24413), .O(n7543[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_7 (.CI(n24413), .I0(n7557[4]), .I1(n472_adj_4371), 
            .CO(n24414));
    SB_LUT4 add_3450_6_lut (.I0(GND_net), .I1(n7557[3]), .I2(n399_adj_4370), 
            .I3(n24412), .O(n7543[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_6 (.CI(n24412), .I0(n7557[3]), .I1(n399_adj_4370), 
            .CO(n24413));
    SB_LUT4 add_3450_5_lut (.I0(GND_net), .I1(n7557[2]), .I2(n326_adj_4369), 
            .I3(n24411), .O(n7543[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_5 (.CI(n24411), .I0(n7557[2]), .I1(n326_adj_4369), 
            .CO(n24412));
    SB_LUT4 add_3450_4_lut (.I0(GND_net), .I1(n7557[1]), .I2(n253_adj_4368), 
            .I3(n24410), .O(n7543[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_4 (.CI(n24410), .I0(n7557[1]), .I1(n253_adj_4368), 
            .CO(n24411));
    SB_LUT4 add_3450_3_lut (.I0(GND_net), .I1(n7557[0]), .I2(n180_adj_4367), 
            .I3(n24409), .O(n7543[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_3 (.CI(n24409), .I0(n7557[0]), .I1(n180_adj_4367), 
            .CO(n24410));
    SB_LUT4 add_3450_2_lut (.I0(GND_net), .I1(n38_adj_4366), .I2(n107_adj_4365), 
            .I3(GND_net), .O(n7543[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3450_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3450_2 (.CI(GND_net), .I0(n38_adj_4366), .I1(n107_adj_4365), 
            .CO(n24409));
    SB_LUT4 add_3449_14_lut (.I0(GND_net), .I1(n7543[11]), .I2(n980_adj_4363), 
            .I3(n24408), .O(n7528[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3449_13_lut (.I0(GND_net), .I1(n7543[10]), .I2(n907_adj_4362), 
            .I3(n24407), .O(n7528[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4267));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3449_13 (.CI(n24407), .I0(n7543[10]), .I1(n907_adj_4362), 
            .CO(n24408));
    SB_LUT4 add_3440_10_lut (.I0(GND_net), .I1(n7372[7]), .I2(n661), .I3(n24229), 
            .O(n7348[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_10 (.CI(n24229), .I0(n7372[7]), .I1(n661), .CO(n24230));
    SB_LUT4 add_3440_9_lut (.I0(GND_net), .I1(n7372[6]), .I2(n588), .I3(n24228), 
            .O(n7348[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3442_17_lut (.I0(GND_net), .I1(n7417[14]), .I2(GND_net), 
            .I3(n24299), .O(n7395[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_17 (.CI(n24299), .I0(n7417[14]), .I1(GND_net), .CO(n24300));
    SB_LUT4 add_3442_16_lut (.I0(GND_net), .I1(n7417[13]), .I2(n1105_adj_4360), 
            .I3(n24298), .O(n7395[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_16 (.CI(n24298), .I0(n7417[13]), .I1(n1105_adj_4360), 
            .CO(n24299));
    SB_LUT4 add_3442_15_lut (.I0(GND_net), .I1(n7417[12]), .I2(n1032_adj_4359), 
            .I3(n24297), .O(n7395[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3449_12_lut (.I0(GND_net), .I1(n7543[9]), .I2(n834_adj_4358), 
            .I3(n24406), .O(n7528[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_15 (.CI(n24297), .I0(n7417[12]), .I1(n1032_adj_4359), 
            .CO(n24298));
    SB_CARRY add_3440_9 (.CI(n24228), .I0(n7372[6]), .I1(n588), .CO(n24229));
    SB_LUT4 add_3440_8_lut (.I0(GND_net), .I1(n7372[5]), .I2(n515), .I3(n24227), 
            .O(n7348[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3442_14_lut (.I0(GND_net), .I1(n7417[11]), .I2(n959_adj_4357), 
            .I3(n24296), .O(n7395[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_12 (.CI(n24406), .I0(n7543[9]), .I1(n834_adj_4358), 
            .CO(n24407));
    SB_LUT4 add_3449_11_lut (.I0(GND_net), .I1(n7543[8]), .I2(n761_adj_4356), 
            .I3(n24405), .O(n7528[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_14 (.CI(n24296), .I0(n7417[11]), .I1(n959_adj_4357), 
            .CO(n24297));
    SB_CARRY add_3440_8 (.CI(n24227), .I0(n7372[5]), .I1(n515), .CO(n24228));
    SB_LUT4 add_3442_13_lut (.I0(GND_net), .I1(n7417[10]), .I2(n886_adj_4355), 
            .I3(n24295), .O(n7395[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3440_7_lut (.I0(GND_net), .I1(n7372[4]), .I2(n442), .I3(n24226), 
            .O(n7348[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_7 (.CI(n24226), .I0(n7372[4]), .I1(n442), .CO(n24227));
    SB_DFFE \PID_CONTROLLER.integral_1193__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[1]));   // verilog/motorControl.v(32[21:33])
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE \PID_CONTROLLER.integral_1193__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[2]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[3]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[4]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[5]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[6]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[7]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[8]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[9]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[10]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[11]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[12]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[13]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[14]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[15]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[16]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[17]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[18]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[19]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[20]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[21]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[22]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1193__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3624 ), .D(n28[23]));   // verilog/motorControl.v(32[21:33])
    SB_LUT4 i25369_4_lut (.I0(n21_adj_4391), .I1(n19_adj_4385), .I2(n17_adj_4386), 
            .I3(n9_adj_4384), .O(n31200));
    defparam i25369_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i25363_4_lut (.I0(n27_adj_4399), .I1(n15_adj_4387), .I2(n13_adj_4377), 
            .I3(n11_adj_4383), .O(n31194));
    defparam i25363_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3440_6_lut (.I0(GND_net), .I1(n7372[3]), .I2(n369), .I3(n24225), 
            .O(n7348[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_6 (.CI(n24225), .I0(n7372[3]), .I1(n369), .CO(n24226));
    SB_CARRY add_3442_13 (.CI(n24295), .I0(n7417[10]), .I1(n886_adj_4355), 
            .CO(n24296));
    SB_LUT4 add_3442_12_lut (.I0(GND_net), .I1(n7417[9]), .I2(n813_adj_4240), 
            .I3(n24294), .O(n7395[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_12 (.CI(n24294), .I0(n7417[9]), .I1(n813_adj_4240), 
            .CO(n24295));
    SB_LUT4 add_3442_11_lut (.I0(GND_net), .I1(n7417[8]), .I2(n740_adj_4239), 
            .I3(n24293), .O(n7395[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_11 (.CI(n24405), .I0(n7543[8]), .I1(n761_adj_4356), 
            .CO(n24406));
    SB_LUT4 add_3449_10_lut (.I0(GND_net), .I1(n7543[7]), .I2(n688), .I3(n24404), 
            .O(n7528[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_10 (.CI(n24404), .I0(n7543[7]), .I1(n688), .CO(n24405));
    SB_LUT4 add_3449_9_lut (.I0(GND_net), .I1(n7543[6]), .I2(n615), .I3(n24403), 
            .O(n7528[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_9 (.CI(n24403), .I0(n7543[6]), .I1(n615), .CO(n24404));
    SB_LUT4 add_3449_8_lut (.I0(GND_net), .I1(n7543[5]), .I2(n542), .I3(n24402), 
            .O(n7528[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_8 (.CI(n24402), .I0(n7543[5]), .I1(n542), .CO(n24403));
    SB_LUT4 add_3449_7_lut (.I0(GND_net), .I1(n7543[4]), .I2(n469), .I3(n24401), 
            .O(n7528[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_7 (.CI(n24401), .I0(n7543[4]), .I1(n469), .CO(n24402));
    SB_LUT4 add_3449_6_lut (.I0(GND_net), .I1(n7543[3]), .I2(n396), .I3(n24400), 
            .O(n7528[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18744_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n7638[0]));   // verilog/motorControl.v(34[17:23])
    defparam i18744_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_3449_6 (.CI(n24400), .I0(n7543[3]), .I1(n396), .CO(n24401));
    SB_LUT4 add_3449_5_lut (.I0(GND_net), .I1(n7543[2]), .I2(n323), .I3(n24399), 
            .O(n7528[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_5 (.CI(n24399), .I0(n7543[2]), .I1(n323), .CO(n24400));
    SB_LUT4 add_3449_4_lut (.I0(GND_net), .I1(n7543[1]), .I2(n250), .I3(n24398), 
            .O(n7528[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_4 (.CI(n24398), .I0(n7543[1]), .I1(n250), .CO(n24399));
    SB_LUT4 add_3449_3_lut (.I0(GND_net), .I1(n7543[0]), .I2(n177), .I3(n24397), 
            .O(n7528[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3449_3 (.CI(n24397), .I0(n7543[0]), .I1(n177), .CO(n24398));
    SB_LUT4 add_3449_2_lut (.I0(GND_net), .I1(n35), .I2(n104_adj_4211), 
            .I3(GND_net), .O(n7528[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3449_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_11 (.CI(n24293), .I0(n7417[8]), .I1(n740_adj_4239), 
            .CO(n24294));
    SB_LUT4 add_3440_5_lut (.I0(GND_net), .I1(n7372[2]), .I2(n296), .I3(n24224), 
            .O(n7348[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_5 (.CI(n24224), .I0(n7372[2]), .I1(n296), .CO(n24225));
    SB_LUT4 add_3440_4_lut (.I0(GND_net), .I1(n7372[1]), .I2(n223), .I3(n24223), 
            .O(n7348[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_4 (.CI(n24223), .I0(n7372[1]), .I1(n223), .CO(n24224));
    SB_CARRY add_3449_2 (.CI(GND_net), .I0(n35), .I1(n104_adj_4211), .CO(n24397));
    SB_LUT4 i2_4_lut_adj_1483 (.I0(n4_adj_4505), .I1(\Kp[3] ), .I2(n7633[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n7627[2]));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1483.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4569));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1484 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12_adj_4588));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1484.LUT_INIT = 16'h9c50;
    SB_LUT4 add_3448_15_lut (.I0(GND_net), .I1(n7528[12]), .I2(n1050), 
            .I3(n24396), .O(n7512[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18680_4_lut (.I0(n7627[2]), .I1(\Kp[4] ), .I2(n6_adj_4507), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_4589));   // verilog/motorControl.v(34[17:23])
    defparam i18680_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1485 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_4590));   // verilog/motorControl.v(34[17:23])
    defparam i1_4_lut_adj_1485.LUT_INIT = 16'h6ca0;
    SB_LUT4 i18711_4_lut (.I0(n7633[1]), .I1(\Kp[3] ), .I2(n4_adj_4505), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_4591));   // verilog/motorControl.v(34[17:23])
    defparam i18711_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_3448_14_lut (.I0(GND_net), .I1(n7528[11]), .I2(n977), 
            .I3(n24395), .O(n7512[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_14 (.CI(n24395), .I0(n7528[11]), .I1(n977), .CO(n24396));
    SB_LUT4 add_3448_13_lut (.I0(GND_net), .I1(n7528[10]), .I2(n904), 
            .I3(n24394), .O(n7512[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_13 (.CI(n24394), .I0(n7528[10]), .I1(n904), .CO(n24395));
    SB_LUT4 add_3448_12_lut (.I0(GND_net), .I1(n7528[9]), .I2(n831), .I3(n24393), 
            .O(n7512[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18746_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n23275));   // verilog/motorControl.v(34[17:23])
    defparam i18746_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1486 (.I0(n6_adj_4591), .I1(n11_adj_4590), .I2(n8_adj_4589), 
            .I3(n12_adj_4588), .O(n18_adj_4592));   // verilog/motorControl.v(34[17:23])
    defparam i8_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_CARRY add_3448_12 (.CI(n24393), .I0(n7528[9]), .I1(n831), .CO(n24394));
    SB_LUT4 add_3442_10_lut (.I0(GND_net), .I1(n7417[7]), .I2(n667_adj_4202), 
            .I3(n24292), .O(n7395[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_10 (.CI(n24292), .I0(n7417[7]), .I1(n667_adj_4202), 
            .CO(n24293));
    SB_LUT4 i3_4_lut_adj_1487 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13_adj_4593));   // verilog/motorControl.v(34[17:23])
    defparam i3_4_lut_adj_1487.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_3440_3_lut (.I0(GND_net), .I1(n7372[0]), .I2(n150), .I3(n24222), 
            .O(n7348[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3440_3 (.CI(n24222), .I0(n7372[0]), .I1(n150), .CO(n24223));
    SB_LUT4 i9_4_lut_adj_1488 (.I0(n13_adj_4593), .I1(n18_adj_4592), .I2(n23275), 
            .I3(n4_adj_4502), .O(n29930));   // verilog/motorControl.v(34[17:23])
    defparam i9_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 add_3448_11_lut (.I0(GND_net), .I1(n7528[8]), .I2(n758), .I3(n24392), 
            .O(n7512[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_11 (.CI(n24392), .I0(n7528[8]), .I1(n758), .CO(n24393));
    SB_LUT4 add_3442_9_lut (.I0(GND_net), .I1(n7417[6]), .I2(n594_adj_4194), 
            .I3(n24291), .O(n7395[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3448_10_lut (.I0(GND_net), .I1(n7528[7]), .I2(n685), .I3(n24391), 
            .O(n7512[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_9 (.CI(n24291), .I0(n7417[6]), .I1(n594_adj_4194), 
            .CO(n24292));
    SB_LUT4 add_3440_2_lut (.I0(GND_net), .I1(n8_adj_4190), .I2(n77), 
            .I3(GND_net), .O(n7348[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3440_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3442_8_lut (.I0(GND_net), .I1(n7417[5]), .I2(n521_adj_4188), 
            .I3(n24290), .O(n7395[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_8 (.CI(n24290), .I0(n7417[5]), .I1(n521_adj_4188), 
            .CO(n24291));
    SB_LUT4 add_3442_7_lut (.I0(GND_net), .I1(n7417[4]), .I2(n448_adj_4187), 
            .I3(n24289), .O(n7395[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_10 (.CI(n24391), .I0(n7528[7]), .I1(n685), .CO(n24392));
    SB_CARRY add_3440_2 (.CI(GND_net), .I0(n8_adj_4190), .I1(n77), .CO(n24222));
    SB_CARRY add_3442_7 (.CI(n24289), .I0(n7417[4]), .I1(n448_adj_4187), 
            .CO(n24290));
    SB_LUT4 add_3442_6_lut (.I0(GND_net), .I1(n7417[3]), .I2(n375_adj_4185), 
            .I3(n24288), .O(n7395[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_6 (.CI(n24288), .I0(n7417[3]), .I1(n375_adj_4185), 
            .CO(n24289));
    SB_LUT4 add_3442_5_lut (.I0(GND_net), .I1(n7417[2]), .I2(n302_adj_4184), 
            .I3(n24287), .O(n7395[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3448_9_lut (.I0(GND_net), .I1(n7528[6]), .I2(n612), .I3(n24390), 
            .O(n7512[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_9 (.CI(n24390), .I0(n7528[6]), .I1(n612), .CO(n24391));
    SB_LUT4 add_3448_8_lut (.I0(GND_net), .I1(n7528[5]), .I2(n539), .I3(n24389), 
            .O(n7512[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_8 (.CI(n24389), .I0(n7528[5]), .I1(n539), .CO(n24390));
    SB_LUT4 add_3448_7_lut (.I0(GND_net), .I1(n7528[4]), .I2(n466), .I3(n24388), 
            .O(n7512[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_7 (.CI(n24388), .I0(n7528[4]), .I1(n466), .CO(n24389));
    SB_LUT4 add_3448_6_lut (.I0(GND_net), .I1(n7528[3]), .I2(n393), .I3(n24387), 
            .O(n7512[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_6 (.CI(n24387), .I0(n7528[3]), .I1(n393), .CO(n24388));
    SB_LUT4 add_3448_5_lut (.I0(GND_net), .I1(n7528[2]), .I2(n320), .I3(n24386), 
            .O(n7512[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_5 (.CI(n24386), .I0(n7528[2]), .I1(n320), .CO(n24387));
    SB_LUT4 add_3448_4_lut (.I0(GND_net), .I1(n7528[1]), .I2(n247), .I3(n24385), 
            .O(n7512[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_5 (.CI(n24287), .I0(n7417[2]), .I1(n302_adj_4184), 
            .CO(n24288));
    SB_CARRY add_3448_4 (.CI(n24385), .I0(n7528[1]), .I1(n247), .CO(n24386));
    SB_LUT4 add_3442_4_lut (.I0(GND_net), .I1(n7417[1]), .I2(n229_adj_4182), 
            .I3(n24286), .O(n7395[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3448_3_lut (.I0(GND_net), .I1(n7528[0]), .I2(n174), .I3(n24384), 
            .O(n7512[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_4 (.CI(n24286), .I0(n7417[1]), .I1(n229_adj_4182), 
            .CO(n24287));
    SB_CARRY add_3448_3 (.CI(n24384), .I0(n7528[0]), .I1(n174), .CO(n24385));
    SB_LUT4 add_3448_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n7512[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3448_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3442_3_lut (.I0(GND_net), .I1(n7417[0]), .I2(n156), .I3(n24285), 
            .O(n7395[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3448_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n24384));
    SB_LUT4 add_3447_16_lut (.I0(GND_net), .I1(n7512[13]), .I2(n1120), 
            .I3(n24383), .O(n7495[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3447_15_lut (.I0(GND_net), .I1(n7512[12]), .I2(n1047), 
            .I3(n24382), .O(n7495[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_15 (.CI(n24382), .I0(n7512[12]), .I1(n1047), .CO(n24383));
    SB_CARRY add_3442_3 (.CI(n24285), .I0(n7417[0]), .I1(n156), .CO(n24286));
    SB_LUT4 add_3447_14_lut (.I0(GND_net), .I1(n7512[11]), .I2(n974), 
            .I3(n24381), .O(n7495[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_14 (.CI(n24381), .I0(n7512[11]), .I1(n974), .CO(n24382));
    SB_LUT4 add_3442_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n7395[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3442_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3447_13_lut (.I0(GND_net), .I1(n7512[10]), .I2(n901), 
            .I3(n24380), .O(n7495[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3442_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n24285));
    SB_CARRY add_3447_13 (.CI(n24380), .I0(n7512[10]), .I1(n901), .CO(n24381));
    SB_LUT4 add_3441_22_lut (.I0(GND_net), .I1(n7395[19]), .I2(GND_net), 
            .I3(n24284), .O(n7372[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3447_12_lut (.I0(GND_net), .I1(n7512[9]), .I2(n828), .I3(n24379), 
            .O(n7495[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_12 (.CI(n24379), .I0(n7512[9]), .I1(n828), .CO(n24380));
    SB_LUT4 add_3441_21_lut (.I0(GND_net), .I1(n7395[18]), .I2(GND_net), 
            .I3(n24283), .O(n7372[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3447_11_lut (.I0(GND_net), .I1(n7512[8]), .I2(n755), .I3(n24378), 
            .O(n7495[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_11 (.CI(n24378), .I0(n7512[8]), .I1(n755), .CO(n24379));
    SB_CARRY add_3441_21 (.CI(n24283), .I0(n7395[18]), .I1(GND_net), .CO(n24284));
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4568));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3447_10_lut (.I0(GND_net), .I1(n7512[7]), .I2(n682), .I3(n24377), 
            .O(n7495[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_10 (.CI(n24377), .I0(n7512[7]), .I1(n682), .CO(n24378));
    SB_LUT4 add_3447_9_lut (.I0(GND_net), .I1(n7512[6]), .I2(n609), .I3(n24376), 
            .O(n7495[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_9 (.CI(n24376), .I0(n7512[6]), .I1(n609), .CO(n24377));
    SB_LUT4 add_3447_8_lut (.I0(GND_net), .I1(n7512[5]), .I2(n536), .I3(n24375), 
            .O(n7495[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_8 (.CI(n24375), .I0(n7512[5]), .I1(n536), .CO(n24376));
    SB_LUT4 add_3447_7_lut (.I0(GND_net), .I1(n7512[4]), .I2(n463), .I3(n24374), 
            .O(n7495[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_7 (.CI(n24374), .I0(n7512[4]), .I1(n463), .CO(n24375));
    SB_LUT4 add_3447_6_lut (.I0(GND_net), .I1(n7512[3]), .I2(n390), .I3(n24373), 
            .O(n7495[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_6 (.CI(n24373), .I0(n7512[3]), .I1(n390), .CO(n24374));
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4567));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3447_5_lut (.I0(GND_net), .I1(n7512[2]), .I2(n317), .I3(n24372), 
            .O(n7495[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4566));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3447_5 (.CI(n24372), .I0(n7512[2]), .I1(n317), .CO(n24373));
    SB_LUT4 add_3447_4_lut (.I0(GND_net), .I1(n7512[1]), .I2(n244), .I3(n24371), 
            .O(n7495[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_20_lut (.I0(GND_net), .I1(n7395[17]), .I2(GND_net), 
            .I3(n24282), .O(n7372[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_4 (.CI(n24371), .I0(n7512[1]), .I1(n244), .CO(n24372));
    SB_LUT4 i25418_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n31249));   // verilog/motorControl.v(36[10:25])
    defparam i25418_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_3441_20 (.CI(n24282), .I0(n7395[17]), .I1(GND_net), .CO(n24283));
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_4497));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_3447_3_lut (.I0(GND_net), .I1(n7512[0]), .I2(n171), .I3(n24370), 
            .O(n7495[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4565));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4564));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3447_3 (.CI(n24370), .I0(n7512[0]), .I1(n171), .CO(n24371));
    SB_LUT4 add_3447_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n7495[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3447_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3447_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n24370));
    SB_LUT4 add_3446_17_lut (.I0(GND_net), .I1(n7495[14]), .I2(GND_net), 
            .I3(n24369), .O(n7477[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4563));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4562));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4561));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3441_19_lut (.I0(GND_net), .I1(n7395[16]), .I2(GND_net), 
            .I3(n24281), .O(n7372[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_16_lut (.I0(GND_net), .I1(n7495[13]), .I2(n1117), 
            .I3(n24368), .O(n7477[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4560));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4559));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4558));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_16 (.CI(n24368), .I0(n7495[13]), .I1(n1117), .CO(n24369));
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4557));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3446_15_lut (.I0(GND_net), .I1(n7495[12]), .I2(n1044), 
            .I3(n24367), .O(n7477[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_15 (.CI(n24367), .I0(n7495[12]), .I1(n1044), .CO(n24368));
    SB_LUT4 add_3446_14_lut (.I0(GND_net), .I1(n7495[11]), .I2(n971), 
            .I3(n24366), .O(n7477[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4556));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4555));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_14 (.CI(n24366), .I0(n7495[11]), .I1(n971), .CO(n24367));
    SB_LUT4 add_3446_13_lut (.I0(GND_net), .I1(n7495[10]), .I2(n898), 
            .I3(n24365), .O(n7477[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_19 (.CI(n24281), .I0(n7395[16]), .I1(GND_net), .CO(n24282));
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4554));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4553));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_13 (.CI(n24365), .I0(n7495[10]), .I1(n898), .CO(n24366));
    SB_LUT4 add_3441_18_lut (.I0(GND_net), .I1(n7395[15]), .I2(GND_net), 
            .I3(n24280), .O(n7372[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_12_lut (.I0(GND_net), .I1(n7495[9]), .I2(n825_adj_4594), 
            .I3(n24364), .O(n7477[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_12 (.CI(n24364), .I0(n7495[9]), .I1(n825_adj_4594), 
            .CO(n24365));
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4552));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4551));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4550));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3446_11_lut (.I0(GND_net), .I1(n7495[8]), .I2(n752_adj_4595), 
            .I3(n24363), .O(n7477[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4549));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4548));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_11 (.CI(n24363), .I0(n7495[8]), .I1(n752_adj_4595), 
            .CO(n24364));
    SB_LUT4 add_3446_10_lut (.I0(GND_net), .I1(n7495[7]), .I2(n679_adj_4596), 
            .I3(n24362), .O(n7477[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_10 (.CI(n24362), .I0(n7495[7]), .I1(n679_adj_4596), 
            .CO(n24363));
    SB_LUT4 add_3446_9_lut (.I0(GND_net), .I1(n7495[6]), .I2(n606_adj_4597), 
            .I3(n24361), .O(n7477[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_9 (.CI(n24361), .I0(n7495[6]), .I1(n606_adj_4597), 
            .CO(n24362));
    SB_LUT4 add_3446_8_lut (.I0(GND_net), .I1(n7495[5]), .I2(n533_adj_4598), 
            .I3(n24360), .O(n7477[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_8 (.CI(n24360), .I0(n7495[5]), .I1(n533_adj_4598), 
            .CO(n24361));
    SB_LUT4 add_3446_7_lut (.I0(GND_net), .I1(n7495[4]), .I2(n460_adj_4599), 
            .I3(n24359), .O(n7477[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_7 (.CI(n24359), .I0(n7495[4]), .I1(n460_adj_4599), 
            .CO(n24360));
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4547));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3446_6_lut (.I0(GND_net), .I1(n7495[3]), .I2(n387_adj_4600), 
            .I3(n24358), .O(n7477[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_6 (.CI(n24358), .I0(n7495[3]), .I1(n387_adj_4600), 
            .CO(n24359));
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4546));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4545));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3446_5_lut (.I0(GND_net), .I1(n7495[2]), .I2(n314_adj_4601), 
            .I3(n24357), .O(n7477[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4544));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_5 (.CI(n24357), .I0(n7495[2]), .I1(n314_adj_4601), 
            .CO(n24358));
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4543));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4542));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4541));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3446_4_lut (.I0(GND_net), .I1(n7495[1]), .I2(n241_adj_4602), 
            .I3(n24356), .O(n7477[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_4 (.CI(n24356), .I0(n7495[1]), .I1(n241_adj_4602), 
            .CO(n24357));
    SB_LUT4 add_3446_3_lut (.I0(GND_net), .I1(n7495[0]), .I2(n168_adj_4603), 
            .I3(n24355), .O(n7477[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4540));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4538));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_3 (.CI(n24355), .I0(n7495[0]), .I1(n168_adj_4603), 
            .CO(n24356));
    SB_LUT4 add_3446_2_lut (.I0(GND_net), .I1(n26_adj_4604), .I2(n95_adj_4605), 
            .I3(GND_net), .O(n7477[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4537));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_2 (.CI(GND_net), .I0(n26_adj_4604), .I1(n95_adj_4605), 
            .CO(n24355));
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4536));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3445_18_lut (.I0(GND_net), .I1(n7477[15]), .I2(GND_net), 
            .I3(n24354), .O(n7458[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3445_17_lut (.I0(GND_net), .I1(n7477[14]), .I2(GND_net), 
            .I3(n24353), .O(n7458[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_17 (.CI(n24353), .I0(n7477[14]), .I1(GND_net), .CO(n24354));
    SB_LUT4 add_3445_16_lut (.I0(GND_net), .I1(n7477[13]), .I2(n1114_adj_4606), 
            .I3(n24352), .O(n7458[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3445_16 (.CI(n24352), .I0(n7477[13]), .I1(n1114_adj_4606), 
            .CO(n24353));
    SB_LUT4 add_3445_15_lut (.I0(GND_net), .I1(n7477[12]), .I2(n1041), 
            .I3(n24351), .O(n7458[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3445_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4534));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4533));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4606));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4532));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4531));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4530));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4605));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4604));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4529));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4528));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4603));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4602));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4527));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4601));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4526));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4525));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4600));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4524));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4523));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4522));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4599));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4521));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4520));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4598));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4597));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4596));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4595));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4594));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_out_frame[11] , \data_out_frame[6] , GND_net, \data_out_frame[8] , 
            \data_out_frame[24] , \data_out_frame[10] , \data_out_frame[9] , 
            \data_out_frame[5] , rx_data, rx_data_ready, \data_out_frame[7] , 
            n15783, IntegralLimit, clk32MHz, n15782, \data_out_frame[12] , 
            n15781, \data_out_frame[14] , \data_out_frame[15] , \data_out_frame[16] , 
            \data_out_frame[17] , \data_out_frame[18] , \data_out_frame[19] , 
            \data_out_frame[23] , \data_out_frame[20] , \data_out_frame[13] , 
            n15780, n15779, n15778, n15777, n15776, n15775, \FRAME_MATCHER.state[1] , 
            n14318, n63, n3303, n15774, n15773, n15772, n4452, 
            \FRAME_MATCHER.state[0] , n14295, n23, \data_in_frame[2] , 
            \data_in_frame[1] , \data_in[3][3] , \data_in[0] , \data_in[2] , 
            \data_in[3][6] , \data_in[3][1] , \data_in[1] , \data_in[3][0] , 
            \data_in[3][4] , \data_in[3][2] , \data_in[3][7] , \data_out_frame[25] , 
            n771, n15771, n15770, n15769, \data_in_frame[11] , \data_in_frame[12] , 
            \data_in_frame[5] , setpoint, \data_in_frame[10] , n11643, 
            \data_in_frame[3] , \data_in_frame[8] , n4727, \data_in_frame[13] , 
            n15768, n15767, \data_in_frame[9] , \data_in_frame[4] , 
            \data_in_frame[6] , n15766, n15765, n4725, n29573, n63_adj_3, 
            n14309, n123, DE_c, LED_c, n14328, n32531, n32532, 
            n16232, PWMLimit, n16231, n16230, n16229, n16228, n16227, 
            n16226, n16225, n16224, n16223, n16222, n16221, n16220, 
            n16219, n16218, n16217, n16216, n16215, n16214, n16213, 
            n16212, n16211, n16210, n16209, control_mode, n16208, 
            n16207, n16206, n16205, n16204, n16199, tx_active, n27831, 
            n16023, neopxl_color, n16022, n16021, n16020, n16019, 
            n16018, n16017, n16016, n16015, n16014, n16013, n16012, 
            n16011, n16010, n16009, n16008, n16007, n16006, n16005, 
            n16004, n16003, n16002, n16001, n16000, n15999, n15998, 
            n15997, n15996, n15995, n15994, n15993, n15992, n15991, 
            n15990, n15989, n15988, n15987, n15986, n15985, n15984, 
            n15983, n15982, n15981, n15980, n15979, n15978, n15977, 
            n15976, n15975, n15974, n15973, n15972, n15971, n15970, 
            n15969, n15968, n15967, n15966, n15965, n15964, n15963, 
            n15962, n15961, n15960, n15959, n15958, n15957, n15956, 
            n15955, n15954, n15953, n15952, n15951, n15950, n15949, 
            n15948, n15947, n15946, n15945, n15944, n15943, n15942, 
            n15941, n15940, n15939, n15938, n15937, n15936, n15935, 
            n15934, n15933, n15932, n15931, n15930, n15929, n15928, 
            n15927, n15926, n15925, n15924, n15923, n15922, n15921, 
            n15920, n15919, n15918, n15917, n15916, n15915, n15914, 
            n15913, n15912, n15911, n15910, n15909, n15908, n15907, 
            n15906, n15905, n15904, n15903, n15902, n15901, \FRAME_MATCHER.state_31__N_2668[1] , 
            n15900, n15899, n15898, n15897, n15896, n15895, n8515, 
            n122, n5, n32898, n30290, n27243, n15719, n15894, 
            n15893, n15892, n15891, n15890, n15889, n15888, n15887, 
            n15886, n15885, n15884, n15883, n15882, n15881, n15880, 
            n15879, n15878, n15877, n15876, n15875, n15874, n15873, 
            n15872, n15871, n15870, n15869, n15868, n15867, n15866, 
            n15865, n15864, n15863, n15862, n15718, n15716, n15715, 
            \Ki[0] , n15714, \Kp[0] , n15713, n15861, n15860, n15859, 
            n15858, n15857, n15856, n15855, n15705, n15854, n15853, 
            n15852, n15851, n15850, n15849, n15848, \Ki[15] , n15847, 
            \Ki[14] , n15846, \Ki[13] , n15845, \Ki[12] , n15844, 
            \Ki[11] , n15843, \Ki[10] , n15842, \Ki[9] , n15841, 
            \Ki[8] , n15840, \Ki[7] , n15839, \Ki[6] , n15838, \Ki[5] , 
            n15837, \Ki[4] , n15836, \Ki[3] , n15835, \Ki[2] , n15834, 
            \Ki[1] , n15833, \Kp[15] , n15832, \Kp[14] , n15831, 
            \Kp[13] , n15830, \Kp[12] , n15829, \Kp[11] , n15828, 
            \Kp[10] , n15827, \Kp[9] , n15826, \Kp[8] , n15825, 
            \Kp[7] , n15824, \Kp[6] , n15823, \Kp[5] , n15822, \Kp[4] , 
            n15821, \Kp[3] , n15820, \Kp[2] , n15819, \Kp[1] , n15818, 
            n15817, n15815, n15814, n15813, n15812, n15811, n15810, 
            n15809, n15807, n15806, n15805, n15804, n15803, n15802, 
            n15801, n15800, n15799, n15798, n15797, n15796, n15795, 
            n15794, n15793, n15792, n15791, n15790, n15789, n15788, 
            n15787, n15786, n15785, n15784, n28749, n28775, VCC_net, 
            r_SM_Main, n8353, tx_o, \r_SM_Main_2__N_3493[1] , \r_Bit_Index[0] , 
            n4, n15730, n32553, n15722, tx_enable, n15548, n15643, 
            \r_SM_Main_2__N_3422[2] , r_SM_Main_adj_11, n27820, r_Rx_Data, 
            n19238, n4_adj_7, n4_adj_8, \r_Bit_Index[0]_adj_9 , n14287, 
            RX_N_2, n14282, n4_adj_10, n27405, n15764, n16203, n15712, 
            n15711, n15710, n15709, n15708, n15707, n15706) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[6] ;
    input GND_net;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[24] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]rx_data;
    output rx_data_ready;
    output [7:0]\data_out_frame[7] ;
    input n15783;
    output [23:0]IntegralLimit;
    input clk32MHz;
    input n15782;
    output [7:0]\data_out_frame[12] ;
    input n15781;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[13] ;
    input n15780;
    input n15779;
    input n15778;
    input n15777;
    input n15776;
    input n15775;
    output \FRAME_MATCHER.state[1] ;
    output n14318;
    output n63;
    output n3303;
    input n15774;
    input n15773;
    input n15772;
    output n4452;
    output \FRAME_MATCHER.state[0] ;
    output n14295;
    output n23;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[1] ;
    output \data_in[3][3] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[2] ;
    output \data_in[3][6] ;
    output \data_in[3][1] ;
    output [7:0]\data_in[1] ;
    output \data_in[3][0] ;
    output \data_in[3][4] ;
    output \data_in[3][2] ;
    output \data_in[3][7] ;
    output [7:0]\data_out_frame[25] ;
    output n771;
    input n15771;
    input n15770;
    input n15769;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[5] ;
    output [23:0]setpoint;
    output [7:0]\data_in_frame[10] ;
    output n11643;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[8] ;
    output n4727;
    output [7:0]\data_in_frame[13] ;
    input n15768;
    input n15767;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[6] ;
    input n15766;
    input n15765;
    output n4725;
    output n29573;
    output n63_adj_3;
    output n14309;
    output n123;
    output DE_c;
    output LED_c;
    output n14328;
    input n32531;
    input n32532;
    input n16232;
    output [23:0]PWMLimit;
    input n16231;
    input n16230;
    input n16229;
    input n16228;
    input n16227;
    input n16226;
    input n16225;
    input n16224;
    input n16223;
    input n16222;
    input n16221;
    input n16220;
    input n16219;
    input n16218;
    input n16217;
    input n16216;
    input n16215;
    input n16214;
    input n16213;
    input n16212;
    input n16211;
    input n16210;
    input n16209;
    output [7:0]control_mode;
    input n16208;
    input n16207;
    input n16206;
    input n16205;
    input n16204;
    input n16199;
    output tx_active;
    output n27831;
    input n16023;
    output [23:0]neopxl_color;
    input n16022;
    input n16021;
    input n16020;
    input n16019;
    input n16018;
    input n16017;
    input n16016;
    input n16015;
    input n16014;
    input n16013;
    input n16012;
    input n16011;
    input n16010;
    input n16009;
    input n16008;
    input n16007;
    input n16006;
    input n16005;
    input n16004;
    input n16003;
    input n16002;
    input n16001;
    input n16000;
    input n15999;
    input n15998;
    input n15997;
    input n15996;
    input n15995;
    input n15994;
    input n15993;
    input n15992;
    input n15991;
    input n15990;
    input n15989;
    input n15988;
    input n15987;
    input n15986;
    input n15985;
    input n15984;
    input n15983;
    input n15982;
    input n15981;
    input n15980;
    input n15979;
    input n15978;
    input n15977;
    input n15976;
    input n15975;
    input n15974;
    input n15973;
    input n15972;
    input n15971;
    input n15970;
    input n15969;
    input n15968;
    input n15967;
    input n15966;
    input n15965;
    input n15964;
    input n15963;
    input n15962;
    input n15961;
    input n15960;
    input n15959;
    input n15958;
    input n15957;
    input n15956;
    input n15955;
    input n15954;
    input n15953;
    input n15952;
    input n15951;
    input n15950;
    input n15949;
    input n15948;
    input n15947;
    input n15946;
    input n15945;
    input n15944;
    input n15943;
    input n15942;
    input n15941;
    input n15940;
    input n15939;
    input n15938;
    input n15937;
    input n15936;
    input n15935;
    input n15934;
    input n15933;
    input n15932;
    input n15931;
    input n15930;
    input n15929;
    input n15928;
    input n15927;
    input n15926;
    input n15925;
    input n15924;
    input n15923;
    input n15922;
    input n15921;
    input n15920;
    input n15919;
    input n15918;
    input n15917;
    input n15916;
    input n15915;
    input n15914;
    input n15913;
    input n15912;
    input n15911;
    input n15910;
    input n15909;
    input n15908;
    input n15907;
    input n15906;
    input n15905;
    input n15904;
    input n15903;
    input n15902;
    input n15901;
    output \FRAME_MATCHER.state_31__N_2668[1] ;
    input n15900;
    input n15899;
    input n15898;
    input n15897;
    input n15896;
    input n15895;
    output n8515;
    output n122;
    output n5;
    output n32898;
    output n30290;
    input n27243;
    input n15719;
    input n15894;
    input n15893;
    input n15892;
    input n15891;
    input n15890;
    input n15889;
    input n15888;
    input n15887;
    input n15886;
    input n15885;
    input n15884;
    input n15883;
    input n15882;
    input n15881;
    input n15880;
    input n15879;
    input n15878;
    input n15877;
    input n15876;
    input n15875;
    input n15874;
    input n15873;
    input n15872;
    input n15871;
    input n15870;
    input n15869;
    input n15868;
    input n15867;
    input n15866;
    input n15865;
    input n15864;
    input n15863;
    input n15862;
    input n15718;
    input n15716;
    input n15715;
    output \Ki[0] ;
    input n15714;
    output \Kp[0] ;
    input n15713;
    input n15861;
    input n15860;
    input n15859;
    input n15858;
    input n15857;
    input n15856;
    input n15855;
    input n15705;
    input n15854;
    input n15853;
    input n15852;
    input n15851;
    input n15850;
    input n15849;
    input n15848;
    output \Ki[15] ;
    input n15847;
    output \Ki[14] ;
    input n15846;
    output \Ki[13] ;
    input n15845;
    output \Ki[12] ;
    input n15844;
    output \Ki[11] ;
    input n15843;
    output \Ki[10] ;
    input n15842;
    output \Ki[9] ;
    input n15841;
    output \Ki[8] ;
    input n15840;
    output \Ki[7] ;
    input n15839;
    output \Ki[6] ;
    input n15838;
    output \Ki[5] ;
    input n15837;
    output \Ki[4] ;
    input n15836;
    output \Ki[3] ;
    input n15835;
    output \Ki[2] ;
    input n15834;
    output \Ki[1] ;
    input n15833;
    output \Kp[15] ;
    input n15832;
    output \Kp[14] ;
    input n15831;
    output \Kp[13] ;
    input n15830;
    output \Kp[12] ;
    input n15829;
    output \Kp[11] ;
    input n15828;
    output \Kp[10] ;
    input n15827;
    output \Kp[9] ;
    input n15826;
    output \Kp[8] ;
    input n15825;
    output \Kp[7] ;
    input n15824;
    output \Kp[6] ;
    input n15823;
    output \Kp[5] ;
    input n15822;
    output \Kp[4] ;
    input n15821;
    output \Kp[3] ;
    input n15820;
    output \Kp[2] ;
    input n15819;
    output \Kp[1] ;
    input n15818;
    input n15817;
    input n15815;
    input n15814;
    input n15813;
    input n15812;
    input n15811;
    input n15810;
    input n15809;
    input n15807;
    input n15806;
    input n15805;
    input n15804;
    input n15803;
    input n15802;
    input n15801;
    input n15800;
    input n15799;
    input n15798;
    input n15797;
    input n15796;
    input n15795;
    input n15794;
    input n15793;
    input n15792;
    input n15791;
    input n15790;
    input n15789;
    input n15788;
    input n15787;
    input n15786;
    input n15785;
    input n15784;
    output n28749;
    output n28775;
    input VCC_net;
    output [2:0]r_SM_Main;
    output n8353;
    output tx_o;
    output \r_SM_Main_2__N_3493[1] ;
    output \r_Bit_Index[0] ;
    output n4;
    input n15730;
    input n32553;
    input n15722;
    output tx_enable;
    output n15548;
    output n15643;
    output \r_SM_Main_2__N_3422[2] ;
    output [2:0]r_SM_Main_adj_11;
    input n27820;
    output r_Rx_Data;
    output n19238;
    output n4_adj_7;
    output n4_adj_8;
    output \r_Bit_Index[0]_adj_9 ;
    output n14287;
    input RX_N_2;
    output n14282;
    output n4_adj_10;
    input n27405;
    input n15764;
    input n16203;
    input n15712;
    input n15711;
    input n15710;
    input n15709;
    input n15708;
    input n15707;
    input n15706;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n6, n27949, n28307, n28333, n28226, n28227, n28370, n30004, 
        n28288, n28014, n14895, n29701, n28324, n28003, n1581, 
        n28542, n1174, n1178;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    
    wire n15816, n27970, n28313, n26015, n26375, n28466, n28508, 
        n12, n1180, n28216, n14018, n12528, n15395, n14978, n28533, 
        n28485, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n28348, n24, n22, n28282, n18, n26, n26359, n15383, 
        n29447, n28295, n28548, n28210, n26281, n6_adj_3879, n29737, 
        n28536, n28086, n28, n14719, n28438, n38, n36, n42, 
        n40, n14401, n28511, n41, n26451, n39, n30149, n12524, 
        n28244, n1260, n28041, n10, n1291, n28165, n10_adj_3880, 
        n30022;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n16, n17, n31098, n31097, n16_adj_3881, n1265, n6_adj_3882, 
        n17_adj_3883, n25814, n25290, n31152, n31151, n28020, n16_adj_3884, 
        n17_adj_3885, n31116, n31115, n16_adj_3886, n17_adj_3887, 
        n31110, n31109, n16_adj_3888, n17_adj_3889, n31107, n31106, 
        n29994, n16_adj_3890, n17_adj_3891, n31104, n31103, n28213, 
        n8, n28120, n28376, n6_adj_3892, n15008, n28224, n28903, 
        n25712, n2_adj_3893, n23549, n2028, n2_adj_3894, n23548, 
        n2_adj_3895, n23547, n2_adj_3896, n23546, n2_adj_3897, n23545, 
        n2_adj_3898, n23544, n2_adj_3899, n23543, n2_adj_3900, n23542, 
        n2_adj_3901, n23541, n26471, n26444, n28204, n2_adj_3902, 
        n23540, n2_adj_3903, n23539, n2_adj_3904, n23538, n2_adj_3905, 
        n23537, n2_adj_3906, n23536, n2_adj_3907, n23535, n2_adj_3908, 
        n23534, n2649, n3_adj_3909, n2_adj_3910, n23533, n3_adj_3911, 
        n2_adj_3912, n23532, n2_adj_3913, n23531, n2_adj_3914, n23530, 
        n3_adj_3915, n2_adj_3916, n23529, n3_adj_3917, n3_adj_3918, 
        n2_adj_3919, n23528, n3_adj_3920, n3_adj_3921, n2_adj_3922, 
        n23527, n2_adj_3923, n23526, n3_adj_3924, n3_adj_3925, n3_adj_3926, 
        n3_adj_3927, n2_adj_3928, n23525, n3_adj_3929, n3_adj_3930, 
        n2_adj_3931, n23524, n3_adj_3932, n2_adj_3933, n23523, n2_adj_3934, 
        n23522, n3_adj_3935, n2_adj_3936, n23521, n3_adj_3937, n3_adj_3938, 
        n3_adj_3939, n3_adj_3940, n3_adj_3941, n2_adj_3942, n23520, 
        n3_adj_3943, n3_adj_3944, n3_adj_3945, n3_adj_3946, n3_adj_3947, 
        n3_adj_3948, n3_adj_3949, n2_adj_3950, n23519, n3_adj_3951, 
        n3_adj_3952;
    wire [7:0]n8825;
    
    wire n15481, n15614, n3_adj_3953, n3_adj_3954, n161, n28141, 
        n26279, n14352, n25280, n25, n16_adj_3955, n17_adj_3956, 
        n31101, n31100, n6_adj_3957, n5_c, n31008, n7, n31954, 
        n32008, n14, n32056, n31099, n6_adj_3958, n5_adj_3959, n7_adj_3960, 
        n31948, n32080, n14_adj_3961, n32062, n31102, n31353, n5_adj_3962, 
        n7_adj_3963, n32200, n32212, n14_adj_3964, n32068, n31105, 
        n31346, n5_adj_3965, n7_adj_3966, n32194, n32230, n14_adj_3967, 
        n32074, n31108, n31582, n5_adj_3968, n7_adj_3969, n32182, 
        n32164, n14_adj_3970, n32086, n31112, n6_adj_3971, n5_adj_3972, 
        n7_adj_3973, n32032, n32116, n14_adj_3974, n32092, n31150, 
        n6_adj_3975, n5_adj_3976, n7_adj_3977, n32026, n32014, n14_adj_3978, 
        n32044, n31089, n30398, n32206, n31585, n6_adj_3979, n5_adj_3980, 
        n7_adj_3981, n32002, n32188, n14_adj_3982, n32050, n31095, 
        n27, n26_adj_3983, n28_adj_3984, n14454, n28763;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n4626, n14279, n5_adj_3985, n6_adj_3986, n27796, n4561, 
        n28769, n9, n27187, n27833, n27846, n27189, n27847, n27191, 
        n27848, n27193, n27849, n27195, n27850, n27197, n27851, 
        n29088, n27159, n27852, n9_adj_3987, n27233, n27841, n27235, 
        n27842, n41_adj_3988, n1, n11605, n27027, n27843, n18546, 
        n14313, n4_c, n1_adj_3989, n14307, n4_adj_3990, n7_adj_3991, 
        n27237, n27844, n27203, n27845, n27199, n27853, n27201, 
        n27854, n27205, n27834, n27855, n27209, n27836, n19835, 
        n6_adj_3992, tx_transmit_N_3393, n27207, n27835, n27211, n27837, 
        n27213, n27838, n27215, n27839, n19144, n11873, n3_adj_3993, 
        n14316, n28168, n12_adj_3994, n6_adj_3995, n27139, n27840, 
        n8_adj_3996, n14174, n8_adj_3997, n14292;
    wire [0:0]n3505;
    wire [2:0]r_SM_Main_2__N_3496;
    
    wire n28649, n14304, n43, n9411, n30064, \FRAME_MATCHER.rx_data_ready_prev , 
        n18_adj_3998, n24_adj_3999, n27757, n22_adj_4000, n14030, 
        n26429, n6_adj_4001, n14548, n26_adj_4002, n15026;
    wire [31:0]\FRAME_MATCHER.state_31__N_2604 ;
    
    wire n14335, n44, n42_adj_4003, n43_adj_4004, n14738, n10_adj_4005, 
        n28034, n28414, n41_adj_4006, n40_adj_4007, n39_adj_4008, 
        n50, n45, n14158, n14_adj_4009, n15, n14_adj_4010, n14310, 
        n15_adj_4011, n10_adj_4012, n10_adj_4013, n14_adj_4014, n33;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n13, n10_adj_4015, n14_adj_4016, n14320, n18_adj_4017, n20, 
        n15_adj_4018, n28117, n28271, n28207, n20_adj_4019, n19, 
        n30349, n5_adj_4020, n14327, n77, n81, n7_adj_4021, n27219, 
        n9_adj_4022, n7_adj_4023, n26419, n29867, n28247, n29802, 
        n28233, n25305, n29643, n28423, n6_adj_4024, n29188, n28330, 
        n25268, n14060, n26270, n26288;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n14967;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n28364, n26343, n28518, n8_adj_4025, n7_adj_4026, n29713;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n28514, n28171, n28873, n28071, n27925, n26365, n6_adj_4027, 
        n28499, n14845, n28463, n26457, n28256, n10_adj_4028, n19172, 
        n28259, n28232, n26326, n2076, n28405, n30041, n28420, 
        n29699, n27905, n28479, n28253, n15279, n14_adj_4029, n14627, 
        n10_adj_4030, n28195, n28162, n39_adj_4031, n28476, n6_adj_4032, 
        n26455, n28432, n38_adj_4033, n26337, n36_adj_4034, n28451, 
        n26352, n28179, n37, n28530, n35, n4524, n15507, n44_adj_4035, 
        n14395, n14434, n28_adj_4036, n4_adj_4037, n1835, n43_adj_4038, 
        n32, n15253, n28408, n30, n31, n26341, n14437, n29, 
        n28502, n28426, n7_adj_4039, n26348, n26335, n6_adj_4040, 
        n28488, n14515, n15145, n26272, n16_adj_4041, n15_adj_4042, 
        n17_adj_4043, n14_adj_4044, n26491, n28198, n28075, n28367, 
        n28_adj_4045, n27994, n21, n14727, n28156, n20_adj_4046, 
        n18_adj_4047, n24_adj_4048, n29407, n30_adj_4049, n28104, 
        n25251, n31_adj_4050, n27908, n29_adj_4051, n32_adj_4052, 
        n28444, n25359, n20_adj_4053, n19_adj_4054, n29012, n21_adj_4055, 
        n14617, n14499, n28124, n4040, n29993, n31_adj_4056, n12002, 
        n4523, n14987, n27984, Kp_23__N_810, n12_adj_4057, n28030, 
        n28321, n28230, n14368, n28847, n14588, n15085, n8_adj_4058, 
        n27_adj_4059, n14756, n8_adj_4060, n28145, n30312, n14662, 
        n8_adj_4061, n28301, n19_adj_4062, n14593, n24_adj_4063, n14819, 
        n30_adj_4064, n14542, n8_adj_4065, n10_adj_4066, n14648, n25_adj_4067, 
        n31_adj_4068, n11435, n28101, n28851, n14_adj_4069, n19871, 
        n10_adj_4070;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n29704, n29748, n23580, n23579, n23578, n23577, n14164, 
        n23576, n23575, n14_adj_4071, n20_adj_4072, n22_adj_4073, 
        n21_adj_4074, n6_adj_4075, n10_adj_4076, n27894, n27747, n27859, 
        n14332, n14338, n26290, n23574, n7_adj_4077, n26304, n28241, 
        n28110, n30114, n27911, n25261, n10_adj_4078, n13958, n14931, 
        n29581, n28382;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n28539;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n27957, n14705, n14521, n15096, n28482, n27929;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n57, n27915, n28262, n28318, n28037, n64, n29381, n26346, 
        n68, n28393, n66, n28238, n28011, n28127, n67, n28189, 
        n28527, n65, n62, n10_adj_4079, n14357, n14687, n72, n28261, 
        n28185, n28235, n28061, n70, n28429, n27918, n28545, n71, 
        n69, n80, n28053, n8_adj_4080, n25004, n10_adj_4081, n73, 
        n14518, n25952, n28292, n29640, n26333, n25294, n28417, 
        n6_adj_4082, n16_adj_4083, n28457, n17_adj_4084, n15_adj_4085, 
        n28379, n15416, n10_adj_4086, n14612, n81_adj_4087, n12_adj_4088, 
        n74, n29577, n28133, n29657, n28095, n15111, n29658, n27981, 
        n12_adj_4089, n28027, n28201, n26318, n28385, n15048, n14_adj_4090, 
        n10_adj_4091, n14459, n28491, n15021, n28521, Kp_23__N_1201, 
        n28250, n28345, n6_adj_4092, n28880, n6_adj_4093, n28472, 
        n28080, n28285, n15015, Kp_23__N_973, n14908, n6_adj_4094, 
        n7_adj_4095, n29382, Kp_23__N_976, n27991, n14632, n12_adj_4096, 
        n15317, n14505, Kp_23__N_1446, n14344, n27963, n14561, n14_adj_4097, 
        n28114, n9_adj_4098, n29900, n12_adj_4099, n6_adj_4100, n6_adj_4101, 
        n26276, n29862, n26383, Kp_23__N_1094, n14645, Kp_23__N_1378, 
        n15_adj_4102, n14_adj_4103, n28441, n27960, n14363, n28402, 
        n10_adj_4104, n28083, n27932, n12_adj_4105, n27974, Kp_23__N_1443, 
        n10_adj_4106, n28493, n28221, n14_adj_4107, n10_adj_4108, 
        n28356, n15039, n10_adj_4109, n28068, n14693, n12_adj_4110, 
        n27988, n28373, n26397, n28802, n13989, n26296, n7_adj_4111, 
        n14942, n15114, n15034, n28057, n28469, n15247, n8_adj_4112, 
        n28089, Kp_23__N_868, n28496, n27946, n22_adj_4113, n19686, 
        n7_adj_4114, n8_adj_4115, n8_adj_4116, n27867;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n16191, n16192, n16193, n16194, n29733, n16195, n28209, 
        n16196, n28351, n25_adj_4117, n28298, n16_adj_4118, n27935, 
        n28454, n24_adj_4119, n16197, n16198, n28_adj_4120, n25278, 
        n28049, n28390, n26320, n14917, n18_adj_4121, n28411, n14493, 
        n24_adj_4122, n22_adj_4123, n26_adj_4124, n28265, n29131, 
        n27921, Kp_23__N_944, n6_adj_4126, n15336, n12761, n16_adj_4127, 
        n17_adj_4128, n15120, n28336, n3_adj_4129, n28361, Kp_23__N_979, 
        n8_adj_4130;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n16183, n16184, n28159, n6_adj_4131, Kp_23__N_1186, n28396, 
        n20_adj_4132, n19_adj_4133, n14638, n21_adj_4134, n14378, 
        n10_adj_4135, n6_adj_4136, n14536, n16185, n28017, n32227, 
        n28399, n6_adj_4137, n31966, n32221;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n28460, n16186, n16187, n16188, n16189, n12_adj_4138, n32215, 
        n32209, n6_adj_4139, n32203, n32197, n32610, n32191, n32612, 
        n32185, n28505, n28310, n10_adj_4140, n32179, n32613, n12_adj_4141, 
        n16190, n8_adj_4142, n16175, n32_adj_4143, n16176, n16177, 
        n32609, n32161, n12_adj_4144, n31972, n32155, n6_adj_4145, 
        n31978, n32149, n29711, n31984, n32143, n32598, n31990, 
        n32137, n14_adj_4146, n31996, n32131, n15_adj_4147, n32104, 
        n32125, n10_adj_4148, n30020, n32113, n9_adj_4149, n11, 
        n32101, n29270, n12_adj_4150;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n32089, n29351, n32083, n29325, n32077, n29156, n32071, 
        n29303, n32065, n16178, n1_adj_4151, n16179, n87, n88, 
        n28448, n16_adj_4152, n32059, n17_adj_4153, n32053, n29740, 
        n32047, n32041, n29675, n28896, n32029, n29177, n32023, 
        n22_adj_4154, n29624, n28_adj_4155, n32011, n29199, n19123, 
        n16180, n16181, n19125, n16182, n19127, n19157, n7_adj_4156, 
        n8_adj_4157, n8_adj_4158, n27906, n16167, n16168, n16169, 
        n16170, n16171, n6_adj_4159, n29496, n16172, n16173, n29910, 
        n15514, n16174, n8_adj_4160, n16159, n28293, n28105, n28199, 
        n18_adj_4161, n27137, n8_adj_4162, n8_adj_4163, n19636, n19638, 
        n19642, n19660, n8_adj_4164, n29468, n16160, n16161, n16162, 
        n16163, n16164, n16165, n16166, n14347, n15605, n29767, 
        n16151, n16152, n32005, n16153, n16154, n16155, n16156, 
        n16157, n16158, n19694, n27883, n16143, n16144, n16145, 
        n16146, n16147, n16148, n16149, n16150, n26_adj_4165, n27874, 
        n8_adj_4166, n16135, n16136, n16137, n16138, n16139, n16140, 
        n16141, n16142, n16127, n16128, n16129, n16130, n16131, 
        n16132, n16133, n16134, n16119, n16120, n16121, n16122, 
        n16123, n16124, n16125, n16126, n16111, n16112, n16113, 
        n16114, n16115, n16116, n30_adj_4167, n31999, n17_adj_4168, 
        n31993, n31987, n16117, n31981, n31975, n31969, n31963, 
        n4525, n16118, n16103, n31951, n4526, n31945, n16104, 
        n16105, n16106, n16107, n16108, n16109, n16110, n4527, 
        n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, 
        n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
        n4544, n4545, n4546, n4547, n16095, n16096, n16097, n16098, 
        n16099, n16100, n16101, n16102, n16094, n16093, n16092, 
        n16091, n16090, n16089, n16088, n16087, n16086, n16085, 
        n16084, n16083, n16082, n16081, n16080, n16079, n16078, 
        n16077, n16076, n16075, n16074, n16073, n16072, n16071, 
        n16070, n16069, n16068, n16067, n16066, n16065, n16064, 
        n16063, n16062, n16061, n16060, n16059, n16058, n16057, 
        n16056, n16055, n16054, n16053, n16052, n16051, n16050, 
        n16049, n16048, n16047, n16046, n16045, n16044, n16043, 
        n16042, n16041, n16040, n16039, n16038, n16037, n16036, 
        n16035, n16034, n16033, n16032, n16031, n16030, n16029, 
        n16028, n16027, n16026, n16025, n16024, n15717, n15808;
    
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n27949), .I1(\data_out_frame[8] [4]), .I2(n28307), 
            .I3(n6), .O(n28333));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut (.I0(n28226), .I1(n28227), .I2(n28370), .I3(\data_out_frame[24] [0]), 
            .O(n30004));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[6] [2]), 
            .I2(n28288), .I3(\data_out_frame[6] [4]), .O(n28014));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(n28014), .I1(n28333), .I2(n14895), .I3(GND_net), 
            .O(n29701));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[11] [2]), .I1(n28324), .I2(n28003), 
            .I3(\data_out_frame[9] [1]), .O(n1581));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_848 (.I0(n1581), .I1(n29701), .I2(GND_net), .I3(GND_net), 
            .O(n28542));
    defparam i1_2_lut_adj_848.LUT_INIT = 16'h9999;
    SB_LUT4 i386_2_lut (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1174));   // verilog/coms.v(72[16:27])
    defparam i386_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i389_2_lut (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1178));   // verilog/coms.v(73[16:27])
    defparam i389_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14052_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15816));   // verilog/coms.v(90[7:20])
    defparam i14052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_849 (.I0(\data_out_frame[9] [3]), .I1(n27970), 
            .I2(n1178), .I3(\data_out_frame[11] [5]), .O(n28313));
    defparam i3_4_lut_adj_849.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_850 (.I0(n26015), .I1(n26375), .I2(GND_net), 
            .I3(GND_net), .O(n28466));
    defparam i1_2_lut_adj_850.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut (.I0(n28466), .I1(n28508), .I2(\data_out_frame[11] [7]), 
            .I3(n28313), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(n1180), .I1(n12), .I2(n28542), .I3(n28216), 
            .O(n14018));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_851 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n12528));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_851.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_852 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n15395));
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_853 (.I0(\data_out_frame[6] [7]), .I1(n27970), 
            .I2(n15395), .I3(GND_net), .O(n14978));
    defparam i2_3_lut_adj_853.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n15783));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_854 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n27949));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_854.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_855 (.I0(\data_out_frame[8] [1]), .I1(n27949), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n28533));
    defparam i2_3_lut_adj_855.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_856 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28485));
    defparam i1_2_lut_adj_856.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n15782));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i10_4_lut (.I0(n28348), .I1(n14978), .I2(\data_out_frame[5] [5]), 
            .I3(\data_out_frame[12] [0]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n28485), .I1(\data_out_frame[5] [0]), .I2(\data_out_frame[7] [4]), 
            .I3(\data_out_frame[11] [5]), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n28282), .I1(n24), .I2(n18), .I3(n14018), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n26359), .I1(n26), .I2(n22), .I3(n15383), 
            .O(n29447));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_857 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n28295));
    defparam i2_3_lut_adj_857.LUT_INIT = 16'h9696;
    SB_LUT4 i392_2_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1180));   // verilog/coms.v(74[16:27])
    defparam i392_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28216));
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_859 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n28548));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_859.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_860 (.I0(\data_out_frame[10] [0]), .I1(n28548), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n28210));
    defparam i2_3_lut_adj_860.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_861 (.I0(\data_out_frame[7] [6]), .I1(n26281), 
            .I2(\data_out_frame[5] [4]), .I3(n6_adj_3879), .O(n29737));
    defparam i4_4_lut_adj_861.LUT_INIT = 16'h9669;
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n15781));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_862 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28536));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_863 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28086));
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h6666;
    SB_LUT4 i5_2_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut (.I0(n28536), .I1(n14719), .I2(n28438), .I3(n29737), 
            .O(n38));
    defparam i15_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_864 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[14] [6]), 
            .I2(n28086), .I3(\data_out_frame[15] [0]), .O(n36));
    defparam i13_4_lut_adj_864.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n28295), .I1(n38), .I2(n28), .I3(n29447), 
            .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[12] [4]), .O(n40));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(n12528), .I1(n36), .I2(n14401), .I3(n28511), 
            .O(n41));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[10] [4]), 
            .I2(\data_out_frame[14] [7]), .I3(n26451), .O(n39));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n30149));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_865 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n28282));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_865.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_866 (.I0(\data_out_frame[10] [5]), .I1(n28282), 
            .I2(\data_out_frame[8] [4]), .I3(n12524), .O(n14895));
    defparam i3_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_867 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[12] [5]), 
            .I2(n14895), .I3(GND_net), .O(n28244));
    defparam i2_3_lut_adj_867.LUT_INIT = 16'h9696;
    SB_LUT4 i472_2_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1260));   // verilog/coms.v(85[17:28])
    defparam i472_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_868 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15383));
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_869 (.I0(n15383), .I1(\data_out_frame[5] [6]), 
            .I2(n28041), .I3(\data_out_frame[5] [7]), .O(n10));
    defparam i4_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_LUT4 i503_2_lut (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1291));   // verilog/coms.v(71[16:27])
    defparam i503_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_870 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[9] [7]), .O(n28348));
    defparam i3_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_871 (.I0(\data_out_frame[5] [4]), .I1(n1291), .I2(\data_out_frame[10] [2]), 
            .I3(n28165), .O(n10_adj_3880));
    defparam i4_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[5] [6]), .I1(n10_adj_3880), .I2(\data_out_frame[8] [0]), 
            .I3(GND_net), .O(n30022));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25534_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31098));
    defparam i25534_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25501_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31097));
    defparam i25501_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3881));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_872 (.I0(n1265), .I1(n28348), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_3882));
    defparam i1_2_lut_adj_872.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3883));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_873 (.I0(n25814), .I1(n25290), .I2(n28041), .I3(n6_adj_3882), 
            .O(n26281));
    defparam i4_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 i25502_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31152));
    defparam i25502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25504_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31151));
    defparam i25504_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_874 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28020));
    defparam i1_2_lut_adj_874.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3884));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3885));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25511_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31116));
    defparam i25511_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_875 (.I0(\data_out_frame[8] [1]), .I1(n25814), 
            .I2(GND_net), .I3(GND_net), .O(n28165));
    defparam i1_2_lut_adj_875.LUT_INIT = 16'h6666;
    SB_LUT4 i25574_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31115));
    defparam i25574_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3886));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_876 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[6] [0]), .O(n14719));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_876.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3887));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25514_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31110));
    defparam i25514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25518_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31109));
    defparam i25518_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3888));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3889));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25521_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31107));
    defparam i25521_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25524_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31106));
    defparam i25524_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_877 (.I0(n26281), .I1(\data_out_frame[10] [1]), 
            .I2(n30022), .I3(GND_net), .O(n29994));
    defparam i2_3_lut_adj_877.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3890));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3891));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25525_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31104));
    defparam i25525_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25527_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31103));
    defparam i25527_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[14] [6]), 
            .I2(n28213), .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_878 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[14] [5]), 
            .I2(n8), .I3(\data_out_frame[12] [5]), .O(n28120));
    defparam i1_4_lut_adj_878.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_879 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28376));
    defparam i1_2_lut_adj_879.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_880 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[13] [0]), 
            .I2(n26451), .I3(n6_adj_3892), .O(n15008));
    defparam i4_4_lut_adj_880.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_881 (.I0(\data_out_frame[19] [3]), .I1(n15008), 
            .I2(n28376), .I3(n28120), .O(n28224));
    defparam i3_4_lut_adj_881.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_882 (.I0(\data_out_frame[19] [2]), .I1(n28224), 
            .I2(n28903), .I3(GND_net), .O(n25712));
    defparam i2_3_lut_adj_882.LUT_INIT = 16'h6969;
    SB_LUT4 add_43_33_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n23549), .O(n2_adj_3893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_32_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n23548), .O(n2_adj_3894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n23548), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n23549));
    SB_LUT4 add_43_31_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n23547), .O(n2_adj_3895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n23547), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n23548));
    SB_LUT4 add_43_30_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n23546), .O(n2_adj_3896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_30 (.CI(n23546), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n23547));
    SB_LUT4 add_43_29_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n23545), .O(n2_adj_3897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_29 (.CI(n23545), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n23546));
    SB_LUT4 add_43_28_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n23544), .O(n2_adj_3898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_28 (.CI(n23544), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n23545));
    SB_LUT4 add_43_27_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n23543), .O(n2_adj_3899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_27 (.CI(n23543), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n23544));
    SB_LUT4 add_43_26_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n23542), .O(n2_adj_3900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_26 (.CI(n23542), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n23543));
    SB_LUT4 add_43_25_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n23541), .O(n2_adj_3901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_883 (.I0(n26471), .I1(\data_out_frame[23] [6]), 
            .I2(n26444), .I3(n28226), .O(n28204));
    defparam i3_4_lut_adj_883.LUT_INIT = 16'h9669;
    SB_CARRY add_43_25 (.CI(n23541), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n23542));
    SB_LUT4 add_43_24_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n23540), .O(n2_adj_3902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n23540), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n23541));
    SB_LUT4 add_43_23_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n23539), .O(n2_adj_3903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n23539), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n23540));
    SB_LUT4 add_43_22_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n23538), .O(n2_adj_3904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_22 (.CI(n23538), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n23539));
    SB_LUT4 add_43_21_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n23537), .O(n2_adj_3905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_21 (.CI(n23537), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n23538));
    SB_LUT4 add_43_20_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n23536), .O(n2_adj_3906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n23536), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n23537));
    SB_LUT4 add_43_19_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n23535), .O(n2_adj_3907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_19 (.CI(n23535), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n23536));
    SB_LUT4 add_43_18_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n23534), .O(n2_adj_3908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3909));
    defparam select_338_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_18 (.CI(n23534), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n23535));
    SB_LUT4 add_43_17_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n23533), .O(n2_adj_3910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3911));
    defparam select_338_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_17 (.CI(n23533), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n23534));
    SB_LUT4 add_43_16_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n23532), .O(n2_adj_3912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n23532), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n23533));
    SB_LUT4 add_43_15_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n23531), .O(n2_adj_3913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_15 (.CI(n23531), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n23532));
    SB_LUT4 add_43_14_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n23530), .O(n2_adj_3914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3915));
    defparam select_338_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_14 (.CI(n23530), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n23531));
    SB_LUT4 add_43_13_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n23529), .O(n2_adj_3916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3917));
    defparam select_338_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_13 (.CI(n23529), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n23530));
    SB_LUT4 select_338_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3918));
    defparam select_338_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_12_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n23528), .O(n2_adj_3919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3920));
    defparam select_338_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_12 (.CI(n23528), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n23529));
    SB_LUT4 select_338_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3921));
    defparam select_338_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_11_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n23527), .O(n2_adj_3922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_11 (.CI(n23527), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n23528));
    SB_LUT4 add_43_10_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n23526), .O(n2_adj_3923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n23526), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n23527));
    SB_LUT4 select_338_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3924));
    defparam select_338_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3925));
    defparam select_338_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3926));
    defparam select_338_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3927));
    defparam select_338_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_9_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n23525), .O(n2_adj_3928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3929));
    defparam select_338_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3930));
    defparam select_338_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_9 (.CI(n23525), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n23526));
    SB_LUT4 add_43_8_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n23524), .O(n2_adj_3931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3932));
    defparam select_338_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_8 (.CI(n23524), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n23525));
    SB_LUT4 add_43_7_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n23523), .O(n2_adj_3933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n23523), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n23524));
    SB_LUT4 add_43_6_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n23522), .O(n2_adj_3934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3935));
    defparam select_338_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_6 (.CI(n23522), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n23523));
    SB_LUT4 add_43_5_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n23521), .O(n2_adj_3936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3937));
    defparam select_338_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3938));
    defparam select_338_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n15780));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_338_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3939));
    defparam select_338_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3940));
    defparam select_338_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_5 (.CI(n23521), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n23522));
    SB_LUT4 select_338_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3941));
    defparam select_338_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_4_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n23520), .O(n2_adj_3942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_4 (.CI(n23520), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n23521));
    SB_LUT4 select_338_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3943));
    defparam select_338_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3944));
    defparam select_338_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3945));
    defparam select_338_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3946));
    defparam select_338_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3947));
    defparam select_338_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3948));
    defparam select_338_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3949));
    defparam select_338_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_3_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n23519), .O(n2_adj_3950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_338_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3951));
    defparam select_338_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_338_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3952));
    defparam select_338_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n15481), .D(n8825[7]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n15481), .D(n8825[6]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n15481), .D(n8825[5]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n15481), .D(n8825[4]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n15779));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_338_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3953));
    defparam select_338_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_3 (.CI(n23519), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n23520));
    SB_LUT4 select_338_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3954));
    defparam select_338_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_2_lut (.I0(n2028), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n15778));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n23519));
    SB_LUT4 i9_4_lut (.I0(n28141), .I1(n26279), .I2(n14352), .I3(n25280), 
            .O(n25));   // verilog/coms.v(85[17:70])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3955));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3956));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25530_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31101));
    defparam i25530_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25532_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31100));
    defparam i25532_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3957));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut (.I0(n5_c), .I1(n6_adj_3957), 
            .I2(n31008), .I3(GND_net), .O(n7));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1539849_i1_3_lut (.I0(n31954), .I1(n32008), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14));
    defparam i1539849_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25535_2_lut (.I0(n32056), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31099));
    defparam i25535_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3958));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3959));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut (.I0(n5_adj_3959), 
            .I1(n6_adj_3958), .I2(n31008), .I3(GND_net), .O(n7_adj_3960));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1540452_i1_3_lut (.I0(n31948), .I1(n32080), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3961));
    defparam i1540452_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25531_2_lut (.I0(n32062), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31102));
    defparam i25531_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n31353));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3962));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_4_lut (.I0(n5_adj_3962), 
            .I1(byte_transmit_counter[0]), .I2(n31008), .I3(n31353), .O(n7_adj_3963));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1541055_i1_3_lut (.I0(n32200), .I1(n32212), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3964));
    defparam i1541055_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25526_2_lut (.I0(n32068), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31105));
    defparam i25526_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i25515_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n31346));   // verilog/coms.v(106[34:55])
    defparam i25515_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3965));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_4_lut (.I0(n5_adj_3965), 
            .I1(n31346), .I2(n31008), .I3(byte_transmit_counter[0]), .O(n7_adj_3966));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1541658_i1_3_lut (.I0(n32194), .I1(n32230), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3967));
    defparam i1541658_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25523_2_lut (.I0(n32074), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31108));
    defparam i25523_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i25749_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n31582));   // verilog/coms.v(106[34:55])
    defparam i25749_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3968));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_4_lut (.I0(n5_adj_3968), 
            .I1(n31582), .I2(n31008), .I3(byte_transmit_counter[0]), .O(n7_adj_3969));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1542261_i1_3_lut (.I0(n32182), .I1(n32164), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3970));
    defparam i1542261_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25507_2_lut (.I0(n32086), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31112));
    defparam i25507_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n6_adj_3971));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hb0bc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3972));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut (.I0(n5_adj_3972), 
            .I1(n6_adj_3971), .I2(n31008), .I3(GND_net), .O(n7_adj_3973));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1543467_i1_3_lut (.I0(n32032), .I1(n32116), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3974));
    defparam i1543467_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25564_2_lut (.I0(n32092), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31150));
    defparam i25564_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i25167_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n31008));   // verilog/coms.v(106[34:55])
    defparam i25167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i6_3_lut (.I0(\data_out_frame[5] [1]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n6_adj_3975));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3976));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut (.I0(n5_adj_3976), 
            .I1(n6_adj_3975), .I2(n31008), .I3(GND_net), .O(n7_adj_3977));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1538643_i1_3_lut (.I0(n32026), .I1(n32014), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3978));
    defparam i1538643_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25568_2_lut (.I0(n32044), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31089));
    defparam i25568_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i24567_4_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n30398));
    defparam i24567_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i25752_3_lut (.I0(n32206), .I1(n30398), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n31585));
    defparam i25752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n6_adj_3979));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hb0b3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3980));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_4_lut (.I0(n5_adj_3980), 
            .I1(n6_adj_3979), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n7_adj_3981));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1539246_i1_3_lut (.I0(n32002), .I1(n32188), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3982));
    defparam i1539246_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25541_2_lut (.I0(n32050), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n31095));
    defparam i25541_2_lut.LUT_INIT = 16'h2222;
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n15777));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n15776));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n15775));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_884 (.I0(n25), .I1(n27), .I2(n26_adj_3983), 
            .I3(n28_adj_3984), .O(n14454));   // verilog/coms.v(85[17:70])
    defparam i15_4_lut_adj_884.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(n28763), .I1(\FRAME_MATCHER.state [3]), .I2(n4626), 
            .I3(GND_net), .O(n14279));
    defparam i1_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i26087_4_lut (.I0(n14279), .I1(n4626), .I2(n5_adj_3985), .I3(n6_adj_3986), 
            .O(n27796));
    defparam i26087_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i26042_4_lut (.I0(n28763), .I1(\FRAME_MATCHER.state [3]), .I2(n4561), 
            .I3(n4626), .O(n28769));
    defparam i26042_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i26039_2_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4561));   // verilog/coms.v(145[4] 299[11])
    defparam i26039_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_885 (.I0(\FRAME_MATCHER.state [29]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27187));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_886 (.I0(\FRAME_MATCHER.state [29]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27846));
    defparam i1_2_lut_adj_886.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_887 (.I0(\FRAME_MATCHER.state [28]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27189));
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_888 (.I0(\FRAME_MATCHER.state [28]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27847));
    defparam i1_2_lut_adj_888.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_889 (.I0(\FRAME_MATCHER.state [27]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27191));
    defparam i1_2_lut_adj_889.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_890 (.I0(\FRAME_MATCHER.state [27]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27848));
    defparam i1_2_lut_adj_890.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_891 (.I0(\FRAME_MATCHER.state [26]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27193));
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_892 (.I0(\FRAME_MATCHER.state [26]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27849));
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_893 (.I0(\FRAME_MATCHER.state [25]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27195));
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_894 (.I0(\FRAME_MATCHER.state [25]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27850));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_895 (.I0(\FRAME_MATCHER.state [24]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27197));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_896 (.I0(\FRAME_MATCHER.state [24]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27851));
    defparam i1_2_lut_adj_896.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_897 (.I0(\FRAME_MATCHER.state [23]), .I1(n29088), 
            .I2(GND_net), .I3(GND_net), .O(n27159));
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\FRAME_MATCHER.state [23]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27852));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_899 (.I0(\FRAME_MATCHER.state [22]), .I1(n9_adj_3987), 
            .I2(GND_net), .I3(GND_net), .O(n27233));
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\FRAME_MATCHER.state [22]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27841));
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\FRAME_MATCHER.state [21]), .I1(n9_adj_3987), 
            .I2(GND_net), .I3(GND_net), .O(n27235));
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_902 (.I0(\FRAME_MATCHER.state [21]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27842));
    defparam i1_2_lut_adj_902.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n41_adj_3988), .I1(n14318), .I2(n1), .I3(n11605), 
            .O(n29088));   // verilog/coms.v(115[11:12])
    defparam i2_4_lut.LUT_INIT = 16'hfbfa;
    SB_LUT4 i1_2_lut_adj_903 (.I0(\FRAME_MATCHER.state [20]), .I1(n29088), 
            .I2(GND_net), .I3(GND_net), .O(n27027));
    defparam i1_2_lut_adj_903.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\FRAME_MATCHER.state [20]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27843));
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_905 (.I0(n63), .I1(n18546), .I2(n14313), .I3(GND_net), 
            .O(n4_c));   // verilog/coms.v(142[4] 144[7])
    defparam i1_3_lut_adj_905.LUT_INIT = 16'ha8a8;
    SB_LUT4 i2_3_lut_adj_906 (.I0(n1_adj_3989), .I1(n4_c), .I2(n3303), 
            .I3(GND_net), .O(n11605));   // verilog/coms.v(227[9:54])
    defparam i2_3_lut_adj_906.LUT_INIT = 16'h0808;
    SB_LUT4 i1_4_lut_adj_907 (.I0(n1), .I1(n14307), .I2(n4_adj_3990), 
            .I3(n7_adj_3991), .O(n9_adj_3987));
    defparam i1_4_lut_adj_907.LUT_INIT = 16'hbbba;
    SB_LUT4 i1_2_lut_adj_908 (.I0(\FRAME_MATCHER.state [19]), .I1(n9_adj_3987), 
            .I2(GND_net), .I3(GND_net), .O(n27237));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_909 (.I0(\FRAME_MATCHER.state [19]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27844));
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_910 (.I0(\FRAME_MATCHER.state [18]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27203));
    defparam i1_2_lut_adj_910.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_911 (.I0(\FRAME_MATCHER.state [18]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27845));
    defparam i1_2_lut_adj_911.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_912 (.I0(\FRAME_MATCHER.state [16]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27199));
    defparam i1_2_lut_adj_912.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\FRAME_MATCHER.state [16]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27853));
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_914 (.I0(\FRAME_MATCHER.state [15]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27201));
    defparam i1_2_lut_adj_914.LUT_INIT = 16'h8888;
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n15481), .D(n8825[3]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_915 (.I0(\FRAME_MATCHER.state [15]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27854));
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_916 (.I0(\FRAME_MATCHER.state [11]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27205));
    defparam i1_2_lut_adj_916.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_917 (.I0(\FRAME_MATCHER.state [11]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27834));
    defparam i1_2_lut_adj_917.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_918 (.I0(\FRAME_MATCHER.state [10]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27855));
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_919 (.I0(\FRAME_MATCHER.state [9]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27209));
    defparam i1_2_lut_adj_919.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\FRAME_MATCHER.state [9]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27836));
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h8888;
    SB_LUT4 i26052_2_lut (.I0(n19835), .I1(n6_adj_3992), .I2(GND_net), 
            .I3(GND_net), .O(tx_transmit_N_3393));
    defparam i26052_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_921 (.I0(\FRAME_MATCHER.state [8]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27207));
    defparam i1_2_lut_adj_921.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_922 (.I0(\FRAME_MATCHER.state [8]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27835));
    defparam i1_2_lut_adj_922.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\FRAME_MATCHER.state [7]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27211));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_924 (.I0(\FRAME_MATCHER.state [7]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27837));
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_925 (.I0(\FRAME_MATCHER.state [6]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27213));
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\FRAME_MATCHER.state [6]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27838));
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_927 (.I0(\FRAME_MATCHER.state [5]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27215));
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h8888;
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n15774));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n15773));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_928 (.I0(\FRAME_MATCHER.state [5]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27839));
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_929 (.I0(n19144), .I1(n11873), .I2(n3_adj_3993), 
            .I3(n14316), .O(n27833));
    defparam i1_4_lut_adj_929.LUT_INIT = 16'ha0a8;
    SB_LUT4 i5_4_lut_3_lut_4_lut (.I0(\data_out_frame[11] [7]), .I1(n28168), 
            .I2(\data_out_frame[14] [3]), .I3(\data_out_frame[16] [4]), 
            .O(n12_adj_3994));
    defparam i5_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_930 (.I0(n1), .I1(n14307), .I2(n4_adj_3990), 
            .I3(n6_adj_3995), .O(n9));
    defparam i1_4_lut_adj_930.LUT_INIT = 16'hbbba;
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n15772));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n15481), .D(n8825[2]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_931 (.I0(\FRAME_MATCHER.state [4]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n27139));
    defparam i1_2_lut_adj_931.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_932 (.I0(\FRAME_MATCHER.state [4]), .I1(n27833), 
            .I2(GND_net), .I3(GND_net), .O(n27840));
    defparam i1_2_lut_adj_932.LUT_INIT = 16'h8888;
    SB_LUT4 i14714_4_lut (.I0(n8_adj_3996), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n14174), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i14714_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i14715_4_lut (.I0(n8_adj_3997), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n14292), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i14715_4_lut.LUT_INIT = 16'h3230;
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3496[0]), .C(clk32MHz), 
            .D(n3505[0]), .R(n28763));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i49_4_lut (.I0(n28649), .I1(n14304), .I2(\FRAME_MATCHER.state [3]), 
            .I3(\FRAME_MATCHER.state [2]), .O(n43));
    defparam i49_4_lut.LUT_INIT = 16'h0735;
    SB_LUT4 i15263_3_lut_4_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(\FRAME_MATCHER.state[1] ), .I2(n14295), .I3(n14318), .O(n2649));
    defparam i15263_3_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_adj_933 (.I0(n9411), .I1(n23), .I2(GND_net), .I3(GND_net), 
            .O(n1));   // verilog/coms.v(227[6] 229[9])
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_934 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[1] [7]), .O(n30064));
    defparam i3_4_lut_adj_934.LUT_INIT = 16'hfffe;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_2_lut (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3998));
    defparam i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10_4_lut_adj_935 (.I0(\data_in_frame[1] [4]), .I1(n30064), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[2] [6]), .O(n24_adj_3999));
    defparam i10_4_lut_adj_935.LUT_INIT = 16'h0020;
    SB_LUT4 i8_4_lut_adj_936 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[1] [2]), 
            .I2(n27757), .I3(\data_in_frame[2] [1]), .O(n22_adj_4000));
    defparam i8_4_lut_adj_936.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut (.I0(n14030), .I1(\data_out_frame[20] [4]), .I2(\data_out_frame[20] [3]), 
            .I3(n26429), .O(n6_adj_4001));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_937 (.I0(\data_in_frame[1] [6]), .I1(n24_adj_3999), 
            .I2(n18_adj_3998), .I3(n14548), .O(n26_adj_4002));
    defparam i12_4_lut_adj_937.LUT_INIT = 16'h0080;
    SB_LUT4 i13_4_lut_adj_938 (.I0(n15026), .I1(n26_adj_4002), .I2(n22_adj_4000), 
            .I3(\data_in_frame[1] [1]), .O(\FRAME_MATCHER.state_31__N_2604 [3]));
    defparam i13_4_lut_adj_938.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_adj_939 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n14335));   // verilog/coms.v(161[5:29])
    defparam i1_2_lut_adj_939.LUT_INIT = 16'hbbbb;
    SB_LUT4 i18_4_lut_adj_940 (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [30]), 
            .I2(\FRAME_MATCHER.i [23]), .I3(\FRAME_MATCHER.i [24]), .O(n44));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut_adj_940.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_941 (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [15]), .O(n42_adj_4003));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut_adj_941.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_942 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [29]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [18]), .O(n43_adj_4004));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut_adj_942.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[13] [6]), .I1(n14738), .I2(n14018), 
            .I3(GND_net), .O(n10_adj_4005));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_943 (.I0(\data_out_frame[13] [6]), .I1(n14738), 
            .I2(n28034), .I3(\data_out_frame[16] [0]), .O(n28414));
    defparam i2_3_lut_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_944 (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [7]), .I3(\FRAME_MATCHER.i [20]), .O(n41_adj_4006));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut_adj_944.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [11]), .O(n40_adj_4007));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i [19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4008));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41_adj_4006), .I1(n43_adj_4004), .I2(n42_adj_4003), 
            .I3(n44), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_945 (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [8]), 
            .I2(\FRAME_MATCHER.i [17]), .I3(\FRAME_MATCHER.i [5]), .O(n45));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut_adj_945.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39_adj_4008), .I3(n40_adj_4007), 
            .O(n14292));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_946 (.I0(\FRAME_MATCHER.i [4]), .I1(n14292), .I2(GND_net), 
            .I3(GND_net), .O(n14174));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_946.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut_adj_947 (.I0(\data_in[3][3] ), .I1(\data_in[0] [7]), 
            .I2(n14158), .I3(GND_net), .O(n14_adj_4009));
    defparam i5_3_lut_adj_947.LUT_INIT = 16'hfdfd;
    SB_LUT4 i6_4_lut_adj_948 (.I0(\data_in[2] [1]), .I1(\data_in[0] [2]), 
            .I2(\data_in[3][6] ), .I3(\data_in[2] [3]), .O(n15));
    defparam i6_4_lut_adj_948.LUT_INIT = 16'hf7ff;
    SB_LUT4 i8_4_lut_adj_949 (.I0(n15), .I1(\data_in[3][1] ), .I2(n14_adj_4009), 
            .I3(\data_in[3] [5]), .O(n18546));
    defparam i8_4_lut_adj_949.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_adj_950 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4010));
    defparam i5_3_lut_adj_950.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_951 (.I0(\data_in[0] [6]), .I1(n14310), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_4011));
    defparam i6_4_lut_adj_951.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_952 (.I0(n15_adj_4011), .I1(\data_in[3][0] ), .I2(n14_adj_4010), 
            .I3(\data_in[2] [2]), .O(n14158));
    defparam i8_4_lut_adj_952.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_953 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4012));
    defparam i4_4_lut_adj_953.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_954 (.I0(\data_in[3][4] ), .I1(n10_adj_4012), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n14310));
    defparam i5_3_lut_adj_954.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [0]), .I1(\data_in[0] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4013));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_955 (.I0(\data_in[1] [2]), .I1(\data_in[1] [3]), 
            .I2(\data_in[3][2] ), .I3(\data_in[1] [6]), .O(n14_adj_4014));
    defparam i6_4_lut_adj_955.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut (.I0(\data_in[3][7] ), .I1(n14_adj_4014), .I2(n10_adj_4013), 
            .I3(\data_in[0] [5]), .O(n33));
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i5_4_lut_adj_956 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[0] [1]), .O(n13));
    defparam i5_4_lut_adj_956.LUT_INIT = 16'h2000;
    SB_LUT4 i2_2_lut_adj_957 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4015));
    defparam i2_2_lut_adj_957.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_958 (.I0(\data_in[0] [2]), .I1(\data_in[3][3] ), 
            .I2(\data_in[3][1] ), .I3(\data_in[0] [7]), .O(n14_adj_4016));
    defparam i6_4_lut_adj_958.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_959 (.I0(\data_in[3][6] ), .I1(n14_adj_4016), .I2(n10_adj_4015), 
            .I3(\data_in[2] [1]), .O(n14320));
    defparam i7_4_lut_adj_959.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_960 (.I0(\data_in[2] [4]), .I1(n14320), .I2(\data_in[1] [5]), 
            .I3(n14313), .O(n18_adj_4017));
    defparam i7_4_lut_adj_960.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_961 (.I0(\data_in[0] [6]), .I1(n18_adj_4017), .I2(\data_in[3][0] ), 
            .I3(n14310), .O(n20));
    defparam i9_4_lut_adj_961.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_962 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4018));
    defparam i4_2_lut_adj_962.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_963 (.I0(n15_adj_4018), .I1(n20), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n1_adj_3989));
    defparam i10_4_lut_adj_963.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_964 (.I0(\data_out_frame[20] [3]), .I1(n28117), 
            .I2(\data_out_frame[25] [0]), .I3(n28271), .O(n28207));
    defparam i2_3_lut_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_965 (.I0(n14158), .I1(n14320), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [5]), .O(n20_adj_4019));
    defparam i8_4_lut_adj_965.LUT_INIT = 16'hefff;
    SB_LUT4 i7_4_lut_adj_966 (.I0(\data_in[2] [5]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3][7] ), .I3(\data_in[2] [6]), .O(n19));
    defparam i7_4_lut_adj_966.LUT_INIT = 16'hfffd;
    SB_LUT4 i24518_4_lut (.I0(\data_in[2] [0]), .I1(\data_in[0] [1]), .I2(\data_in[3][2] ), 
            .I3(\data_in[1] [2]), .O(n30349));
    defparam i24518_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n30349), .I1(n19), .I2(n20_adj_4019), .I3(GND_net), 
            .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i14664_4_lut (.I0(n5_adj_4020), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i14664_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_967 (.I0(n11873), .I1(n14327), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_adj_967.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_968 (.I0(\FRAME_MATCHER.state [3]), .I1(n81), .I2(n41_adj_3988), 
            .I3(n77), .O(n7_adj_4021));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_4_lut_adj_969 (.I0(n14295), .I1(n7_adj_4021), .I2(n14335), 
            .I3(\FRAME_MATCHER.state_31__N_2604 [3]), .O(n27219));
    defparam i1_4_lut_adj_969.LUT_INIT = 16'hcdcc;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n15771));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_970 (.I0(n13), .I1(n9_adj_4022), .I2(\data_in_frame[0] [5]), 
            .I3(\data_in_frame[0] [6]), .O(n27757));
    defparam i7_4_lut_adj_970.LUT_INIT = 16'h0002;
    SB_LUT4 i2_2_lut_adj_971 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4023));
    defparam i2_2_lut_adj_971.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_972 (.I0(n7_adj_4023), .I1(n26419), .I2(n29867), 
            .I3(n28247), .O(n29802));
    defparam i4_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_973 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(n28233), .I3(n25305), .O(n29643));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_974 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[24] [7]), 
            .I2(n28423), .I3(n6_adj_4024), .O(n29188));
    defparam i4_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_975 (.I0(\data_out_frame[20] [4]), .I1(n28330), 
            .I2(n25268), .I3(GND_net), .O(n14060));
    defparam i2_3_lut_adj_975.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n15481), .D(n8825[1]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n15770));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_976 (.I0(n26471), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28247));
    defparam i1_2_lut_adj_976.LUT_INIT = 16'h9999;
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n15769));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_977 (.I0(n26270), .I1(n28330), .I2(\data_out_frame[24] [7]), 
            .I3(n6_adj_4001), .O(n26288));
    defparam i4_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_978 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [4]), 
            .I2(n14454), .I3(GND_net), .O(n14967));   // verilog/coms.v(72[16:41])
    defparam i2_3_lut_adj_978.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28364));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_980 (.I0(n26343), .I1(n14030), .I2(n28518), .I3(GND_net), 
            .O(n8_adj_4025));
    defparam i3_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_981 (.I0(n26288), .I1(n28207), .I2(n7_adj_4026), 
            .I3(n8_adj_4025), .O(n29713));
    defparam i2_4_lut_adj_981.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_982 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28514));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_983 (.I0(n28171), .I1(n28414), .I2(n28873), .I3(GND_net), 
            .O(n26343));
    defparam i2_3_lut_adj_983.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28071));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27925));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_986 (.I0(n26270), .I1(n26365), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4027));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_987 (.I0(\data_in_frame[5] [4]), .I1(n28499), .I2(n14845), 
            .I3(GND_net), .O(n28463));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_987.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_988 (.I0(n26429), .I1(n26457), .I2(n28256), .I3(n6_adj_4027), 
            .O(n25268));
    defparam i4_4_lut_adj_988.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_989 (.I0(n26365), .I1(\data_out_frame[20] [6]), 
            .I2(n28873), .I3(\data_out_frame[19] [0]), .O(n10_adj_4028));
    defparam i4_4_lut_adj_989.LUT_INIT = 16'h9669;
    SB_LUT4 i14645_2_lut_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(n161), .I2(n14295), .I3(n14318), .O(n19172));
    defparam i14645_2_lut_2_lut_4_lut_4_lut.LUT_INIT = 16'h08cc;
    SB_LUT4 i1_2_lut_adj_990 (.I0(n29867), .I1(n25305), .I2(GND_net), 
            .I3(GND_net), .O(n28259));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_991 (.I0(\data_out_frame[23] [2]), .I1(n25268), 
            .I2(GND_net), .I3(GND_net), .O(n28232));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_992 (.I0(n26326), .I1(n2076), .I2(n26365), .I3(n28405), 
            .O(n26457));
    defparam i3_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_993 (.I0(n30041), .I1(\data_out_frame[24] [6]), 
            .I2(\data_out_frame[24] [7]), .I3(GND_net), .O(n28271));
    defparam i2_3_lut_adj_993.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_994 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28420));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_995 (.I0(n29699), .I1(\data_out_frame[18] [3]), 
            .I2(\data_out_frame[18] [2]), .I3(GND_net), .O(n28171));
    defparam i2_3_lut_adj_995.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_996 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27905));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'h6666;
    SB_LUT4 i1288_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(85[17:28])
    defparam i1288_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_997 (.I0(n28479), .I1(n26015), .I2(n28253), .I3(n15279), 
            .O(n14_adj_4029));
    defparam i6_4_lut_adj_997.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_998 (.I0(\data_out_frame[16] [2]), .I1(n14_adj_4029), 
            .I2(n10_adj_4005), .I3(n14627), .O(n28873));
    defparam i7_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[16] [1]), .I1(n14627), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[18] [4]), .O(n10_adj_4030));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_999 (.I0(n28195), .I1(\data_out_frame[15] [4]), 
            .I2(n28162), .I3(n28873), .O(n39_adj_4031));
    defparam i16_4_lut_adj_999.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1000 (.I0(\data_out_frame[16] [1]), .I1(n14627), 
            .I2(\data_out_frame[13] [7]), .I3(n28476), .O(n6_adj_4032));
    defparam i1_2_lut_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1001 (.I0(n26455), .I1(n28466), .I2(\data_out_frame[16] [1]), 
            .I3(n28432), .O(n38_adj_4033));
    defparam i15_4_lut_adj_1001.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1002 (.I0(n29699), .I1(n26337), .I2(n28244), 
            .I3(\data_out_frame[16] [0]), .O(n36_adj_4034));
    defparam i13_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1003 (.I0(n28451), .I1(n26352), .I2(n28179), 
            .I3(n26281), .O(n37));
    defparam i14_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i12_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [3]), 
            .I2(n28530), .I3(GND_net), .O(n35));
    defparam i12_3_lut.LUT_INIT = 16'h9696;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n15507), .D(n4524));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i21_4_lut (.I0(n35), .I1(n37), .I2(n36_adj_4034), .I3(n38_adj_4033), 
            .O(n44_adj_4035));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1004 (.I0(n14395), .I1(\data_out_frame[19] [4]), 
            .I2(n14434), .I3(\data_out_frame[19] [5]), .O(n28_adj_4036));
    defparam i10_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n39_adj_4031), .I1(n4_adj_4037), .I2(n14401), 
            .I3(n1835), .O(n43_adj_4038));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1005 (.I0(n43_adj_4038), .I1(n28_adj_4036), .I2(\data_out_frame[18] [0]), 
            .I3(n44_adj_4035), .O(n32));
    defparam i14_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1006 (.I0(n15253), .I1(\data_out_frame[17] [3]), 
            .I2(n28408), .I3(\data_out_frame[17] [0]), .O(n30));
    defparam i12_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1007 (.I0(n28476), .I1(\data_out_frame[17] [4]), 
            .I2(n28376), .I3(\data_out_frame[18] [3]), .O(n31));
    defparam i13_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(\data_out_frame[19] [3]), .I1(n26341), .I2(n14437), 
            .I3(\data_out_frame[18] [1]), .O(n29));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1008 (.I0(n29), .I1(n31), .I2(n30), .I3(n32), 
            .O(n28502));
    defparam i17_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1009 (.I0(\data_out_frame[19] [0]), .I1(n28426), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4039));
    defparam i2_2_lut_adj_1009.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1010 (.I0(n7_adj_4039), .I1(\data_out_frame[18] [5]), 
            .I2(n26348), .I3(n28502), .O(n26335));
    defparam i4_4_lut_adj_1010.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1011 (.I0(n28502), .I1(\data_out_frame[18] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4040));
    defparam i2_2_lut_adj_1011.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(\data_out_frame[20] [7]), .I1(n26326), 
            .I2(n6_adj_4040), .I3(n28488), .O(n26365));
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n14515));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1014 (.I0(\data_out_frame[14] [1]), .I1(n29447), 
            .I2(n14895), .I3(GND_net), .O(n28253));
    defparam i2_3_lut_adj_1014.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1015 (.I0(\data_out_frame[9] [5]), .I1(n15145), 
            .I2(n26272), .I3(n28213), .O(n16_adj_4041));
    defparam i6_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1016 (.I0(\data_out_frame[7] [5]), .I1(n26375), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4042));
    defparam i5_2_lut_adj_1016.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1017 (.I0(\data_out_frame[12] [1]), .I1(n28253), 
            .I2(n28451), .I3(n28168), .O(n17_adj_4043));
    defparam i7_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1018 (.I0(\data_out_frame[16] [3]), .I1(n17_adj_4043), 
            .I2(n15_adj_4042), .I3(n16_adj_4041), .O(n28426));
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1019 (.I0(n28426), .I1(n15145), .I2(\data_out_frame[18] [3]), 
            .I3(\data_out_frame[15] [7]), .O(n14_adj_4044));
    defparam i6_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1020 (.I0(\data_out_frame[20] [5]), .I1(n14_adj_4044), 
            .I2(n10_adj_4030), .I3(n26491), .O(n26429));
    defparam i7_4_lut_adj_1020.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28198));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1022 (.I0(n28075), .I1(\data_out_frame[25] [1]), 
            .I2(n28367), .I3(n28198), .O(n28_adj_4045));   // verilog/coms.v(71[16:27])
    defparam i10_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1023 (.I0(n14515), .I1(\data_out_frame[20] [7]), 
            .I2(n27994), .I3(n28117), .O(n21));
    defparam i8_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(n14727), .I1(n28156), .I2(\data_out_frame[20] [0]), 
            .I3(GND_net), .O(n20_adj_4046));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1024 (.I0(n21), .I1(n26348), .I2(n18_adj_4047), 
            .I3(\data_out_frame[20] [6]), .O(n24_adj_4048));
    defparam i11_4_lut_adj_1024.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1025 (.I0(n26335), .I1(n24_adj_4048), .I2(n20_adj_4046), 
            .I3(n28171), .O(n29407));
    defparam i12_4_lut_adj_1025.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1026 (.I0(n29407), .I1(n28420), .I2(n26365), 
            .I3(n28271), .O(n30_adj_4049));   // verilog/coms.v(71[16:27])
    defparam i12_4_lut_adj_1026.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1027 (.I0(n28104), .I1(\data_out_frame[23] [7]), 
            .I2(n26419), .I3(n25251), .O(n31_adj_4050));   // verilog/coms.v(71[16:27])
    defparam i13_4_lut_adj_1027.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1028 (.I0(\data_out_frame[23] [1]), .I1(n28423), 
            .I2(n27908), .I3(n28204), .O(n29_adj_4051));   // verilog/coms.v(71[16:27])
    defparam i11_4_lut_adj_1028.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1029 (.I0(n29_adj_4051), .I1(n31_adj_4050), .I2(n30_adj_4049), 
            .I3(n32_adj_4052), .O(n28444));   // verilog/coms.v(71[16:27])
    defparam i17_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1030 (.I0(n26343), .I1(\data_out_frame[20] [4]), 
            .I2(n26429), .I3(GND_net), .O(n30041));
    defparam i2_3_lut_adj_1030.LUT_INIT = 16'h6969;
    SB_LUT4 i8_4_lut_adj_1031 (.I0(n30041), .I1(n28444), .I2(n25359), 
            .I3(n28256), .O(n20_adj_4053));
    defparam i8_4_lut_adj_1031.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1032 (.I0(n28232), .I1(n26471), .I2(\data_out_frame[24] [5]), 
            .I3(n28259), .O(n19_adj_4054));
    defparam i7_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1033 (.I0(n26457), .I1(\data_out_frame[23] [4]), 
            .I2(\data_out_frame[25] [0]), .I3(n29012), .O(n21_adj_4055));
    defparam i9_4_lut_adj_1033.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1034 (.I0(n14617), .I1(n14499), .I2(\data_in_frame[10] [1]), 
            .I3(GND_net), .O(n28124));
    defparam i2_3_lut_adj_1034.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1035 (.I0(\FRAME_MATCHER.state_31__N_2604 [3]), .I1(n4040), 
            .I2(\FRAME_MATCHER.state[1] ), .I3(GND_net), .O(n11643));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_adj_1035.LUT_INIT = 16'h8080;
    SB_LUT4 i11_3_lut_adj_1036 (.I0(n21_adj_4055), .I1(n19_adj_4054), .I2(n20_adj_4053), 
            .I3(GND_net), .O(n29993));
    defparam i11_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1037 (.I0(\FRAME_MATCHER.state[1] ), .I1(n31_adj_4056), 
            .I2(n12002), .I3(GND_net), .O(n4523));
    defparam i2_3_lut_adj_1037.LUT_INIT = 16'h0202;
    SB_LUT4 i3_4_lut_adj_1038 (.I0(n14987), .I1(n28438), .I2(n1180), .I3(\data_out_frame[14] [0]), 
            .O(n14627));
    defparam i3_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28476));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1040 (.I0(\data_in_frame[3] [6]), .I1(n27984), 
            .I2(Kp_23__N_810), .I3(\data_in_frame[1] [3]), .O(n12_adj_4057));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1041 (.I0(n28030), .I1(n28034), .I2(n28321), 
            .I3(n6_adj_4032), .O(n14030));
    defparam i4_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1042 (.I0(\data_in_frame[8] [1]), .I1(n12_adj_4057), 
            .I2(n28230), .I3(n14368), .O(n28847));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(n14030), .I1(n25359), .I2(GND_net), 
            .I3(GND_net), .O(n28117));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1044 (.I0(n28847), .I1(n14588), .I2(n15085), 
            .I3(n8_adj_4058), .O(n27_adj_4059));
    defparam i11_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i24482_4_lut (.I0(\data_in_frame[8] [0]), .I1(n14756), .I2(n8_adj_4060), 
            .I3(n28145), .O(n30312));
    defparam i24482_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_4_lut_adj_1045 (.I0(n26365), .I1(n26335), .I2(n26444), 
            .I3(\data_out_frame[23] [3]), .O(n29867));
    defparam i2_3_lut_4_lut_adj_1045.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1046 (.I0(n14499), .I1(n14662), .I2(n8_adj_4061), 
            .I3(n28301), .O(n19_adj_4062));
    defparam i3_4_lut_adj_1046.LUT_INIT = 16'hb77b;
    SB_LUT4 i14_4_lut_adj_1047 (.I0(n27_adj_4059), .I1(n14593), .I2(n24_adj_4063), 
            .I3(n14819), .O(n30_adj_4064));
    defparam i14_4_lut_adj_1047.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1048 (.I0(n14542), .I1(n8_adj_4065), .I2(n10_adj_4066), 
            .I3(n14648), .O(n25_adj_4067));
    defparam i9_4_lut_adj_1048.LUT_INIT = 16'hfeff;
    SB_LUT4 i15_4_lut_adj_1049 (.I0(n25_adj_4067), .I1(n30_adj_4064), .I2(n19_adj_4062), 
            .I3(n30312), .O(n31_adj_4056));
    defparam i15_4_lut_adj_1049.LUT_INIT = 16'hfeff;
    SB_LUT4 i1634_3_lut (.I0(n31_adj_4068), .I1(n31_adj_4056), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(GND_net), .O(n11435));
    defparam i1634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(n26365), .I1(n26335), .I2(\data_out_frame[23] [1]), 
            .I3(GND_net), .O(n28256));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1050 (.I0(n28101), .I1(n28367), .I2(\data_out_frame[24] [4]), 
            .I3(GND_net), .O(n28851));
    defparam i2_3_lut_adj_1050.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1051 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [0]), .O(n14_adj_4069));
    defparam i6_4_lut_adj_1051.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1052 (.I0(n9_adj_4022), .I1(n14_adj_4069), .I2(\data_in_frame[0] [5]), 
            .I3(\data_in_frame[0] [2]), .O(n12002));
    defparam i7_4_lut_adj_1052.LUT_INIT = 16'hfeff;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(71[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1053 (.I0(\FRAME_MATCHER.state[0] ), .I1(n12002), 
            .I2(n19871), .I3(\FRAME_MATCHER.state [3]), .O(n10_adj_4070));
    defparam i4_4_lut_adj_1053.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(\data_out_frame[9] [4]), .I1(n28313), 
            .I2(GND_net), .I3(GND_net), .O(n15145));
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'h6666;
    SB_LUT4 i26023_3_lut (.I0(n11435), .I1(n10_adj_4070), .I2(\FRAME_MATCHER.state [2]), 
            .I3(GND_net), .O(n15507));
    defparam i26023_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 mux_1051_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4523), .I3(GND_net), .O(n4524));
    defparam mux_1051_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1055 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[15] [4]), .I3(n28414), .O(n27994));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28321));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1057 (.I0(\data_out_frame[20] [2]), .I1(n28321), 
            .I2(n27994), .I3(n29704), .O(n25359));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1057.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1058 (.I0(\data_out_frame[19] [7]), .I1(n25359), 
            .I2(n29748), .I3(GND_net), .O(n29012));
    defparam i2_3_lut_adj_1058.LUT_INIT = 16'h6969;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n23580), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n23579), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1059 (.I0(\data_out_frame[24] [3]), .I1(n29012), 
            .I2(\data_out_frame[24] [4]), .I3(GND_net), .O(n28104));
    defparam i2_3_lut_adj_1059.LUT_INIT = 16'h6969;
    SB_CARRY add_3971_8 (.CI(n23579), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n23580));
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n23578), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_7 (.CI(n23578), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n23579));
    SB_LUT4 i14618_2_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n19144));
    defparam i14618_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n14307));   // verilog/coms.v(222[5:21])
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'hbbbb;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n23577), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_6 (.CI(n23577), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n23578));
    SB_LUT4 i2_3_lut_adj_1061 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n14164), .I3(GND_net), .O(n14295));   // verilog/coms.v(254[5:25])
    defparam i2_3_lut_adj_1061.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_out_frame[13] [5]), .I1(n26375), 
            .I2(GND_net), .I3(GND_net), .O(n26491));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n23576), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1063 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[15] [6]), .I3(n26455), .O(n28156));
    defparam i3_4_lut_adj_1063.LUT_INIT = 16'h9669;
    SB_CARRY add_3971_5 (.CI(n23576), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n23577));
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n23575), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_4 (.CI(n23575), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n23576));
    SB_LUT4 i3_4_lut_adj_1064 (.I0(n31_adj_4056), .I1(n14335), .I2(n27757), 
            .I3(n14316), .O(n4727));
    defparam i3_4_lut_adj_1064.LUT_INIT = 16'h0010;
    SB_LUT4 select_338_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2649), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_338_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_1065 (.I0(\FRAME_MATCHER.state [7]), .I1(\FRAME_MATCHER.state [5]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4071));   // verilog/coms.v(201[5:24])
    defparam i2_2_lut_adj_1065.LUT_INIT = 16'heeee;
    SB_LUT4 i8_4_lut_adj_1066 (.I0(\FRAME_MATCHER.state [6]), .I1(\FRAME_MATCHER.state [24]), 
            .I2(\FRAME_MATCHER.state [27]), .I3(\FRAME_MATCHER.state [23]), 
            .O(n20_adj_4072));   // verilog/coms.v(201[5:24])
    defparam i8_4_lut_adj_1066.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1067 (.I0(\FRAME_MATCHER.state [4]), .I1(n20_adj_4072), 
            .I2(n14_adj_4071), .I3(\FRAME_MATCHER.state [16]), .O(n22_adj_4073));   // verilog/coms.v(201[5:24])
    defparam i10_4_lut_adj_1067.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1068 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [22]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [21]), 
            .O(n21_adj_4074));   // verilog/coms.v(201[5:24])
    defparam i9_4_lut_adj_1068.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1069 (.I0(n21_adj_4074), .I1(\FRAME_MATCHER.state [28]), 
            .I2(n22_adj_4073), .I3(\FRAME_MATCHER.state [26]), .O(n6_adj_4075));
    defparam i1_4_lut_adj_1069.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1070 (.I0(\FRAME_MATCHER.state [18]), .I1(\FRAME_MATCHER.state [19]), 
            .I2(\FRAME_MATCHER.state [25]), .I3(\FRAME_MATCHER.state [30]), 
            .O(n10_adj_4076));
    defparam i4_4_lut_adj_1070.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1071 (.I0(\FRAME_MATCHER.state [20]), .I1(n10_adj_4076), 
            .I2(\FRAME_MATCHER.state [17]), .I3(GND_net), .O(n27894));
    defparam i5_3_lut_adj_1071.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1072 (.I0(\FRAME_MATCHER.state [8]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(\FRAME_MATCHER.state [11]), .I3(\FRAME_MATCHER.state [15]), 
            .O(n27747));
    defparam i3_4_lut_adj_1072.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1073 (.I0(\FRAME_MATCHER.state [10]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [14]), .I3(\FRAME_MATCHER.state [13]), 
            .O(n27859));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n14332));   // verilog/coms.v(146[5:9])
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1075 (.I0(n27859), .I1(n27747), .I2(n27894), 
            .I3(n6_adj_4075), .O(n14164));   // verilog/coms.v(201[5:24])
    defparam i4_4_lut_adj_1075.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1076 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n14338));   // verilog/coms.v(263[5:27])
    defparam i1_2_lut_adj_1076.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_1077 (.I0(\data_out_frame[18] [0]), .I1(n28156), 
            .I2(n14395), .I3(n26290), .O(n29748));
    defparam i3_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n14434));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n23574), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1079 (.I0(n7_adj_4077), .I1(n29748), .I2(n26304), 
            .I3(n28241), .O(n28101));
    defparam i4_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1080 (.I0(n28370), .I1(n28110), .I2(n28101), 
            .I3(GND_net), .O(n25251));
    defparam i2_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1081 (.I0(n25251), .I1(\data_out_frame[24] [2]), 
            .I2(\data_out_frame[24] [3]), .I3(GND_net), .O(n30114));
    defparam i2_3_lut_adj_1081.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1082 (.I0(\data_out_frame[13] [4]), .I1(n28324), 
            .I2(n27911), .I3(n25261), .O(n10_adj_4078));
    defparam i4_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1083 (.I0(n28295), .I1(n10_adj_4078), .I2(n13958), 
            .I3(GND_net), .O(n29699));
    defparam i5_3_lut_adj_1083.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1084 (.I0(n26290), .I1(n14931), .I2(\data_out_frame[17] [6]), 
            .I3(GND_net), .O(n26341));
    defparam i2_3_lut_adj_1084.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1085 (.I0(\data_out_frame[20] [0]), .I1(n26341), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n28241));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1085.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1086 (.I0(n14727), .I1(n28241), .I2(n14395), 
            .I3(GND_net), .O(n29581));
    defparam i2_3_lut_adj_1086.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1087 (.I0(n29581), .I1(\data_out_frame[24] [2]), 
            .I2(\data_out_frame[24] [1]), .I3(GND_net), .O(n27908));
    defparam i2_3_lut_adj_1087.LUT_INIT = 16'h6969;
    SB_CARRY add_3971_3 (.CI(n23574), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n23575));
    SB_LUT4 i1_2_lut_adj_1088 (.I0(n1581), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28030));
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1089 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4022));
    defparam i1_2_lut_adj_1089.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28382));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1091 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[18] [1]), .O(n28539));
    defparam i3_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1092 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n28499));
    defparam i2_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1093 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[16] [3]), 
            .I2(n14454), .I3(\data_in_frame[16] [2]), .O(n27957));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1094 (.I0(n14705), .I1(n14521), .I2(\data_in_frame[5] [4]), 
            .I3(\data_in_frame[7] [6]), .O(n14662));
    defparam i3_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(n14648), .I1(n14662), .I2(GND_net), 
            .I3(GND_net), .O(n15096));
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1096 (.I0(\data_in_frame[15] [4]), .I1(n28482), 
            .I2(\data_in_frame[15] [5]), .I3(GND_net), .O(n27929));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1096.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut_adj_1097 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[17] [0]), .I3(\data_in_frame[18] [5]), .O(n57));
    defparam i15_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1098 (.I0(n27915), .I1(n28262), .I2(n28318), 
            .I3(n28037), .O(n64));
    defparam i22_4_lut_adj_1098.LUT_INIT = 16'h9669;
    SB_LUT4 i26_4_lut (.I0(n29381), .I1(\data_in_frame[8] [5]), .I2(n15096), 
            .I3(n26346), .O(n68));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1099 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[17] [4]), 
            .I2(\data_in_frame[11] [3]), .I3(n28393), .O(n66));
    defparam i24_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1100 (.I0(n28238), .I1(n28011), .I2(n28127), 
            .I3(n27929), .O(n67));
    defparam i25_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(\data_in_frame[10] [1]), .I1(n28189), .I2(n28527), 
            .I3(n27957), .O(n65));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_2_lut (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n62));
    defparam i20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1101 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[19] [4]), 
            .I2(\data_in_frame[19] [2]), .I3(GND_net), .O(n10_adj_4079));
    defparam i3_3_lut_adj_1101.LUT_INIT = 16'h9696;
    SB_LUT4 i30_4_lut (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[10] [3]), 
            .I2(n14357), .I3(n14687), .O(n72));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n28261), .I1(n28185), .I2(n28235), .I3(n28061), 
            .O(n70));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n57), .I1(n28429), .I2(n27918), .I3(n28545), 
            .O(n71));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(\data_in_frame[18] [3]), .I1(n28499), .I2(n28539), 
            .I3(n28382), .O(n69));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i38_4_lut (.I0(n65), .I1(n67), .I2(n66), .I3(n68), .O(n80));
    defparam i38_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(n14931), .I1(\data_out_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28053));
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1103 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[17] [4]), 
            .I2(n28053), .I3(n26304), .O(n28370));
    defparam i1_4_lut_adj_1103.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_1104 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[24] [1]), 
            .I2(n25712), .I3(GND_net), .O(n8_adj_4080));
    defparam i3_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n15768));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1105 (.I0(n28110), .I1(n30004), .I2(n8_adj_4080), 
            .I3(n28227), .O(n25004));
    defparam i3_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1106 (.I0(\data_out_frame[13] [2]), .I1(n28333), 
            .I2(n28003), .I3(\data_out_frame[9] [0]), .O(n10_adj_4081));
    defparam i4_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(n29704), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28179));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h9999;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3393), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31_4_lut (.I0(\data_in_frame[16] [7]), .I1(n62), .I2(\data_in_frame[13] [3]), 
            .I3(\data_in_frame[16] [6]), .O(n73));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[17] [4]), .I1(n15253), 
            .I2(GND_net), .I3(GND_net), .O(n14518));
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1109 (.I0(\data_out_frame[19] [5]), .I1(n14518), 
            .I2(\data_out_frame[17] [3]), .I3(n15008), .O(n14727));
    defparam i3_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_out_frame[23] [7]), .I1(n14727), 
            .I2(GND_net), .I3(GND_net), .O(n28227));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_out_frame[24] [0]), .I1(n25952), 
            .I2(GND_net), .I3(GND_net), .O(n28075));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(n25712), .I1(\data_out_frame[23] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26419));
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1113 (.I0(n26419), .I1(n28292), .I2(n28075), 
            .I3(\data_out_frame[25] [7]), .O(n29640));
    defparam i3_4_lut_adj_1113.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1114 (.I0(\data_out_frame[12] [7]), .I1(n29701), 
            .I2(\data_out_frame[13] [1]), .I3(GND_net), .O(n26333));
    defparam i2_3_lut_adj_1114.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1115 (.I0(\data_out_frame[15] [2]), .I1(n25294), 
            .I2(n26333), .I3(\data_out_frame[13] [0]), .O(n26304));
    defparam i3_4_lut_adj_1115.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(n26304), .I1(n30149), .I2(GND_net), 
            .I3(GND_net), .O(n28162));
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14437));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1118 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(n26429), .I3(GND_net), .O(n28417));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1118.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1119 (.I0(n14437), .I1(n28903), .I2(\data_out_frame[17] [0]), 
            .I3(n6_adj_4082), .O(n25952));
    defparam i4_4_lut_adj_1119.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1120 (.I0(\data_out_frame[5] [3]), .I1(n26015), 
            .I2(n1178), .I3(n28216), .O(n16_adj_4083));
    defparam i6_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1121 (.I0(n14978), .I1(n28457), .I2(n28548), 
            .I3(\data_out_frame[5] [7]), .O(n17_adj_4084));
    defparam i7_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1122 (.I0(n29994), .I1(n17_adj_4084), .I2(n15_adj_4085), 
            .I3(n16_adj_4083), .O(n4_adj_4037));
    defparam i1_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1123 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[12] [3]), 
            .I2(\data_out_frame[14] [4]), .I3(\data_out_frame[12] [1]), 
            .O(n28530));
    defparam i3_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1124 (.I0(n15279), .I1(n28530), .I2(\data_out_frame[14] [3]), 
            .I3(GND_net), .O(n28488));
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(n28120), .I1(n28488), .I2(GND_net), 
            .I3(GND_net), .O(n28379));
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15416));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1127 (.I0(\data_out_frame[7] [3]), .I1(n26337), 
            .I2(n28511), .I3(\data_out_frame[9] [6]), .O(n10_adj_4086));
    defparam i4_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28432));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1129 (.I0(n15416), .I1(n12_adj_3994), .I2(n28508), 
            .I3(n14612), .O(n26348));
    defparam i6_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_out_frame[19] [0]), .I1(n26348), 
            .I2(GND_net), .I3(GND_net), .O(n28405));
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1131 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[17] [2]), 
            .I2(n28162), .I3(\data_out_frame[17] [3]), .O(n28110));
    defparam i3_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(n28110), .I1(n28224), .I2(GND_net), 
            .I3(GND_net), .O(n28226));
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3393), 
            .CO(n23574));
    SB_LUT4 i1_2_lut_adj_1133 (.I0(\data_out_frame[23] [4]), .I1(n25952), 
            .I2(GND_net), .I3(GND_net), .O(n26444));
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n15767));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i39_4_lut (.I0(n69), .I1(n71), .I2(n70), .I3(n72), .O(n81_adj_4087));
    defparam i39_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1134 (.I0(\data_in_frame[19] [6]), .I1(n10_adj_4079), 
            .I2(\data_in_frame[19] [1]), .I3(\data_in_frame[19] [5]), .O(n12_adj_4088));
    defparam i5_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i41_4_lut (.I0(n81_adj_4087), .I1(n73), .I2(n80), .I3(n74), 
            .O(n29577));
    defparam i41_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1135 (.I0(n29577), .I1(n12_adj_4088), .I2(n28133), 
            .I3(\data_in_frame[19] [7]), .O(n29657));
    defparam i6_4_lut_adj_1135.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1136 (.I0(\data_in_frame[19] [0]), .I1(n29657), 
            .I2(GND_net), .I3(GND_net), .O(n28095));
    defparam i1_2_lut_adj_1136.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1137 (.I0(\data_in_frame[14] [4]), .I1(n25280), 
            .I2(\data_in_frame[12] [2]), .I3(GND_net), .O(n28189));
    defparam i2_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1138 (.I0(\data_in_frame[12] [3]), .I1(n28189), 
            .I2(n15111), .I3(GND_net), .O(n29658));
    defparam i2_3_lut_adj_1138.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1139 (.I0(\data_in_frame[2] [6]), .I1(n27981), 
            .I2(\data_in_frame[7] [4]), .I3(\data_in_frame[0] [4]), .O(n12_adj_4089));   // verilog/coms.v(76[16:27])
    defparam i5_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1140 (.I0(\data_in_frame[3] [0]), .I1(n12_adj_4089), 
            .I2(n28027), .I3(\data_in_frame[5] [2]), .O(n14648));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1141 (.I0(\data_in_frame[11] [6]), .I1(n14648), 
            .I2(\data_in_frame[9] [5]), .I3(n14756), .O(n28261));
    defparam i3_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\data_in_frame[13] [7]), .I1(n28201), 
            .I2(GND_net), .I3(GND_net), .O(n26318));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1143 (.I0(n28385), .I1(n15048), .I2(\data_in_frame[16] [0]), 
            .I3(\data_in_frame[14] [0]), .O(n14_adj_4090));
    defparam i6_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1144 (.I0(n28127), .I1(n14_adj_4090), .I2(n10_adj_4091), 
            .I3(n14459), .O(n28491));
    defparam i7_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14459));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1146 (.I0(n15021), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[11] [0]), .I3(n14459), .O(n28521));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1147 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[17] [5]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n28482));
    defparam i2_3_lut_adj_1147.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1148 (.I0(Kp_23__N_1201), .I1(n28250), .I2(n28345), 
            .I3(n6_adj_4092), .O(n28880));
    defparam i4_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28037));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1150 (.I0(\data_out_frame[19] [1]), .I1(n28379), 
            .I2(\data_out_frame[18] [6]), .I3(n6_adj_4093), .O(n26471));
    defparam i4_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28472));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28080));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1153 (.I0(\data_in_frame[4] [1]), .I1(n28285), 
            .I2(n28080), .I3(n15015), .O(Kp_23__N_973));   // verilog/coms.v(70[16:69])
    defparam i3_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1154 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[6] [2]), 
            .I2(n14908), .I3(n6_adj_4094), .O(n27918));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1155 (.I0(\data_in_frame[6] [3]), .I1(n28071), 
            .I2(n27918), .I3(Kp_23__N_973), .O(n15021));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1156 (.I0(n7_adj_4095), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n19871), .I3(GND_net), .O(n4040));
    defparam i2_3_lut_adj_1156.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(n29737), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26272));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28195));
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1159 (.I0(n26352), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[14] [4]), .I3(n30022), .O(n29382));
    defparam i3_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1160 (.I0(n14352), .I1(Kp_23__N_973), .I2(Kp_23__N_976), 
            .I3(\data_in_frame[8] [5]), .O(n14593));
    defparam i3_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28511));
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28318));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n14401));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1164 (.I0(n27991), .I1(n28318), .I2(n14632), 
            .I3(\data_in_frame[10] [6]), .O(n12_adj_4096));   // verilog/coms.v(76[16:43])
    defparam i5_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1165 (.I0(\data_in_frame[15] [1]), .I1(n12_adj_4096), 
            .I2(n28472), .I3(n15317), .O(n14505));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28250));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1167 (.I0(\data_in_frame[13] [5]), .I1(Kp_23__N_1446), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n14344));
    defparam i2_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1168 (.I0(\data_in_frame[13] [4]), .I1(n27963), 
            .I2(n14561), .I3(\data_in_frame[13] [3]), .O(n14_adj_4097));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\data_in_frame[15] [5]), .I1(n28114), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4098));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1170 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n27911));
    defparam i2_3_lut_adj_1170.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1171 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n29900));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1171.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1172 (.I0(n28020), .I1(n28288), .I2(\data_out_frame[9] [3]), 
            .I3(n27911), .O(n12_adj_4099));
    defparam i5_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1173 (.I0(\data_out_frame[9] [1]), .I1(n12_adj_4099), 
            .I2(n28533), .I3(n29900), .O(n28457));
    defparam i6_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1174 (.I0(n15395), .I1(n1174), .I2(n1260), .I3(n6_adj_4100), 
            .O(n14738));
    defparam i4_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1175 (.I0(n25261), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[9] [1]), .I3(GND_net), .O(n26359));
    defparam i2_3_lut_adj_1175.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1176 (.I0(\data_out_frame[6] [6]), .I1(n26359), 
            .I2(\data_out_frame[8] [7]), .I3(n13958), .O(n6_adj_4101));
    defparam i1_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1177 (.I0(n14738), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(n6_adj_4101), .O(n26375));
    defparam i4_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1178 (.I0(n9_adj_4098), .I1(n14_adj_4097), .I2(n26276), 
            .I3(n29862), .O(n26383));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1178.LUT_INIT = 16'h9669;
    SB_LUT4 equal_1188_i8_2_lut (.I0(Kp_23__N_1094), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4058));   // verilog/coms.v(236[9:81])
    defparam equal_1188_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1179 (.I0(n10_adj_4066), .I1(n15085), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n14645));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1179.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(Kp_23__N_1201), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n27963));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1181 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[13] [4]), .I3(GND_net), .O(n28385));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_17__7__I_0_3899_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1378));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_17__7__I_0_3899_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1182 (.I0(\data_in_frame[11] [4]), .I1(n27963), 
            .I2(n14645), .I3(GND_net), .O(Kp_23__N_1446));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1182.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1183 (.I0(n28457), .I1(\data_out_frame[7] [1]), 
            .I2(n25290), .I3(n28210), .O(n15_adj_4102));
    defparam i6_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1184 (.I0(n15_adj_4102), .I1(\data_out_frame[8] [0]), 
            .I2(n14_adj_4103), .I3(n15395), .O(n26015));
    defparam i8_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1185 (.I0(n28485), .I1(n28536), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n28003));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1185.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28288));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1187 (.I0(n8_adj_4065), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[12] [6]), .I3(GND_net), .O(n28441));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1188 (.I0(n28301), .I1(n27960), .I2(n14363), 
            .I3(n28402), .O(n10_adj_4104));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_in_frame[10] [5]), .I1(n14542), 
            .I2(GND_net), .I3(GND_net), .O(n28083));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27932));
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1191 (.I0(n14687), .I1(n28441), .I2(n27932), 
            .I3(n28083), .O(n12_adj_4105));
    defparam i5_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1192 (.I0(\data_in_frame[13] [0]), .I1(n12_adj_4105), 
            .I2(\data_in_frame[17] [4]), .I3(n28364), .O(n27974));
    defparam i6_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1193 (.I0(Kp_23__N_1443), .I1(Kp_23__N_1446), .I2(Kp_23__N_1378), 
            .I3(n28385), .O(n10_adj_4106));
    defparam i4_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1194 (.I0(n26383), .I1(n10_adj_4106), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n28493));
    defparam i5_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1195 (.I0(\data_in_frame[11] [4]), .I1(n14561), 
            .I2(\data_in_frame[11] [5]), .I3(GND_net), .O(n28221));
    defparam i2_3_lut_adj_1195.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1196 (.I0(n27984), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[5] [0]), .I3(\data_in_frame[7] [1]), .O(n14_adj_4107));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1197 (.I0(\data_in_frame[2] [6]), .I1(n14_adj_4107), 
            .I2(n10_adj_4108), .I3(\data_in_frame[4] [5]), .O(n10_adj_4066));   // verilog/coms.v(70[16:27])
    defparam i7_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1198 (.I0(n28356), .I1(\data_in_frame[4] [6]), 
            .I2(n15039), .I3(\data_in_frame[6] [6]), .O(n10_adj_4109));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1199 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[8] [7]), 
            .I2(n28068), .I3(\data_in_frame[8] [6]), .O(n15048));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n15766));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n15765));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1200 (.I0(\data_out_frame[23] [0]), .I1(n26457), 
            .I2(n26429), .I3(GND_net), .O(n28423));
    defparam i1_2_lut_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1201 (.I0(n28238), .I1(n28441), .I2(n14593), 
            .I3(n14693), .O(n12_adj_4110));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_in_frame[9] [0]), .I1(n15048), 
            .I2(GND_net), .I3(GND_net), .O(n27988));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1203 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[18] [0]), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n28373));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1204 (.I0(\data_in_frame[13] [6]), .I1(n28221), 
            .I2(n26397), .I3(\data_in_frame[16] [0]), .O(n29862));
    defparam i3_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1205 (.I0(Kp_23__N_1443), .I1(n28802), .I2(n13989), 
            .I3(n26296), .O(n7_adj_4111));
    defparam i2_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1206 (.I0(n7_adj_4111), .I1(\data_in_frame[13] [4]), 
            .I2(n29862), .I3(n28373), .O(n28133));
    defparam i4_4_lut_adj_1206.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1207 (.I0(\data_out_frame[23] [0]), .I1(n26457), 
            .I2(n26343), .I3(GND_net), .O(n28330));
    defparam i1_2_lut_3_lut_adj_1207.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1208 (.I0(n26471), .I1(n26270), .I2(n28518), 
            .I3(GND_net), .O(n6_adj_4024));
    defparam i1_2_lut_3_lut_adj_1208.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1209 (.I0(\data_in_frame[13] [1]), .I1(n12_adj_4110), 
            .I2(n28514), .I3(\data_in_frame[12] [7]), .O(n14942));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1210 (.I0(n26471), .I1(n26270), .I2(n26335), 
            .I3(n28420), .O(n25305));
    defparam i2_3_lut_4_lut_adj_1210.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1211 (.I0(n14819), .I1(n28124), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n15114));
    defparam i2_3_lut_adj_1211.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1212 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n28429));
    defparam i2_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1213 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[12] [0]), .I3(GND_net), .O(n28235));
    defparam i2_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(n15026), .I1(n14548), .I2(GND_net), 
            .I3(GND_net), .O(n27984));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1215 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27960));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1215.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(n15034), .I1(n28057), .I2(GND_net), 
            .I3(GND_net), .O(n28469));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1217 (.I0(n15247), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n8_adj_4112));
    defparam i3_3_lut_adj_1217.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28089));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1219 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(n28141), .I3(Kp_23__N_868), .O(n28496));
    defparam i3_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1220 (.I0(n27946), .I1(\data_in_frame[2] [1]), 
            .I2(n8_adj_4112), .I3(\data_in_frame[0] [6]), .O(n22_adj_4113));
    defparam i7_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i15147_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n19686));
    defparam i15147_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1221 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n19686), .I3(byte_transmit_counter[2]), .O(n19835));
    defparam i2_4_lut_adj_1221.LUT_INIT = 16'h8880;
    SB_LUT4 i2_3_lut_adj_1222 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n6_adj_3992));
    defparam i2_3_lut_adj_1222.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1223 (.I0(n27747), .I1(n27894), .I2(n27859), 
            .I3(n6_adj_4075), .O(n19871));
    defparam i4_4_lut_adj_1223.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_782_i1_4_lut (.I0(n7_adj_4114), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n4626), .I3(n8_adj_4115), .O(n3505[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_782_i1_4_lut.LUT_INIT = 16'h0c5c;
    SB_LUT4 i2_3_lut_4_lut_adj_1224 (.I0(n14304), .I1(n14338), .I2(n31_adj_4068), 
            .I3(n27757), .O(n4725));   // verilog/coms.v(263[5:27])
    defparam i2_3_lut_4_lut_adj_1224.LUT_INIT = 16'h0100;
    SB_LUT4 i2_3_lut_4_lut_adj_1225 (.I0(n14304), .I1(n14338), .I2(n31_adj_4068), 
            .I3(n12002), .O(n29573));   // verilog/coms.v(263[5:27])
    defparam i2_3_lut_4_lut_adj_1225.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1226 (.I0(n28233), .I1(n14060), .I2(n28259), 
            .I3(n28444), .O(n28518));
    defparam i2_3_lut_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i11652_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n16191));
    defparam i11652_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11653_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n16192));
    defparam i11653_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11654_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n16193));
    defparam i11654_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11655_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n16194));
    defparam i11655_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1227 (.I0(\data_out_frame[25] [1]), .I1(n26288), 
            .I2(\data_out_frame[25] [2]), .I3(n14060), .O(n29733));
    defparam i2_3_lut_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i11656_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n16195));
    defparam i11656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1228 (.I0(\data_out_frame[25] [1]), .I1(n26288), 
            .I2(n28207), .I3(GND_net), .O(n28209));
    defparam i1_2_lut_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(n771), .I1(n9411), .I2(n14295), 
            .I3(GND_net), .O(n4_adj_3990));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'h0404;
    SB_LUT4 i11657_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n16196));
    defparam i11657_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[6] [6]), .I3(n10_adj_4081), .O(n29704));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1230 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n28307));
    defparam i1_2_lut_3_lut_adj_1230.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1231 (.I0(n28496), .I1(n28080), .I2(n28351), 
            .I3(\data_in_frame[5] [6]), .O(n25_adj_4117));
    defparam i10_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(n28298), .I1(n14357), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4118));
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1233 (.I0(\data_in_frame[1] [3]), .I1(n27935), 
            .I2(n28454), .I3(\data_in_frame[5] [3]), .O(n24_adj_4119));
    defparam i9_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i11658_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n16197));
    defparam i11658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11659_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27867), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n16198));
    defparam i11659_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1234 (.I0(n25_adj_4117), .I1(n14908), .I2(n22_adj_4113), 
            .I3(n28469), .O(n28_adj_4120));
    defparam i13_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1235 (.I0(n14363), .I1(n28_adj_4120), .I2(n24_adj_4119), 
            .I3(n16_adj_4118), .O(n25278));
    defparam i14_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_in_frame[5] [1]), .I1(n28049), 
            .I2(GND_net), .I3(GND_net), .O(n28351));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1237 (.I0(\data_in_frame[7] [2]), .I1(n28390), 
            .I2(n28351), .I3(n14548), .O(n15085));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(n15085), .I1(n14756), .I2(GND_net), 
            .I3(GND_net), .O(n26320));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 i4_2_lut_adj_1239 (.I0(n14917), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4121));
    defparam i4_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1240 (.I0(n26320), .I1(n28411), .I2(n14493), 
            .I3(n15034), .O(n24_adj_4122));
    defparam i10_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1241 (.I0(\data_in_frame[14] [1]), .I1(n26279), 
            .I2(\data_in_frame[13] [7]), .I3(n25278), .O(n22_adj_4123));
    defparam i8_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1242 (.I0(\data_in_frame[2] [2]), .I1(n24_adj_4122), 
            .I2(n18_adj_4121), .I3(\data_in_frame[0] [1]), .O(n26_adj_4124));
    defparam i12_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1243 (.I0(n28235), .I1(n26_adj_4124), .I2(n22_adj_4123), 
            .I3(\data_in_frame[9] [2]), .O(n28265));
    defparam i13_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1244 (.I0(\data_in_frame[16] [4]), .I1(n28265), 
            .I2(\data_in_frame[16] [3]), .I3(n29131), .O(n28802));
    defparam i3_4_lut_adj_1244.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27921));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28402));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\data_in_frame[5] [6]), .I1(n14705), 
            .I2(GND_net), .I3(GND_net), .O(n28145));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n27935));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1249 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n14304), .I3(GND_net), .O(n63_adj_3));   // verilog/coms.v(201[5:24])
    defparam i2_3_lut_adj_1249.LUT_INIT = 16'hfbfb;
    SB_LUT4 equal_103_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4116));   // verilog/coms.v(154[7:23])
    defparam equal_103_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_3_lut_adj_1250 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n28324));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1250.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_944));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4126));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1252 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[10] [2]), 
            .I2(\data_in_frame[7] [7]), .I3(n6_adj_4126), .O(n27915));
    defparam i4_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1253 (.I0(\data_in_frame[5] [4]), .I1(n15336), 
            .I2(n12761), .I3(\data_in_frame[3] [5]), .O(n28298));
    defparam i3_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1254 (.I0(n14368), .I1(n28061), .I2(n14917), 
            .I3(GND_net), .O(n14617));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1254.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1255 (.I0(n14617), .I1(n28298), .I2(n27915), 
            .I3(Kp_23__N_944), .O(n15111));
    defparam i3_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1256 (.I0(\data_in_frame[12] [5]), .I1(n15111), 
            .I2(\data_in_frame[14] [6]), .I3(\data_in_frame[12] [4]), .O(n27991));
    defparam i3_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1257 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(\data_in_frame[10] [4]), .I3(\data_in_frame[5] [7]), .O(n16_adj_4127));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1258 (.I0(n28145), .I1(n28402), .I2(\data_in_frame[2] [0]), 
            .I3(n27921), .O(n17_adj_4128));   // verilog/coms.v(78[16:27])
    defparam i7_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1259 (.I0(n17_adj_4128), .I1(\data_in_frame[6] [0]), 
            .I2(n16_adj_4127), .I3(\data_in_frame[6] [2]), .O(n14687));   // verilog/coms.v(78[16:27])
    defparam i9_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(n14687), .I1(n27991), .I2(GND_net), 
            .I3(GND_net), .O(n15120));
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28336));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27946));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1263 (.I0(n3_adj_4129), .I1(n28361), .I2(n28071), 
            .I3(\data_in_frame[2] [0]), .O(Kp_23__N_976));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_976), 
            .I2(GND_net), .I3(GND_net), .O(n28011));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1265 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n15026));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28285));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28454));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1268 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n14548));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1269 (.I0(\data_in_frame[1] [7]), .I1(n28454), 
            .I2(n28285), .I3(n15026), .O(Kp_23__N_979));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\data_in_frame[4] [4]), .I1(n14548), 
            .I2(GND_net), .I3(GND_net), .O(n15039));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h6666;
    SB_LUT4 equal_104_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4130));   // verilog/coms.v(154[7:23])
    defparam equal_104_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i11075_2_lut (.I0(n15481), .I1(n14327), .I2(GND_net), .I3(GND_net), 
            .O(n15614));   // verilog/coms.v(127[12] 300[6])
    defparam i11075_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11644_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n16183));
    defparam i11644_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11645_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n16184));
    defparam i11645_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28159));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1272 (.I0(n15039), .I1(\data_in_frame[4] [5]), 
            .I2(Kp_23__N_979), .I3(n6_adj_4131), .O(Kp_23__N_1094));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(\data_in_frame[7] [7]), .I1(n12761), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n14917));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28356));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14363));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28361));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1277 (.I0(n15096), .I1(Kp_23__N_1186), .I2(\data_in_frame[10] [0]), 
            .I3(GND_net), .O(n25280));
    defparam i2_3_lut_adj_1277.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14352));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1279 (.I0(n28068), .I1(n28527), .I2(\data_in_frame[6] [3]), 
            .I3(n28396), .O(n20_adj_4132));
    defparam i8_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1280 (.I0(n28361), .I1(n14363), .I2(\data_in_frame[9] [6]), 
            .I3(n28463), .O(n19_adj_4133));
    defparam i7_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1281 (.I0(n28356), .I1(n14917), .I2(n27925), 
            .I3(n14638), .O(n21_adj_4134));
    defparam i9_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1282 (.I0(n21_adj_4134), .I1(n19_adj_4133), .I2(n20_adj_4132), 
            .I3(GND_net), .O(n26279));
    defparam i11_3_lut_adj_1282.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28141));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27981));
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14378));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1286 (.I0(\data_in_frame[7] [3]), .I1(n28390), 
            .I2(n28496), .I3(\data_in_frame[5] [1]), .O(n14756));
    defparam i1_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1287 (.I0(n28124), .I1(Kp_23__N_1186), .I2(\data_in_frame[12] [2]), 
            .I3(n28382), .O(n10_adj_4135));
    defparam i4_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_in_frame[5] [5]), .I1(n15336), 
            .I2(GND_net), .I3(GND_net), .O(n14521));
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4136));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1290 (.I0(Kp_23__N_868), .I1(\data_in_frame[3] [0]), 
            .I2(n14378), .I3(n6_adj_4136), .O(n28049));
    defparam i4_4_lut_adj_1290.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14536));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1292 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n14705));
    defparam i2_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_in_frame[4] [5]), .I1(n25278), 
            .I2(GND_net), .I3(GND_net), .O(n28230));
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1294 (.I0(n14705), .I1(n14536), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[3] [3]), .O(n12761));
    defparam i3_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 i11646_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n16185));
    defparam i11646_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1295 (.I0(n29381), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28017));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1295.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1296 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n28057));
    defparam i2_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1297 (.I0(\data_in_frame[7] [4]), .I1(n26346), 
            .I2(n14819), .I3(\data_in_frame[9] [6]), .O(n28_adj_3984));   // verilog/coms.v(85[17:70])
    defparam i12_4_lut_adj_1297.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1298 (.I0(n28049), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[12] [1]), .I3(n28393), .O(n26_adj_3983));   // verilog/coms.v(85[17:70])
    defparam i10_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1299 (.I0(\data_in_frame[11] [7]), .I1(n10_adj_4135), 
            .I2(n26346), .I3(n14638), .O(n29131));
    defparam i5_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n32227));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n32227_bdd_4_lut (.I0(n32227), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n32230));
    defparam n32227_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1300 (.I0(n28399), .I1(\data_in_frame[8] [2]), 
            .I2(\data_in_frame[10] [3]), .I3(\data_in_frame[8] [1]), .O(n6_adj_4137));   // verilog/coms.v(75[16:27])
    defparam i1_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n31966), .I2(n31095), .I3(byte_transmit_counter[4]), .O(n32221));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n32221_bdd_4_lut (.I0(n32221), .I1(n14_adj_3982), .I2(n7_adj_3981), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n32221_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1301 (.I0(n14917), .I1(\data_in_frame[3] [7]), 
            .I2(n28460), .I3(n6_adj_4137), .O(n14693));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1302 (.I0(\data_in_frame[18] [7]), .I1(n29131), 
            .I2(\data_in_frame[16] [5]), .I3(GND_net), .O(n28185));
    defparam i2_3_lut_adj_1302.LUT_INIT = 16'h6969;
    SB_LUT4 i11647_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n16186));
    defparam i11647_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1303 (.I0(n28472), .I1(n28514), .I2(\data_in_frame[17] [1]), 
            .I3(GND_net), .O(n28545));
    defparam i2_3_lut_adj_1303.LUT_INIT = 16'h9696;
    SB_LUT4 i11648_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n16187));
    defparam i11648_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11649_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n16188));
    defparam i11649_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11650_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n16189));
    defparam i11650_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1304 (.I0(n28221), .I1(n28261), .I2(n14344), 
            .I3(n28201), .O(n12_adj_4138));
    defparam i5_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_26341 (.I0(byte_transmit_counter[3]), 
            .I1(n31585), .I2(n31089), .I3(byte_transmit_counter[4]), .O(n32215));
    defparam byte_transmit_counter_3__bdd_4_lut_26341.LUT_INIT = 16'he4aa;
    SB_LUT4 n32215_bdd_4_lut (.I0(n32215), .I1(n14_adj_3978), .I2(n7_adj_3977), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n32215_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1305 (.I0(\data_in_frame[16] [1]), .I1(n12_adj_4138), 
            .I2(n28265), .I3(\data_in_frame[16] [2]), .O(n26296));
    defparam i6_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26346 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n32209));
    defparam byte_transmit_counter_0__bdd_4_lut_26346.LUT_INIT = 16'he4aa;
    SB_LUT4 n32209_bdd_4_lut (.I0(n32209), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n32212));
    defparam n32209_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(n14561), .I1(n27957), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4139));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26331 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n32203));
    defparam byte_transmit_counter_0__bdd_4_lut_26331.LUT_INIT = 16'he4aa;
    SB_LUT4 n32203_bdd_4_lut (.I0(n32203), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n32206));
    defparam n32203_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1307 (.I0(\data_in_frame[14] [0]), .I1(n26318), 
            .I2(n14645), .I3(n6_adj_4139), .O(n13989));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_1307.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26326 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n32197));
    defparam byte_transmit_counter_0__bdd_4_lut_26326.LUT_INIT = 16'he4aa;
    SB_LUT4 n32197_bdd_4_lut (.I0(n32197), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n32200));
    defparam n32197_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_rep_17_2_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32610));   // verilog/coms.v(78[16:27])
    defparam i1_rep_17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26321 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n32191));
    defparam byte_transmit_counter_0__bdd_4_lut_26321.LUT_INIT = 16'he4aa;
    SB_LUT4 n32191_bdd_4_lut (.I0(n32191), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n32194));
    defparam n32191_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_rep_19_2_lut (.I0(n13989), .I1(n26296), .I2(GND_net), .I3(GND_net), 
            .O(n32612));
    defparam i1_rep_19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26316 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n32185));
    defparam byte_transmit_counter_0__bdd_4_lut_26316.LUT_INIT = 16'he4aa;
    SB_LUT4 n32185_bdd_4_lut (.I0(n32185), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n32188));
    defparam n32185_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1308 (.I0(n28505), .I1(n28310), .I2(\data_in_frame[21] [3]), 
            .I3(n28545), .O(n10_adj_4140));
    defparam i4_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26311 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n32179));
    defparam byte_transmit_counter_0__bdd_4_lut_26311.LUT_INIT = 16'he4aa;
    SB_LUT4 n32179_bdd_4_lut (.I0(n32179), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n32182));
    defparam n32179_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_rep_20_2_lut (.I0(n28429), .I1(n28545), .I2(GND_net), .I3(GND_net), 
            .O(n32613));   // verilog/coms.v(76[16:43])
    defparam i1_rep_20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1309 (.I0(n15114), .I1(n32613), .I2(\data_in_frame[19] [4]), 
            .I3(n14942), .O(n12_adj_4141));   // verilog/coms.v(76[16:43])
    defparam i5_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i111_2_lut_3_lut (.I0(n771), .I1(n9411), .I2(n14309), .I3(GND_net), 
            .O(n41_adj_3988));   // verilog/coms.v(157[6] 159[9])
    defparam i111_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2_3_lut_4_lut_adj_1310 (.I0(n26326), .I1(\data_out_frame[17] [0]), 
            .I2(n30149), .I3(\data_out_frame[17] [1]), .O(n28903));
    defparam i2_3_lut_4_lut_adj_1310.LUT_INIT = 16'h9669;
    SB_LUT4 i11651_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27867), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n16190));
    defparam i11651_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11636_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n16175));
    defparam i11636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1311 (.I0(n32_adj_4143), .I1(n1_adj_3989), 
            .I2(\FRAME_MATCHER.state[1] ), .I3(GND_net), .O(n123));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_3_lut_adj_1311.LUT_INIT = 16'h8080;
    SB_LUT4 i11637_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n16176));
    defparam i11637_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1312 (.I0(n32_adj_4143), .I1(n1_adj_3989), 
            .I2(n63), .I3(GND_net), .O(n9411));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_3_lut_adj_1312.LUT_INIT = 16'h8080;
    SB_LUT4 i11638_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n16177));
    defparam i11638_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1313 (.I0(\data_in[2] [5]), .I1(\data_in[2] [6]), 
            .I2(n33), .I3(GND_net), .O(n14313));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1313.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_rep_16_2_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32609));   // verilog/coms.v(72[16:41])
    defparam i1_rep_16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26306 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n32161));
    defparam byte_transmit_counter_0__bdd_4_lut_26306.LUT_INIT = 16'he4aa;
    SB_LUT4 n32161_bdd_4_lut (.I0(n32161), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n32164));
    defparam n32161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1314 (.I0(\data_in_frame[21] [2]), .I1(n32609), 
            .I2(\data_in_frame[16] [7]), .I3(n14967), .O(n12_adj_4144));   // verilog/coms.v(72[16:41])
    defparam i5_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_26336 (.I0(byte_transmit_counter[3]), 
            .I1(n31972), .I2(n31150), .I3(byte_transmit_counter[4]), .O(n32155));
    defparam byte_transmit_counter_3__bdd_4_lut_26336.LUT_INIT = 16'he4aa;
    SB_LUT4 n32155_bdd_4_lut (.I0(n32155), .I1(n14_adj_3974), .I2(n7_adj_3973), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n32155_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1315 (.I0(\data_in_frame[19] [6]), .I1(n28880), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n6_adj_4145));
    defparam i2_3_lut_adj_1315.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_26286 (.I0(byte_transmit_counter[3]), 
            .I1(n31978), .I2(n31112), .I3(byte_transmit_counter[4]), .O(n32149));
    defparam byte_transmit_counter_3__bdd_4_lut_26286.LUT_INIT = 16'he4aa;
    SB_LUT4 n32149_bdd_4_lut (.I0(n32149), .I1(n14_adj_3970), .I2(n7_adj_3969), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n32149_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1316 (.I0(\data_in_frame[19] [0]), .I1(n12_adj_4144), 
            .I2(n28336), .I3(n15120), .O(n29711));   // verilog/coms.v(72[16:41])
    defparam i6_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_26281 (.I0(byte_transmit_counter[3]), 
            .I1(n31984), .I2(n31108), .I3(byte_transmit_counter[4]), .O(n32143));
    defparam byte_transmit_counter_3__bdd_4_lut_26281.LUT_INIT = 16'he4aa;
    SB_LUT4 n32143_bdd_4_lut (.I0(n32143), .I1(n14_adj_3967), .I2(n7_adj_3966), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n32143_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_rep_5_3_lut (.I0(n28802), .I1(n13989), .I2(n26296), .I3(GND_net), 
            .O(n32598));
    defparam i1_rep_5_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_26276 (.I0(byte_transmit_counter[3]), 
            .I1(n31990), .I2(n31105), .I3(byte_transmit_counter[4]), .O(n32137));
    defparam byte_transmit_counter_3__bdd_4_lut_26276.LUT_INIT = 16'he4aa;
    SB_LUT4 n32137_bdd_4_lut (.I0(n32137), .I1(n14_adj_3964), .I2(n7_adj_3963), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n32137_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_1317 (.I0(n28133), .I1(\data_in_frame[20] [0]), 
            .I2(\data_in_frame[19] [7]), .I3(GND_net), .O(n14_adj_4146));
    defparam i5_3_lut_adj_1317.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_26271 (.I0(byte_transmit_counter[3]), 
            .I1(n31996), .I2(n31102), .I3(byte_transmit_counter[4]), .O(n32131));
    defparam byte_transmit_counter_3__bdd_4_lut_26271.LUT_INIT = 16'he4aa;
    SB_LUT4 n32131_bdd_4_lut (.I0(n32131), .I1(n14_adj_3961), .I2(n7_adj_3960), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n32131_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1318 (.I0(n32598), .I1(n28493), .I2(\data_in_frame[19] [6]), 
            .I3(n27974), .O(n15_adj_4147));
    defparam i6_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_26266 (.I0(byte_transmit_counter[3]), 
            .I1(n32104), .I2(n31099), .I3(byte_transmit_counter[4]), .O(n32125));
    defparam byte_transmit_counter_3__bdd_4_lut_26266.LUT_INIT = 16'he4aa;
    SB_LUT4 n32125_bdd_4_lut (.I0(n32125), .I1(n14), .I2(n7), .I3(byte_transmit_counter[4]), 
            .O(tx_data[3]));
    defparam n32125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1319 (.I0(n28429), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[21] [1]), .I3(n28505), .O(n10_adj_4148));
    defparam i4_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1320 (.I0(n15_adj_4147), .I1(\data_in_frame[17] [5]), 
            .I2(n14_adj_4146), .I3(n28880), .O(n30020));
    defparam i8_4_lut_adj_1320.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26291 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n32113));
    defparam byte_transmit_counter_0__bdd_4_lut_26291.LUT_INIT = 16'he4aa;
    SB_LUT4 n32113_bdd_4_lut (.I0(n32113), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n32116));
    defparam n32113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1321 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[21] [4]), 
            .I2(\data_in_frame[16] [6]), .I3(GND_net), .O(n9_adj_4149));
    defparam i2_3_lut_adj_1321.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1322 (.I0(n14505), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[17] [0]), .I3(\data_in_frame[19] [2]), .O(n11));
    defparam i4_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n31100), .I2(n31101), .I3(byte_transmit_counter[2]), .O(n32101));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n32101_bdd_4_lut (.I0(n32101), .I1(n17_adj_3956), .I2(n16_adj_3955), 
            .I3(byte_transmit_counter[2]), .O(n32104));
    defparam n32101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1323 (.I0(n26276), .I1(n27932), .I2(\data_in_frame[13] [2]), 
            .I3(n15317), .O(n29270));
    defparam i3_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1324 (.I0(n29270), .I1(\data_in_frame[19] [4]), 
            .I2(\data_in_frame[21] [6]), .I3(\data_in_frame[15] [3]), .O(n12_adj_4150));
    defparam i5_4_lut_adj_1324.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26252 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n32089));
    defparam byte_transmit_counter_0__bdd_4_lut_26252.LUT_INIT = 16'he4aa;
    SB_LUT4 n32089_bdd_4_lut (.I0(n32089), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n32092));
    defparam n32089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1325 (.I0(\data_in_frame[20] [6]), .I1(n32610), 
            .I2(n28802), .I3(n13989), .O(n29351));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1325.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26233 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n32083));
    defparam byte_transmit_counter_0__bdd_4_lut_26233.LUT_INIT = 16'he4aa;
    SB_LUT4 n32083_bdd_4_lut (.I0(n32083), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n32086));
    defparam n32083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1326 (.I0(n14505), .I1(n12_adj_4150), .I2(n27974), 
            .I3(\data_in_frame[19] [5]), .O(n29325));
    defparam i6_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26228 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n32077));
    defparam byte_transmit_counter_0__bdd_4_lut_26228.LUT_INIT = 16'he4aa;
    SB_LUT4 n32077_bdd_4_lut (.I0(n32077), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n32080));
    defparam n32077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1327 (.I0(\data_in_frame[20] [3]), .I1(n28491), 
            .I2(n26383), .I3(\data_in_frame[18] [1]), .O(n29156));
    defparam i3_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26223 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n32071));
    defparam byte_transmit_counter_0__bdd_4_lut_26223.LUT_INIT = 16'he4aa;
    SB_LUT4 n32071_bdd_4_lut (.I0(n32071), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n32074));
    defparam n32071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1328 (.I0(n11), .I1(n9_adj_4149), .I2(n29658), 
            .I3(n15120), .O(n29303));
    defparam i6_4_lut_adj_1328.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26218 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n32065));
    defparam byte_transmit_counter_0__bdd_4_lut_26218.LUT_INIT = 16'he4aa;
    SB_LUT4 n32065_bdd_4_lut (.I0(n32065), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n32068));
    defparam n32065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11639_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n16178));
    defparam i11639_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state[1] ), .I3(n1_adj_4151), .O(n5_adj_3985));   // verilog/coms.v(145[4] 299[11])
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'h6745;
    SB_LUT4 i11640_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n16179));
    defparam i11640_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n11873), .I1(n14327), .I2(n87), 
            .I3(\FRAME_MATCHER.state [12]), .O(n88));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i6_4_lut_adj_1329 (.I0(n27929), .I1(\data_in_frame[19] [7]), 
            .I2(n28448), .I3(n28114), .O(n16_adj_4152));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26213 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n32059));
    defparam byte_transmit_counter_0__bdd_4_lut_26213.LUT_INIT = 16'he4aa;
    SB_LUT4 n32059_bdd_4_lut (.I0(n32059), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n32062));
    defparam n32059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1330 (.I0(\data_in_frame[9] [1]), .I1(n28373), 
            .I2(n28521), .I3(n27988), .O(n17_adj_4153));   // verilog/coms.v(85[17:70])
    defparam i7_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26208 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n32053));
    defparam byte_transmit_counter_0__bdd_4_lut_26208.LUT_INIT = 16'he4aa;
    SB_LUT4 n32053_bdd_4_lut (.I0(n32053), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n32056));
    defparam n32053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1331 (.I0(\data_in_frame[18] [4]), .I1(n32612), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[18] [3]), .O(n29740));
    defparam i3_4_lut_adj_1331.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26203 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n32047));
    defparam byte_transmit_counter_0__bdd_4_lut_26203.LUT_INIT = 16'he4aa;
    SB_LUT4 n32047_bdd_4_lut (.I0(n32047), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n32050));
    defparam n32047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26198 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n32041));
    defparam byte_transmit_counter_0__bdd_4_lut_26198.LUT_INIT = 16'he4aa;
    SB_LUT4 n32041_bdd_4_lut (.I0(n32041), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n32044));
    defparam n32041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1332 (.I0(\data_in_frame[19] [3]), .I1(n12_adj_4141), 
            .I2(n28310), .I3(\data_in_frame[21] [5]), .O(n29675));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1333 (.I0(\data_in_frame[18] [3]), .I1(n28491), 
            .I2(\data_in_frame[20] [4]), .I3(n26296), .O(n28896));
    defparam i3_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26193 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n32029));
    defparam byte_transmit_counter_0__bdd_4_lut_26193.LUT_INIT = 16'he4aa;
    SB_LUT4 n32029_bdd_4_lut (.I0(n32029), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n32032));
    defparam n32029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1334 (.I0(\data_in_frame[20] [7]), .I1(n28095), 
            .I2(n28802), .I3(\data_in_frame[18] [5]), .O(n29177));
    defparam i3_4_lut_adj_1334.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26184 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n32023));
    defparam byte_transmit_counter_0__bdd_4_lut_26184.LUT_INIT = 16'he4aa;
    SB_LUT4 n32023_bdd_4_lut (.I0(n32023), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n32026));
    defparam n32023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1335 (.I0(n29711), .I1(n14942), .I2(n6_adj_4145), 
            .I3(\data_in_frame[21] [7]), .O(n22_adj_4154));
    defparam i6_4_lut_adj_1335.LUT_INIT = 16'hd77d;
    SB_LUT4 i12_4_lut_adj_1336 (.I0(n28896), .I1(n29675), .I2(n29624), 
            .I3(n29740), .O(n28_adj_4155));
    defparam i12_4_lut_adj_1336.LUT_INIT = 16'hfeff;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26179 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n32011));
    defparam byte_transmit_counter_0__bdd_4_lut_26179.LUT_INIT = 16'he4aa;
    SB_LUT4 n32011_bdd_4_lut (.I0(n32011), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n32014));
    defparam n32011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1337 (.I0(n17_adj_4153), .I1(n15317), .I2(n16_adj_4152), 
            .I3(\data_in_frame[20] [1]), .O(n29199));   // verilog/coms.v(85[17:70])
    defparam i9_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i14599_2_lut_3_lut_4_lut (.I0(n11873), .I1(n14327), .I2(n87), 
            .I3(\FRAME_MATCHER.state [13]), .O(n19123));
    defparam i14599_2_lut_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1338 (.I0(n14164), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n11605), .O(n7_adj_3991));
    defparam i1_2_lut_3_lut_4_lut_adj_1338.LUT_INIT = 16'h1000;
    SB_LUT4 i11641_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n16180));
    defparam i11641_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11642_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n16181));
    defparam i11642_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14600_2_lut_3_lut_4_lut (.I0(n11873), .I1(n14327), .I2(n87), 
            .I3(\FRAME_MATCHER.state [14]), .O(n19125));
    defparam i14600_2_lut_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i11643_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27867), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n16182));
    defparam i11643_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14601_2_lut_3_lut_4_lut (.I0(n11873), .I1(n14327), .I2(n87), 
            .I3(\FRAME_MATCHER.state [17]), .O(n19127));
    defparam i14601_2_lut_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i14630_2_lut_3_lut_4_lut (.I0(n11873), .I1(n14327), .I2(n87), 
            .I3(\FRAME_MATCHER.state [30]), .O(n19157));
    defparam i14630_2_lut_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i15331_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n19871), .O(n4626));
    defparam i15331_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1339 (.I0(n26326), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[19] [0]), .I3(n26348), .O(n6_adj_4093));
    defparam i1_2_lut_3_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1340 (.I0(n11873), .I1(n14327), .I2(n87), 
            .I3(\FRAME_MATCHER.state [31]), .O(n7_adj_4156));
    defparam i1_2_lut_3_lut_4_lut_adj_1340.LUT_INIT = 16'hf200;
    SB_LUT4 i15108_1_lut_3_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), 
            .I1(\FRAME_MATCHER.state[0] ), .I2(n14316), .I3(n14295), .O(n2028));
    defparam i15108_1_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h04cc;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in[2] [5]), .I1(\data_in[2] [6]), 
            .I2(n33), .I3(n18546), .O(n32_adj_4143));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 equal_97_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4142));   // verilog/coms.v(154[7:23])
    defparam equal_97_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1341 (.I0(\data_in_frame[9] [4]), .I1(n15085), 
            .I2(n14756), .I3(n28261), .O(n28262));
    defparam i1_2_lut_3_lut_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1342 (.I0(n14588), .I1(Kp_23__N_1094), 
            .I2(\data_in_frame[8] [7]), .I3(\data_in_frame[18] [2]), .O(n28127));
    defparam i1_2_lut_3_lut_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1343 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[1] [5]), .O(n28301));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1344 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[16] [6]), 
            .I2(n10_adj_4140), .I3(\data_in_frame[19] [2]), .O(n29624));
    defparam i5_3_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 equal_106_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4157));   // verilog/coms.v(154[7:23])
    defparam equal_106_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_4_lut_adj_1345 (.I0(\data_in_frame[18] [7]), .I1(n29131), 
            .I2(\data_in_frame[16] [5]), .I3(n14693), .O(n28505));
    defparam i1_2_lut_4_lut_adj_1345.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1346 (.I0(\data_in_frame[16] [7]), .I1(n15021), 
            .I2(\data_in_frame[10] [5]), .I3(n14542), .O(n28310));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3950), .S(n3_adj_3954));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3942), .S(n3_adj_3953));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1347 (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[5] [5]), 
            .I2(n15336), .I3(n14845), .O(n28393));
    defparam i2_3_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1348 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [2]), .O(n15336));
    defparam i1_2_lut_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1349 (.I0(\data_in_frame[4] [5]), .I1(n25278), 
            .I2(n14493), .I3(n15026), .O(n28396));
    defparam i2_3_lut_4_lut_adj_1349.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1350 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[0] [1]), .I3(n28159), .O(n6_adj_4131));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n3_adj_4129));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n14368));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(n4452), .I1(n9411), .I2(n14295), 
            .I3(GND_net), .O(n3_adj_3993));   // verilog/coms.v(259[6] 261[9])
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(n14316), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n14327));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'hbfbf;
    SB_LUT4 i3_3_lut_adj_1355 (.I0(\data_in_frame[18] [6]), .I1(n29658), 
            .I2(n28095), .I3(GND_net), .O(n8_adj_4158));
    defparam i3_3_lut_adj_1355.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[6] [7]), .I3(GND_net), .O(n28411));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1357 (.I0(n28233), .I1(n14060), .I2(\data_out_frame[25] [3]), 
            .I3(\data_out_frame[25] [2]), .O(n27906));
    defparam i1_2_lut_3_lut_4_lut_adj_1357.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n6_adj_3992), .O(n8_adj_4115));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i11628_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n16167));
    defparam i11628_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11629_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n16168));
    defparam i11629_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1358 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3] [6]), .I3(GND_net), .O(n14908));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1358.LUT_INIT = 16'h9696;
    SB_LUT4 i11630_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n16169));
    defparam i11630_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(\data_in_frame[5] [5]), .I1(n15026), 
            .I2(n14548), .I3(GND_net), .O(n14357));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1360 (.I0(n14561), .I1(\data_in_frame[9] [0]), 
            .I2(n15048), .I3(\data_in_frame[11] [3]), .O(Kp_23__N_1443));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i11631_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n16170));
    defparam i11631_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1361 (.I0(\data_in_frame[6] [7]), .I1(n10_adj_4109), 
            .I2(n15034), .I3(n28057), .O(n14588));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i11632_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n16171));
    defparam i11632_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_in_frame[9] [4]), .I1(n15085), 
            .I2(n14756), .I3(GND_net), .O(n26397));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1363 (.I0(\data_in_frame[20] [2]), .I1(n14588), 
            .I2(n28493), .I3(n6_adj_4159), .O(n29496));
    defparam i4_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[15] [2]), .I3(\data_in_frame[15] [1]), .O(n28238));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i11633_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n16172));
    defparam i11633_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1365 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n14_adj_4103));
    defparam i5_3_lut_4_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i11634_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n16173));
    defparam i11634_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1366 (.I0(n14588), .I1(Kp_23__N_1094), .I2(\data_in_frame[8] [7]), 
            .I3(GND_net), .O(Kp_23__N_1201));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3936), .S(n3_adj_3952));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3934), .S(n3_adj_3951));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3933), .S(n3_adj_3949));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3931), .S(n3_adj_3948));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3928), .S(n3_adj_3947));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3923), .S(n3_adj_3946));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3922), .S(n3_adj_3945));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3919), .S(n3_adj_3944));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3916), .S(n3_adj_3943));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3914), .S(n3_adj_3941));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3913), .S(n3_adj_3940));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3912), .S(n3_adj_3939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3910), .S(n3_adj_3938));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3908), .S(n3_adj_3937));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3907), .S(n3_adj_3935));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3906), .S(n3_adj_3932));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3905), .S(n3_adj_3930));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3904), .S(n3_adj_3929));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3903), .S(n3_adj_3927));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3902), .S(n3_adj_3926));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3901), .S(n3_adj_3925));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3900), .S(n3_adj_3924));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3899), .S(n3_adj_3921));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3898), .S(n3_adj_3920));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3897), .S(n3_adj_3918));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3896), .S(n3_adj_3917));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3895), .S(n3_adj_3915));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3894), .S(n3_adj_3911));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3893), .S(n3_adj_3909));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n15514), .D(n29910));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1367 (.I0(n15015), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [4]), .I3(n28463), .O(n14819));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i11635_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27867), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n16174));
    defparam i11635_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[11] [4]), .I3(GND_net), .O(n6_adj_4100));
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1369 (.I0(n15015), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [4]), .I3(n14536), .O(Kp_23__N_868));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i11620_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n16159));
    defparam i11620_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n15514), .D(n29640));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n15514), .D(n25004));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n15514), .D(n28293));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n15514), .D(n30114));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n15514), .D(n28105));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n15514), .D(n28851));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n15514), .D(n29993));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n15514), .D(n29713));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n15514), .D(n29188));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n15514), .D(n28209));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n15514), .D(n29733));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n15514), .D(n27906));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n15514), .D(n29643));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n15514), .D(n28199));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n15514), .D(n29802));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[13] [5]), 
            .I2(Kp_23__N_1446), .I3(\data_in_frame[15] [7]), .O(n28114));
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1371 (.I0(n30020), .I1(n15114), .I2(n10_adj_4148), 
            .I3(n29657), .O(n18_adj_4161));
    defparam i2_4_lut_adj_1371.LUT_INIT = 16'hbeeb;
    SB_LUT4 i2_3_lut_4_lut_adj_1372 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(n28448), .I3(n14593), .O(n26276));
    defparam i2_3_lut_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(\data_in_frame[10] [7]), .I1(Kp_23__N_1094), 
            .I2(\data_in_frame[8] [7]), .I3(GND_net), .O(n28448));
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n27137), .S(n27219));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n27840), .S(n27139));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n27839), .S(n27215));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n27838), .S(n27213));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n27837), .S(n27211));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n27835), .S(n27207));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n27836), .S(n27209));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n27855), .S(n8_adj_4162));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n27834), .S(n27205));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n88), .S(n8_adj_4163));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n19123), .S(n19636));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n19125), .S(n19638));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n27854), .S(n27201));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n27853), .S(n27199));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n19127), .S(n19642));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n27845), .S(n27203));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n27844), .S(n27237));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n27843), .S(n27027));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n27842), .S(n27235));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n27841), .S(n27233));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n27852), .S(n27159));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n27851), .S(n27197));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n27850), .S(n27195));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n27849), .S(n27193));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n27848), .S(n27191));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n27847), .S(n27189));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n27846), .S(n27187));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n19157), .S(n19660));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_4156), .S(n8_adj_4164));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n15481), .D(n8825[0]), .R(n15614));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .E(n28769), 
            .D(n4561), .R(n29468));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11621_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n16160));
    defparam i11621_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11622_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n16161));
    defparam i11622_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11623_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n16162));
    defparam i11623_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11624_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n16163));
    defparam i11624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11625_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n16164));
    defparam i11625_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(n15021), .I1(\data_in_frame[10] [5]), 
            .I2(n14542), .I3(GND_net), .O(n14632));
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_LUT4 i11626_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n16165));
    defparam i11626_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1375 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[16] [6]), 
            .I2(n29382), .I3(n26272), .O(n26326));
    defparam i2_3_lut_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i11627_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27867), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n16166));
    defparam i11627_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1376 (.I0(\data_out_frame[12] [7]), .I1(n28014), 
            .I2(n14347), .I3(GND_net), .O(n26451));
    defparam i1_2_lut_4_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1377 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(n28014), .I3(n14347), .O(n25294));
    defparam i2_3_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n7_adj_4095));
    defparam i18_4_lut_3_lut.LUT_INIT = 16'h1414;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n27796), .D(n15605), 
            .R(n29767));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n6_adj_4094));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1379 (.I0(n14593), .I1(\data_in_frame[10] [5]), 
            .I2(\data_in_frame[12] [7]), .I3(n14542), .O(n15317));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1380 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [7]), 
            .I2(n14542), .I3(GND_net), .O(n28345));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_LUT4 i11612_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n16151));
    defparam i11612_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1381 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [7]), 
            .I2(n28201), .I3(GND_net), .O(n10_adj_4091));
    defparam i2_2_lut_3_lut_adj_1381.LUT_INIT = 16'h9696;
    SB_LUT4 i11613_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n16152));
    defparam i11613_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1382 (.I0(\data_in_frame[9] [4]), .I1(n26320), 
            .I2(n28261), .I3(\data_in_frame[13] [6]), .O(n28201));
    defparam i1_2_lut_4_lut_adj_1382.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[2] [7]), .I3(GND_net), .O(n28027));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26169 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n32005));
    defparam byte_transmit_counter_0__bdd_4_lut_26169.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1384 (.I0(\data_out_frame[5] [4]), .I1(n10_adj_4086), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[5] [1]), .O(n28168));
    defparam i5_3_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1385 (.I0(\data_out_frame[14] [2]), .I1(n29737), 
            .I2(\data_out_frame[12] [2]), .I3(GND_net), .O(n26337));
    defparam i1_2_lut_3_lut_adj_1385.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(n26471), .I3(\data_out_frame[23] [4]), .O(n7_adj_4026));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(\data_out_frame[18] [7]), .I1(n28120), 
            .I2(n28488), .I3(GND_net), .O(n6_adj_4082));
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'h9696;
    SB_LUT4 i11614_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n16153));
    defparam i11614_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11615_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n16154));
    defparam i11615_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(n26333), .I1(n29704), .I2(\data_out_frame[15] [3]), 
            .I3(GND_net), .O(n15253));
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h6969;
    SB_LUT4 i11616_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n16155));
    defparam i11616_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32_3_lut_4_lut (.I0(\data_in_frame[14] [1]), .I1(n64), .I2(\data_in_frame[17] [7]), 
            .I3(\data_in_frame[17] [6]), .O(n74));
    defparam i32_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11617_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n16156));
    defparam i11617_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(n14164), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n14304));   // verilog/coms.v(263[5:27])
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'hfefe;
    SB_LUT4 i11618_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n16157));
    defparam i11618_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11619_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27867), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n16158));
    defparam i11619_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11604_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n16143));
    defparam i11604_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11605_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n16144));
    defparam i11605_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11606_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n16145));
    defparam i11606_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11607_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n16146));
    defparam i11607_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1389 (.I0(n29581), .I1(\data_out_frame[24] [2]), 
            .I2(\data_out_frame[24] [1]), .I3(n28292), .O(n28293));
    defparam i1_2_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(n4452), .I1(n9411), .I2(n14328), 
            .I3(GND_net), .O(n87));   // verilog/coms.v(259[6] 261[9])
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_4_lut_adj_1391 (.I0(n26333), .I1(n28179), .I2(n14931), 
            .I3(\data_out_frame[17] [5]), .O(n14395));
    defparam i1_2_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i11608_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n16147));
    defparam i11608_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1392 (.I0(n29699), .I1(n1581), .I2(\data_out_frame[13] [3]), 
            .I3(\data_out_frame[15] [5]), .O(n26290));
    defparam i2_3_lut_4_lut_adj_1392.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_4_lut_adj_1393 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[17] [4]), .I3(n15253), .O(n7_adj_4077));
    defparam i2_2_lut_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 n32005_bdd_4_lut (.I0(n32005), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n32008));
    defparam n32005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(n29699), .I1(\data_out_frame[13] [5]), 
            .I2(n26375), .I3(GND_net), .O(n26455));
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'h9696;
    SB_LUT4 i11609_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n16148));
    defparam i11609_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11610_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n16149));
    defparam i11610_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11611_3_lut_4_lut (.I0(n19694), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n16150));
    defparam i11611_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1395 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n14316), .I3(GND_net), .O(n14318));   // verilog/coms.v(222[5:21])
    defparam i1_2_lut_3_lut_adj_1395.LUT_INIT = 16'hfbfb;
    SB_LUT4 i10_4_lut_adj_1396 (.I0(n29303), .I1(n29156), .I2(n29325), 
            .I3(n29351), .O(n26_adj_4165));
    defparam i10_4_lut_adj_1396.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1397 (.I0(n12524), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[10] [4]), .I3(n14719), .O(n14347));
    defparam i2_3_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1398 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n19172), .O(n27874));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1398.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(n14164), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n14316));   // verilog/coms.v(231[5:23])
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_4_lut_adj_1400 (.I0(n14727), .I1(n28241), .I2(n14395), 
            .I3(n28104), .O(n28105));
    defparam i1_2_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1401 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n19172), .O(n27883));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1401.LUT_INIT = 16'hefff;
    SB_LUT4 i11596_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n16135));
    defparam i11596_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_94_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4166));
    defparam equal_94_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1402 (.I0(\data_out_frame[9] [4]), .I1(n28313), 
            .I2(\data_out_frame[15] [7]), .I3(\data_out_frame[15] [6]), 
            .O(n28034));
    defparam i1_2_lut_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut_4_lut (.I0(n15021), .I1(\data_in_frame[5] [5]), .I2(n27984), 
            .I3(n28017), .O(n24_adj_4063));
    defparam i8_3_lut_4_lut.LUT_INIT = 16'hbeeb;
    SB_LUT4 i11597_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n16136));
    defparam i11597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11598_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n16137));
    defparam i11598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1403 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(n28460), .O(n8_adj_4061));   // verilog/coms.v(78[16:27])
    defparam i3_3_lut_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i11599_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n16138));
    defparam i11599_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11600_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n16139));
    defparam i11600_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11601_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n16140));
    defparam i11601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1404 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(n28396), .O(n8_adj_4060));
    defparam i3_3_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(GND_net), .O(n28460));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i11602_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n16141));
    defparam i11602_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1406 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [6]), .I3(n14705), .O(n28399));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i11603_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n16142));
    defparam i11603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11588_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n16127));
    defparam i11588_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11589_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n16128));
    defparam i11589_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15154_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n19694));
    defparam i15154_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i11590_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n16129));
    defparam i11590_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1407 (.I0(\data_out_frame[13] [7]), .I1(n1581), 
            .I2(n29701), .I3(GND_net), .O(n28451));
    defparam i1_2_lut_3_lut_adj_1407.LUT_INIT = 16'h6969;
    SB_LUT4 i11591_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n16130));
    defparam i11591_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1408 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[7] [3]), .O(n27970));
    defparam i1_2_lut_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1409 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[18] [7]), .I3(\data_out_frame[18] [6]), 
            .O(n28408));
    defparam i1_2_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i11592_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n16131));
    defparam i11592_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11593_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n16132));
    defparam i11593_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1410 (.I0(n26326), .I1(n10_adj_4028), .I2(n14515), 
            .I3(n2076), .O(n26270));
    defparam i5_3_lut_4_lut_adj_1410.LUT_INIT = 16'h9669;
    SB_LUT4 i11594_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n16133));
    defparam i11594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1411 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n15015));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i11595_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n16134));
    defparam i11595_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11580_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n16119));
    defparam i11580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1412 (.I0(\data_out_frame[20] [3]), .I1(n14030), 
            .I2(n25359), .I3(\data_out_frame[24] [5]), .O(n28367));
    defparam i1_2_lut_3_lut_4_lut_adj_1412.LUT_INIT = 16'h9669;
    SB_LUT4 i11581_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n16120));
    defparam i11581_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(n26365), .I1(\data_out_frame[23] [2]), 
            .I2(n25268), .I3(GND_net), .O(n28233));
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i11582_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n16121));
    defparam i11582_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11583_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n16122));
    defparam i11583_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11584_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n16123));
    defparam i11584_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1414 (.I0(n29867), .I1(n25305), .I2(\data_out_frame[25] [5]), 
            .I3(\data_out_frame[25] [4]), .O(n28199));
    defparam i1_2_lut_4_lut_adj_1414.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1415 (.I0(\FRAME_MATCHER.state [3]), .I1(n9411), 
            .I2(n23), .I3(n87), .O(n27137));
    defparam i1_3_lut_4_lut_adj_1415.LUT_INIT = 16'haa08;
    SB_LUT4 i1_2_lut_3_lut_adj_1416 (.I0(n14295), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n14309));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_adj_1416.LUT_INIT = 16'hefef;
    SB_LUT4 i11585_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n16124));
    defparam i11585_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1417 (.I0(n19172), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n27867));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1417.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1418 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n14292), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_4020));
    defparam i1_3_lut_4_lut_adj_1418.LUT_INIT = 16'hfefc;
    SB_LUT4 i11586_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n16125));
    defparam i11586_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1519_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_3997));
    defparam i1519_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i11587_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n16126));
    defparam i11587_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11572_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n16111));
    defparam i11572_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11573_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n16112));
    defparam i11573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11574_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n16113));
    defparam i11574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11575_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n16114));
    defparam i11575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11576_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n16115));
    defparam i11576_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11577_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n16116));
    defparam i11577_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1419 (.I0(n29199), .I1(n28_adj_4155), .I2(n22_adj_4154), 
            .I3(n29177), .O(n30_adj_4167));
    defparam i14_4_lut_adj_1419.LUT_INIT = 16'hfeff;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26164 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n31999));
    defparam byte_transmit_counter_0__bdd_4_lut_26164.LUT_INIT = 16'he4aa;
    SB_LUT4 n31999_bdd_4_lut (.I0(n31999), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n32002));
    defparam n31999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1420 (.I0(\data_in_frame[21] [0]), .I1(n29496), 
            .I2(n8_adj_4158), .I3(n14967), .O(n17_adj_4168));
    defparam i1_4_lut_adj_1420.LUT_INIT = 16'hdeed;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_26242 (.I0(byte_transmit_counter[1]), 
            .I1(n31103), .I2(n31104), .I3(byte_transmit_counter[2]), .O(n31993));
    defparam byte_transmit_counter_1__bdd_4_lut_26242.LUT_INIT = 16'he4aa;
    SB_LUT4 n31993_bdd_4_lut (.I0(n31993), .I1(n17_adj_3891), .I2(n16_adj_3890), 
            .I3(byte_transmit_counter[2]), .O(n31996));
    defparam n31993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15_4_lut_adj_1421 (.I0(n17_adj_4168), .I1(n30_adj_4167), .I2(n26_adj_4165), 
            .I3(n18_adj_4161), .O(n31_adj_4068));
    defparam i15_4_lut_adj_1421.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_26154 (.I0(byte_transmit_counter[1]), 
            .I1(n31106), .I2(n31107), .I3(byte_transmit_counter[2]), .O(n31987));
    defparam byte_transmit_counter_1__bdd_4_lut_26154.LUT_INIT = 16'he4aa;
    SB_LUT4 n31987_bdd_4_lut (.I0(n31987), .I1(n17_adj_3889), .I2(n16_adj_3888), 
            .I3(byte_transmit_counter[2]), .O(n31990));
    defparam n31987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11578_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n16117));
    defparam i11578_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_26149 (.I0(byte_transmit_counter[1]), 
            .I1(n31109), .I2(n31110), .I3(byte_transmit_counter[2]), .O(n31981));
    defparam byte_transmit_counter_1__bdd_4_lut_26149.LUT_INIT = 16'he4aa;
    SB_LUT4 n31981_bdd_4_lut (.I0(n31981), .I1(n17_adj_3887), .I2(n16_adj_3886), 
            .I3(byte_transmit_counter[2]), .O(n31984));
    defparam n31981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_26144 (.I0(byte_transmit_counter[1]), 
            .I1(n31115), .I2(n31116), .I3(byte_transmit_counter[2]), .O(n31975));
    defparam byte_transmit_counter_1__bdd_4_lut_26144.LUT_INIT = 16'he4aa;
    SB_LUT4 n31975_bdd_4_lut (.I0(n31975), .I1(n17_adj_3885), .I2(n16_adj_3884), 
            .I3(byte_transmit_counter[2]), .O(n31978));
    defparam n31975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_26139 (.I0(byte_transmit_counter[1]), 
            .I1(n31151), .I2(n31152), .I3(byte_transmit_counter[2]), .O(n31969));
    defparam byte_transmit_counter_1__bdd_4_lut_26139.LUT_INIT = 16'he4aa;
    SB_LUT4 n31969_bdd_4_lut (.I0(n31969), .I1(n17_adj_3883), .I2(n16_adj_3881), 
            .I3(byte_transmit_counter[2]), .O(n31972));
    defparam n31969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_26134 (.I0(byte_transmit_counter[1]), 
            .I1(n31097), .I2(n31098), .I3(byte_transmit_counter[2]), .O(n31963));
    defparam byte_transmit_counter_1__bdd_4_lut_26134.LUT_INIT = 16'he4aa;
    SB_LUT4 n31963_bdd_4_lut (.I0(n31963), .I1(n17), .I2(n16), .I3(byte_transmit_counter[2]), 
            .O(n31966));
    defparam n31963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n15507), .D(n4525));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11579_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n16118));
    defparam i11579_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11564_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n16103));
    defparam i11564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26159 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n31951));
    defparam byte_transmit_counter_0__bdd_4_lut_26159.LUT_INIT = 16'he4aa;
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n15507), .D(n4526));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n31951_bdd_4_lut (.I0(n31951), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n31954));
    defparam n31951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_26121 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n31945));
    defparam byte_transmit_counter_0__bdd_4_lut_26121.LUT_INIT = 16'he4aa;
    SB_LUT4 n31945_bdd_4_lut (.I0(n31945), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n31948));
    defparam n31945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1422 (.I0(n9411), .I1(n3303), .I2(n14316), 
            .I3(GND_net), .O(n6_adj_3995));   // verilog/coms.v(227[6] 229[9])
    defparam i1_2_lut_3_lut_adj_1422.LUT_INIT = 16'h0202;
    SB_LUT4 i11565_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n16104));
    defparam i11565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(n9411), .I1(n3303), .I2(n14318), 
            .I3(GND_net), .O(n81));   // verilog/coms.v(227[6] 229[9])
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h0202;
    SB_LUT4 i11566_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n16105));
    defparam i11566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11567_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n16106));
    defparam i11567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_91_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4160));   // verilog/coms.v(154[7:23])
    defparam equal_91_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i11568_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n16107));
    defparam i11568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_92_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3996));   // verilog/coms.v(154[7:23])
    defparam equal_92_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11569_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n16108));
    defparam i11569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1424 (.I0(n81), .I1(n41_adj_3988), .I2(n1), 
            .I3(\FRAME_MATCHER.state [31]), .O(n8_adj_4164));
    defparam i1_2_lut_4_lut_adj_1424.LUT_INIT = 16'hfe00;
    SB_LUT4 i11570_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n16109));
    defparam i11570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11571_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n16110));
    defparam i11571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n15507), .D(n4527));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n15507), .D(n4528));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n15507), .D(n4529));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n15507), .D(n4530));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n15507), .D(n4531));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n15507), .D(n4532));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n15507), .D(n4533));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n15507), 
            .D(n4534));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n15507), 
            .D(n4535));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n15507), 
            .D(n4536));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n15507), 
            .D(n4537));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n15507), 
            .D(n4538));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n15507), 
            .D(n4539));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n15507), 
            .D(n4540));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n15507), 
            .D(n4541));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n15507), 
            .D(n4542));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n15507), 
            .D(n4543));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n15507), 
            .D(n4544));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n15507), 
            .D(n4545));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n15507), 
            .D(n4546));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n15507), 
            .D(n4547));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1425 (.I0(\data_in_frame[6] [0]), .I1(Kp_23__N_810), 
            .I2(n14548), .I3(GND_net), .O(n14493));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1425.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1426 (.I0(\data_in_frame[6] [0]), .I1(Kp_23__N_810), 
            .I2(n28230), .I3(n12761), .O(n29381));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1426.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_4_lut_adj_1427 (.I0(Kp_23__N_979), .I1(n28011), .I2(\data_in_frame[6] [5]), 
            .I3(\data_in_frame[8] [6]), .O(n8_adj_4065));   // verilog/coms.v(76[16:43])
    defparam i2_2_lut_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1428 (.I0(Kp_23__N_979), .I1(n28011), .I2(\data_in_frame[6] [5]), 
            .I3(Kp_23__N_1094), .O(n28068));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i15121_2_lut_4_lut (.I0(n81), .I1(n41_adj_3988), .I2(n1), 
            .I3(\FRAME_MATCHER.state [30]), .O(n19660));
    defparam i15121_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i15104_2_lut_4_lut (.I0(n81), .I1(n41_adj_3988), .I2(n1), 
            .I3(\FRAME_MATCHER.state [17]), .O(n19642));
    defparam i15104_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i11556_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n16095));
    defparam i11556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11557_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n16096));
    defparam i11557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11558_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n16097));
    defparam i11558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11559_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n16098));
    defparam i11559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n32531));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state[1] ), .C(clk32MHz), 
           .D(n32532));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11560_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n16099));
    defparam i11560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n16232));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n16231));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n16230));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n16229));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11561_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n16100));
    defparam i11561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n16228));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n16227));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n16226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n16225));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n16224));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n16223));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n16222));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n16221));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n16220));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n16219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n16218));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n16217));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n16216));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n16215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n16214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n16213));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11562_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n16101));
    defparam i11562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n16212));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n16211));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n16210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n16209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n16208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n16207));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n16206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n16205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n16204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n16199));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n16198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n16197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n16196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n16195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n16194));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n16193));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n16192));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n16191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n16190));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n16189));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11563_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n16102));
    defparam i11563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n16188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n16187));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n16186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n16185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n16184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n16183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n16182));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n16181));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n16180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n16179));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n16178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n16177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n16176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n16175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n16174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n16173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n16172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n16171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n16170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n16169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n16168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n16167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n16166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n16165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n16164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n16163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n16162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n16161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n16160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n16159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n16158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n16157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n16156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n16155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n16154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n16153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n16152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n16151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n16150));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n16149));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n16148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n16147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n16146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n16145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n16144));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n16143));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n16142));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n16141));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n16140));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n16139));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n16138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n16137));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n16136));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n16135));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n16134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n16133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n16132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n16131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n16130));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n16129));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n16128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n16127));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n16126));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n16125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n16124));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n16123));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n16122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n16121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n16120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n16119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n16118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n16117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n16116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n16115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n16114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n16113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n16112));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n16111));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n16110));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n16109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n16108));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n16107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n16106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n16105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n16104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n16103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n16102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n16101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n16100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n16099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n16098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n16097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n16096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n16095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n16094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n16093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n16092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n16091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n16090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n16089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n16088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n16087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n16086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n16085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n16084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n16083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n16082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n16081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n16080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n16079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n16078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n16077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n16076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n16075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n16074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n16073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n16072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n16071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n16070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n16069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n16068));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1429 (.I0(tx_active), .I1(r_SM_Main_2__N_3496[0]), 
            .I2(n19835), .I3(GND_net), .O(n7_adj_4114));
    defparam i2_2_lut_3_lut_adj_1429.LUT_INIT = 16'hfefe;
    SB_LUT4 i15102_2_lut_4_lut (.I0(n81), .I1(n41_adj_3988), .I2(n1), 
            .I3(\FRAME_MATCHER.state [14]), .O(n19638));
    defparam i15102_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1430 (.I0(tx_active), .I1(r_SM_Main_2__N_3496[0]), 
            .I2(n14327), .I3(tx_transmit_N_3393), .O(n27831));
    defparam i1_2_lut_3_lut_4_lut_adj_1430.LUT_INIT = 16'h0f0e;
    SB_LUT4 i26012_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3496[0]), 
            .I2(n14327), .I3(n63_adj_3), .O(n15481));
    defparam i26012_3_lut_4_lut.LUT_INIT = 16'h01ff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1431 (.I0(tx_active), .I1(r_SM_Main_2__N_3496[0]), 
            .I2(n9411), .I3(tx_transmit_N_3393), .O(n11873));
    defparam i1_2_lut_3_lut_4_lut_adj_1431.LUT_INIT = 16'hf0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1432 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(n28399), .I3(\data_in_frame[1] [4]), .O(n14499));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1433 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[8] [0]), .O(n28061));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1434 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(n15247), .I3(\data_in_frame[0] [5]), .O(n28390));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n15034));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1436 (.I0(n14295), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n14328));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_adj_1436.LUT_INIT = 16'hbfbf;
    SB_LUT4 i22830_2_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n14164), .I3(GND_net), .O(n28649));
    defparam i22830_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n16067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n16066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n16065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n16064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n16063));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n16062));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n16061));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n16060));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n16059));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n16058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n16057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n16056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n16055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n16054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n16053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n16052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n16051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n16050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n16049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n16048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n16047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n16046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n16045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n16044));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n16043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n16042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n16041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n16040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n16039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n16038));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n16037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n16036));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n16035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n16034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n16033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n16032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n16031));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n16030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n16029));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n16028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n16027));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n16026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n16025));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n16024));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n16023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n16022));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n16021));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n16020));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n16019));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n16018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n16017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n16016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n16015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n16014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n16013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n16012));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n16011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n16010));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n16009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n16008));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n16007));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n16006));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n16005));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n16004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n16003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n16002));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n16001));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n16000));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n15999));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n15998));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n15997));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n15996));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n15995));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n15994));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n15993));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n15992));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n15991));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n15990));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n15989));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n15988));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n15987));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n15986));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n15985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n15984));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n15983));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n15982));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n15981));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n15980));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n15979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n15978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n15977));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n15976));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n15975));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n15974));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n15973));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n15972));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n15971));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n15970));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n15969));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n15968));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n15967));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n15966));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n15965));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n15964));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n15963));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n15962));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n15961));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n15960));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n15959));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n15958));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n15957));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n15956));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n15955));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n15954));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n15953));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1437 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[6] [7]), .I3(\data_in_frame[0] [5]), .O(n10_adj_4108));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i11548_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n16087));
    defparam i11548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15101_2_lut_4_lut (.I0(n81), .I1(n41_adj_3988), .I2(n1), 
            .I3(\FRAME_MATCHER.state [13]), .O(n19636));
    defparam i15101_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i11549_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n16088));
    defparam i11549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11550_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n16089));
    defparam i11550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n15952));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n15951));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n15950));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n15949));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n15948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n15947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n15946));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n15945));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n15944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n15943));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11551_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n16090));
    defparam i11551_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n15942));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n15941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n15940));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n15939));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n15938));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n15937));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n15936));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n15935));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11552_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n16091));
    defparam i11552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n15934));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n15933));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n15932));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n15931));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n15930));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n15929));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n15928));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11553_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n16092));
    defparam i11553_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n15927));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n15926));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n15925));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n15924));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n15923));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n15922));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n15921));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n15920));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n15919));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n15918));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n15917));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n15916));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n15915));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n15914));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n15913));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n15912));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n15911));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n15910));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n15909));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n15908));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n15907));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n15906));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1438 (.I0(n81), .I1(n41_adj_3988), .I2(n1), 
            .I3(\FRAME_MATCHER.state [12]), .O(n8_adj_4163));
    defparam i1_2_lut_4_lut_adj_1438.LUT_INIT = 16'hfe00;
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n15905));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n15904));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n15903));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n15902));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n15901));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1439 (.I0(n63), .I1(n3303), .I2(n123), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2668[1] ));
    defparam i2_3_lut_adj_1439.LUT_INIT = 16'hfdfd;
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n15900));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11554_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n16093));
    defparam i11554_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11555_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27883), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n16094));
    defparam i11555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11540_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n16079));
    defparam i11540_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11541_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n16080));
    defparam i11541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1440 (.I0(n81), .I1(n41_adj_3988), .I2(n1), 
            .I3(\FRAME_MATCHER.state [10]), .O(n8_adj_4162));
    defparam i1_2_lut_4_lut_adj_1440.LUT_INIT = 16'hfe00;
    SB_LUT4 i11542_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n16081));
    defparam i11542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n15899));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n15898));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n15897));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n15896));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n15895));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11543_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n16082));
    defparam i11543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11544_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n16083));
    defparam i11544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11545_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n16084));
    defparam i11545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11546_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n16085));
    defparam i11546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11547_3_lut_4_lut (.I0(n19694), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n16086));
    defparam i11547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i26028_4_lut_4_lut (.I0(n14332), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n19871), .I3(n14279), .O(n29767));
    defparam i26028_4_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i4056_2_lut (.I0(n63), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n8515));   // verilog/coms.v(157[6] 159[9])
    defparam i4056_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1441 (.I0(\FRAME_MATCHER.state [2]), .I1(n1_adj_3989), 
            .I2(n32_adj_4143), .I3(GND_net), .O(n122));
    defparam i1_3_lut_adj_1441.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_366_Select_2_i5_4_lut (.I0(n122), .I1(n14318), .I2(n3303), 
            .I3(n63), .O(n5));
    defparam select_366_Select_2_i5_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i14799_rep_305_2_lut (.I0(n122), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n32898));   // verilog/coms.v(142[4] 144[7])
    defparam i14799_rep_305_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26060_3_lut_4_lut (.I0(n14332), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n28763), .I3(\FRAME_MATCHER.state [3]), .O(n29468));
    defparam i26060_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i22938_3_lut_4_lut (.I0(n14332), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n19871), .I3(\FRAME_MATCHER.state [3]), .O(n28763));
    defparam i22938_3_lut_4_lut.LUT_INIT = 16'hfef0;
    SB_LUT4 i1_2_lut_3_lut_adj_1442 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n14638));
    defparam i1_2_lut_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1443 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(n14756), .I3(GND_net), .O(n26346));
    defparam i1_2_lut_3_lut_adj_1443.LUT_INIT = 16'h9696;
    SB_LUT4 i11532_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n16071));
    defparam i11532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11533_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n16072));
    defparam i11533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11534_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n16073));
    defparam i11534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11535_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n16074));
    defparam i11535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11536_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n16075));
    defparam i11536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11537_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n16076));
    defparam i11537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11538_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n16077));
    defparam i11538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11539_3_lut_4_lut (.I0(n8_adj_4166), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n16078));
    defparam i11539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24460_2_lut_4_lut (.I0(n63), .I1(n18546), .I2(n14313), .I3(n1_adj_3989), 
            .O(n30290));
    defparam i24460_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1444 (.I0(n29704), .I1(n1581), .I2(\data_out_frame[13] [3]), 
            .I3(\data_out_frame[15] [4]), .O(n14931));
    defparam i1_2_lut_3_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(n29704), .I1(n1581), .I2(\data_out_frame[13] [3]), 
            .I3(n28417), .O(n18_adj_4047));
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1445 (.I0(\data_in_frame[0] [5]), .I1(Kp_23__N_868), 
            .I2(n28027), .I3(GND_net), .O(n14845));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1445.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1446 (.I0(\data_in_frame[0] [5]), .I1(Kp_23__N_868), 
            .I2(\data_in_frame[2] [6]), .I3(n28089), .O(n15247));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i26065_2_lut_3_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n15605));
    defparam i26065_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i2_4_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state_31__N_2604 [3]), 
            .O(n6_adj_3986));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha0a4;
    SB_LUT4 i14833_2_lut_4_lut (.I0(n12002), .I1(n31_adj_4068), .I2(n31_adj_4056), 
            .I3(\FRAME_MATCHER.state[1] ), .O(n1_adj_4151));
    defparam i14833_2_lut_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i11524_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n16063));
    defparam i11524_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11525_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n16064));
    defparam i11525_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11526_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n16065));
    defparam i11526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11527_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n16066));
    defparam i11527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1447 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[5] [0]), .I3(n13958), .O(n25261));
    defparam i1_2_lut_3_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i11528_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n16067));
    defparam i11528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11529_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n16068));
    defparam i11529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11530_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n16069));
    defparam i11530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11531_3_lut_4_lut (.I0(n8_adj_4116), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n16070));
    defparam i11531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1448 (.I0(n14588), .I1(n10_adj_4066), .I2(\data_in_frame[9] [2]), 
            .I3(GND_net), .O(n14561));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_1448.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1449 (.I0(n14588), .I1(n10_adj_4066), .I2(n26320), 
            .I3(\data_in_frame[9] [4]), .O(n28527));   // verilog/coms.v(72[16:41])
    defparam i1_3_lut_4_lut_adj_1449.LUT_INIT = 16'h9669;
    SB_LUT4 i11516_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n16055));
    defparam i11516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11517_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n16056));
    defparam i11517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11518_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n16057));
    defparam i11518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11519_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n16058));
    defparam i11519_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i26017_2_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n7_adj_4095), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n19871), .O(n15514));   // verilog/coms.v(127[12] 300[6])
    defparam i26017_2_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i11520_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n16059));
    defparam i11520_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(n26352), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[12] [5]), .I3(n14895), .O(n6_adj_3892));
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i11521_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n16060));
    defparam i11521_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n27243));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n15719));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n15894));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n15893));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n15892));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n15891));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n15890));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n15889));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n15888));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n15887));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n15886));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n15885));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1451 (.I0(n26281), .I1(\data_out_frame[10] [1]), 
            .I2(n30022), .I3(n28479), .O(n28213));
    defparam i1_2_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1452 (.I0(n26352), .I1(n12524), .I2(n28020), 
            .I3(n14719), .O(n28479));
    defparam i1_2_lut_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n15884));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n15883));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n15882));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n15881));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n15880));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n15879));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n15878));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n15877));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n15876));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n15875));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n15874));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n15873));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n15872));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n15871));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n15870));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n15869));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n15868));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n15867));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n15866));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n15865));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n15864));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n15863));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n15862));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n15718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n15717));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n15716));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n15715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n15714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n15713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n15861));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n15860));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n15859));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n15858));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n15857));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n15856));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n15855));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11522_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n16061));
    defparam i11522_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n15705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n15854));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n15853));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n15852));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n15851));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n15850));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n15849));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n15848));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n15847));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11523_3_lut_4_lut (.I0(n8_adj_4130), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n16062));
    defparam i11523_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1453 (.I0(n14719), .I1(\data_out_frame[8] [1]), 
            .I2(n25814), .I3(\data_out_frame[10] [3]), .O(n26352));
    defparam i2_3_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n15846));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n15845));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n15844));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n15843));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n15842));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1454 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[1] [3]), .I3(n10_adj_4104), .O(n14542));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1455 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [1]), 
            .I2(n28411), .I3(n28159), .O(Kp_23__N_810));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i11508_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n16047));
    defparam i11508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1456 (.I0(n13958), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[7] [5]), .O(n25290));
    defparam i2_3_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i11509_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n16048));
    defparam i11509_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n28041));
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1458 (.I0(n28224), .I1(\data_out_frame[23] [7]), 
            .I2(n14727), .I3(GND_net), .O(n28292));
    defparam i1_2_lut_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1459 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[7] [4]), .I3(\data_out_frame[9] [4]), .O(n28438));
    defparam i2_3_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i11510_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n16049));
    defparam i11510_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1460 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [2]), .I3(n28210), .O(n6_adj_3879));
    defparam i1_2_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i11511_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n16050));
    defparam i11511_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11512_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n16051));
    defparam i11512_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11513_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n16052));
    defparam i11513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n14316), 
            .I2(n14295), .I3(n43), .O(n23));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hff2a;
    SB_LUT4 i11514_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n16053));
    defparam i11514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1461 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [2]), .I3(GND_net), .O(n14612));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1461.LUT_INIT = 16'h9696;
    SB_LUT4 i11515_3_lut_4_lut (.I0(n8_adj_4142), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n16054));
    defparam i11515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n15841));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1462 (.I0(\data_in_frame[15] [4]), .I1(n28521), 
            .I2(\data_in_frame[13] [3]), .I3(n28539), .O(n6_adj_4159));
    defparam i1_2_lut_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1463 (.I0(\data_in_frame[15] [4]), .I1(n28521), 
            .I2(\data_in_frame[13] [3]), .I3(n28482), .O(n6_adj_4092));
    defparam i1_2_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n15840));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14_3_lut_4_lut (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(n27905), .I3(n28_adj_4045), .O(n32_adj_4052));   // verilog/coms.v(71[16:27])
    defparam i14_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1464 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(n25712), .I3(n28204), .O(n29910));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1464.LUT_INIT = 16'h9669;
    SB_LUT4 i11500_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n16039));
    defparam i11500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11501_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n16040));
    defparam i11501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11502_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n16041));
    defparam i11502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11503_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n16042));
    defparam i11503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[8] [1]), 
            .I2(n27949), .I3(\data_out_frame[8] [2]), .O(n18));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11504_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n16043));
    defparam i11504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11505_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n16044));
    defparam i11505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1465 (.I0(n28057), .I1(\data_in_frame[11] [6]), 
            .I2(n28017), .I3(\data_in_frame[7] [1]), .O(n27));   // verilog/coms.v(85[17:70])
    defparam i11_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut_4_lut_adj_1466 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[6] [0]), 
            .I2(n15416), .I3(n1265), .O(n15_adj_4085));   // verilog/coms.v(85[17:70])
    defparam i5_2_lut_3_lut_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i11506_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n16045));
    defparam i11506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11507_3_lut_4_lut (.I0(n8_adj_4157), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n16046));
    defparam i11507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n15839));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1467 (.I0(\data_out_frame[11] [7]), .I1(n26281), 
            .I2(n4_adj_4037), .I3(GND_net), .O(n15279));
    defparam i2_2_lut_3_lut_adj_1467.LUT_INIT = 16'h9696;
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n15838));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n15837));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n15836));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n15835));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n15834));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n15833));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n15832));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n15831));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n15830));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n15829));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n15828));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n15827));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11492_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n16031));
    defparam i11492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11493_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n16032));
    defparam i11493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11494_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n16033));
    defparam i11494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n15826));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n15825));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n15824));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n15823));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n15822));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n15821));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n15820));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n15819));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3][7] ), .C(clk32MHz), .D(n15818));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11495_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n16034));
    defparam i11495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i31 (.Q(\data_in[3][6] ), .C(clk32MHz), .D(n15817));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n15816));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3][4] ), .C(clk32MHz), .D(n15815));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3][3] ), .C(clk32MHz), .D(n15814));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3][2] ), .C(clk32MHz), .D(n15813));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3][1] ), .C(clk32MHz), .D(n15812));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11496_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n16035));
    defparam i11496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11497_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n16036));
    defparam i11497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11498_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n16037));
    defparam i11498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1468 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(\data_out_frame[5] [7]), .O(n25814));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i25 (.Q(\data_in[3][0] ), .C(clk32MHz), .D(n15811));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n15810));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n15809));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n15808));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n15807));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n15806));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n15805));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n15804));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11499_3_lut_4_lut (.I0(n8_adj_4160), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n16038));
    defparam i11499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n15803));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n15802));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n15801));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n15800));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n15799));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n15798));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n15797));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_3_lut (.I0(\data_out_frame[6] [0]), .I1(n10), 
            .I2(n1265), .I3(GND_net), .O(n13958));   // verilog/coms.v(85[17:70])
    defparam i5_3_lut_4_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11178_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n15717));
    defparam i11178_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n15796));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1469 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [1]), 
            .I2(n1260), .I3(n28307), .O(n1265));
    defparam i2_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i11485_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n16024));
    defparam i11485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n15795));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11486_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n16025));
    defparam i11486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n15794));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n15793));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n15792));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n15791));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1470 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[5] [0]), .O(n28508));
    defparam i1_2_lut_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n15790));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11487_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n16026));
    defparam i11487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n15789));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1471 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n14987));
    defparam i1_2_lut_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1472 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n12524));
    defparam i1_2_lut_3_lut_adj_1472.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n15788));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11488_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n16027));
    defparam i11488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n15787));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n15786));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n15785));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1051_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4523), .I3(GND_net), .O(n4547));
    defparam mux_1051_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n15784));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11489_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n16028));
    defparam i11489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1051_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4523), .I3(GND_net), .O(n4546));
    defparam mux_1051_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4523), .I3(GND_net), .O(n4545));
    defparam mux_1051_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4523), .I3(GND_net), .O(n4544));
    defparam mux_1051_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4523), .I3(GND_net), .O(n4543));
    defparam mux_1051_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4523), .I3(GND_net), .O(n4542));
    defparam mux_1051_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4523), .I3(GND_net), .O(n4541));
    defparam mux_1051_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4523), .I3(GND_net), .O(n4540));
    defparam mux_1051_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11490_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n16029));
    defparam i11490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1051_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4523), .I3(GND_net), .O(n4539));
    defparam mux_1051_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11491_3_lut_4_lut (.I0(n8_adj_3996), .I1(n27874), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n16030));
    defparam i11491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1051_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4523), .I3(GND_net), .O(n4538));
    defparam mux_1051_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4523), .I3(GND_net), .O(n4537));
    defparam mux_1051_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4523), .I3(GND_net), .O(n4536));
    defparam mux_1051_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4523), .I3(GND_net), .O(n4535));
    defparam mux_1051_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4523), .I3(GND_net), .O(n4534));
    defparam mux_1051_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4523), .I3(GND_net), .O(n4533));
    defparam mux_1051_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4523), .I3(GND_net), .O(n4532));
    defparam mux_1051_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4523), .I3(GND_net), .O(n4531));
    defparam mux_1051_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4523), .I3(GND_net), .O(n4530));
    defparam mux_1051_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4523), .I3(GND_net), .O(n4529));
    defparam mux_1051_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4523), .I3(GND_net), .O(n4528));
    defparam mux_1051_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4523), .I3(GND_net), .O(n4527));
    defparam mux_1051_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1186));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1051_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4523), .I3(GND_net), .O(n4526));
    defparam mux_1051_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14049_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15808));   // verilog/coms.v(90[7:20])
    defparam i14049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1051_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4523), .I3(GND_net), .O(n4525));
    defparam mux_1051_i2_3_lut.LUT_INIT = 16'hcaca;
    uart_tx tx (.clk32MHz(clk32MHz), .GND_net(GND_net), .n28749(n28749), 
            .n28775(n28775), .VCC_net(VCC_net), .\r_SM_Main_2__N_3496[0] (r_SM_Main_2__N_3496[0]), 
            .r_SM_Main({r_SM_Main}), .n8353(n8353), .tx_o(tx_o), .tx_data({tx_data}), 
            .\r_SM_Main_2__N_3493[1] (\r_SM_Main_2__N_3493[1] ), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .n4(n4), .n15730(n15730), .n32553(n32553), .n15722(n15722), 
            .tx_active(tx_active), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.n15548(n15548), .clk32MHz(clk32MHz), .n15643(n15643), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\r_SM_Main_2__N_3422[2] (\r_SM_Main_2__N_3422[2] ), 
            .r_SM_Main({r_SM_Main_adj_11}), .n27820(n27820), .r_Rx_Data(r_Rx_Data), 
            .n19238(n19238), .n4(n4_adj_7), .n4_adj_1(n4_adj_8), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_9 ), 
            .n14287(n14287), .RX_N_2(RX_N_2), .n14282(n14282), .n4_adj_2(n4_adj_10), 
            .n27405(n27405), .rx_data_ready(rx_data_ready), .n15764(n15764), 
            .n16203(n16203), .rx_data({rx_data}), .n15712(n15712), .n15711(n15711), 
            .n15710(n15710), .n15709(n15709), .n15708(n15708), .n15707(n15707), 
            .n15706(n15706)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, GND_net, n28749, n28775, VCC_net, \r_SM_Main_2__N_3496[0] , 
            r_SM_Main, n8353, tx_o, tx_data, \r_SM_Main_2__N_3493[1] , 
            \r_Bit_Index[0] , n4, n15730, n32553, n15722, tx_active, 
            tx_enable) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    input GND_net;
    output n28749;
    output n28775;
    input VCC_net;
    input \r_SM_Main_2__N_3496[0] ;
    output [2:0]r_SM_Main;
    output n8353;
    output tx_o;
    input [7:0]tx_data;
    output \r_SM_Main_2__N_3493[1] ;
    output \r_Bit_Index[0] ;
    output n4;
    input n15730;
    input n32553;
    input n15722;
    output tx_active;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n15626, n24020;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n24021, n24019, n24018, n24017, n24016, n24015, n3, n11634;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n9640, n19702, n9639, n32038, n32110, o_Tx_Serial_N_3524, 
        n32107, n32035, n3_adj_3878, n10, n29690, n24022;
    
    SB_DFFESR r_Clock_Count_1197__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n1), .D(n41[8]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1197__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n1), .D(n41[7]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1197__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n1), .D(n41[6]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1197__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n1), .D(n41[5]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1197__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n1), .D(n41[4]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1197__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n1), .D(n41[3]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1197__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n1), .D(n41[2]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 r_Clock_Count_1197_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n24020), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n28749), 
            .D(n307[1]), .R(n28775));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY r_Clock_Count_1197_add_4_8 (.CI(n24020), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n24021));
    SB_LUT4 r_Clock_Count_1197_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n24019), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1197_add_4_7 (.CI(n24019), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n24020));
    SB_LUT4 r_Clock_Count_1197_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n24018), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1197_add_4_6 (.CI(n24018), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n24019));
    SB_LUT4 r_Clock_Count_1197_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n24017), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1197_add_4_5 (.CI(n24017), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n24018));
    SB_LUT4 r_Clock_Count_1197_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n24016), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1197_add_4_4 (.CI(n24016), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n24017));
    SB_LUT4 r_Clock_Count_1197_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n24015), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1197_add_4_3 (.CI(n24015), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n24016));
    SB_LUT4 r_Clock_Count_1197_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1197_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n24015));
    SB_LUT4 i3895_2_lut (.I0(\r_SM_Main_2__N_3496[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n8353));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i3895_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n9640), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3496[0] ), 
            .I3(r_SM_Main[1]), .O(n11634));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n28749), 
            .D(n307[2]), .R(n28775));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1197__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n1), .D(n41[0]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i26079_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3493[1] ), .O(n28749));
    defparam i26079_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n19702));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i26073_3_lut (.I0(n28749), .I1(n19702), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28775));
    defparam i26073_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1295_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1295_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1288_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1288_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5173_4_lut (.I0(\r_SM_Main_2__N_3496[0] ), .I1(n19702), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3493[1] ), .O(n9639));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5173_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i5174_3_lut (.I0(n9639), .I1(\r_SM_Main_2__N_3493[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n9640));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5174_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1542864_i1_3_lut (.I0(n32038), .I1(n32110), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3524));
    defparam i1542864_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3524), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n32107));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n32107_bdd_4_lut (.I0(n32107), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n32110));
    defparam n32107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3493[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_26247 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n32035));
    defparam r_Bit_Index_0__bdd_4_lut_26247.LUT_INIT = 16'he4aa;
    SB_LUT4 n32035_bdd_4_lut (.I0(n32035), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n32038));
    defparam n32035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n11634), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3878), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[3]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n29690));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n29690), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3493[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26049_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3493[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n15626));
    defparam i26049_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n15730));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1197__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n1), .D(n41[1]), .R(n15626));   // verilog/uart_tx.v(118[34:51])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n32553));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n15722));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i7001_2_lut_3_lut (.I0(\r_SM_Main_2__N_3493[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_3878));
    defparam i7001_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 r_Clock_Count_1197_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n24022), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1197_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n24021), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1197_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY r_Clock_Count_1197_add_4_9 (.CI(n24021), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n24022));
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n15548, clk32MHz, n15643, GND_net, VCC_net, \r_SM_Main_2__N_3422[2] , 
            r_SM_Main, n27820, r_Rx_Data, n19238, n4, n4_adj_1, 
            \r_Bit_Index[0] , n14287, RX_N_2, n14282, n4_adj_2, n27405, 
            rx_data_ready, n15764, n16203, rx_data, n15712, n15711, 
            n15710, n15709, n15708, n15707, n15706) /* synthesis syn_module_defined=1 */ ;
    output n15548;
    input clk32MHz;
    output n15643;
    input GND_net;
    input VCC_net;
    output \r_SM_Main_2__N_3422[2] ;
    output [2:0]r_SM_Main;
    input n27820;
    output r_Rx_Data;
    output n19238;
    output n4;
    output n4_adj_1;
    output \r_Bit_Index[0] ;
    output n14287;
    input RX_N_2;
    output n14282;
    output n4_adj_2;
    input n27405;
    output rx_data_ready;
    input n15764;
    input n16203;
    output [7:0]rx_data;
    input n15712;
    input n15711;
    input n15710;
    input n15709;
    input n15708;
    input n15707;
    input n15706;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [7:0]n37;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n24014, n24013, n24012, n24011, n24010, n24009, n24008;
    wire [2:0]r_SM_Main_2__N_3428;
    
    wire n31153, n19789, n14177, n3, r_Rx_Data_R, n28737, n15624, 
        n6, n15509, n27862, n19696, n10, n30355, n19723, n1;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n15548), 
            .D(n326[2]), .R(n15643));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n15548), 
            .D(n326[1]), .R(n15643));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1195_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n24014), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1195_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n24013), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1195_add_4_8 (.CI(n24013), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n24014));
    SB_LUT4 r_Clock_Count_1195_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n24012), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1195_add_4_7 (.CI(n24012), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n24013));
    SB_LUT4 r_Clock_Count_1195_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n24011), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1195_add_4_6 (.CI(n24011), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n24012));
    SB_LUT4 r_Clock_Count_1195_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n24010), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1195_add_4_5 (.CI(n24010), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n24011));
    SB_LUT4 r_Clock_Count_1195_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n24009), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1195_add_4_4 (.CI(n24009), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n24010));
    SB_LUT4 r_Clock_Count_1195_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n24008), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1195_add_4_3 (.CI(n24008), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n24009));
    SB_LUT4 r_Clock_Count_1195_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1195_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1195_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n24008));
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(\r_SM_Main_2__N_3422[2] ), 
            .R(n27820));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i25503_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3428[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n31153));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i25503_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n31153), .I1(\r_SM_Main_2__N_3422[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n19789));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i14710_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n19238));
    defparam i14710_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_119_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_119_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_121_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_121_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(n14177), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n14287));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_2));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i22913_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_3428[0]), 
            .I3(GND_net), .O(n28737));
    defparam i22913_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n28737), .I2(\r_SM_Main_2__N_3422[2] ), 
            .I3(r_SM_Main[1]), .O(n15624));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3428[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i26020_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n15509));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i26020_4_lut.LUT_INIT = 16'h4555;
    SB_DFFESR r_Clock_Count_1195__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n15509), .D(n37[0]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1195__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n15509), .D(n37[3]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i1266_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1266_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_845 (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27862));
    defparam i1_2_lut_adj_845.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n19696));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_846 (.I0(r_Clock_Count[3]), .I1(n27862), .I2(n10), 
            .I3(r_Clock_Count[4]), .O(\r_SM_Main_2__N_3422[2] ));
    defparam i1_4_lut_adj_846.LUT_INIT = 16'heccc;
    SB_LUT4 i11104_3_lut (.I0(n15548), .I1(n19696), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n15643));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11104_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3422[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n15548));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1273_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1273_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFFESR r_Clock_Count_1195__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n15509), .D(n37[2]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1195__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n15509), .D(n37[1]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i24524_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[4]), .O(n30355));
    defparam i24524_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut (.I0(r_Clock_Count[0]), .I1(n30355), .I2(n27862), 
            .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_3428[0]));
    defparam i6_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n19696), .I1(\r_SM_Main_2__N_3422[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n19723));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3428[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n19723), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n19789), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(\r_SM_Main_2__N_3422[2] ), .O(n14177));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_847 (.I0(\r_Bit_Index[0] ), .I1(n14177), .I2(GND_net), 
            .I3(GND_net), .O(n14282));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_847.LUT_INIT = 16'heeee;
    SB_LUT4 equal_123_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_123_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n27405));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n15764));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n16203));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1195__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n15509), .D(n37[7]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n15712));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n15711));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n15710));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n15709));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n15708));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n15707));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n15706));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1195__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n15509), .D(n37[6]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1195__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n15509), .D(n37[5]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1195__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n15509), .D(n37[4]), .R(n15624));   // verilog/uart_rx.v(120[34:51])
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (INHA_c_0, CLK_c, pwm_setpoint, 
            GND_net, \half_duty_new[0] , n1138, VCC_net, \half_duty[0][0] , 
            \half_duty[0][1] , \half_duty[0][2] , \half_duty[0][3] , \half_duty[0][4] , 
            \half_duty[0][5] , \half_duty[0][6] , \half_duty[0][7] , \half_duty_new[1] , 
            \half_duty_new[2] , \half_duty_new[3] , \half_duty_new[4] , 
            \half_duty_new[5] , \half_duty_new[6] , \half_duty_new[7] , 
            n16247, n16246, n16245, n16244, n16243, n16242, n16241, 
            n15724);
    output INHA_c_0;
    input CLK_c;
    input [22:0]pwm_setpoint;
    input GND_net;
    output \half_duty_new[0] ;
    output n1138;
    input VCC_net;
    output \half_duty[0][0] ;
    output \half_duty[0][1] ;
    output \half_duty[0][2] ;
    output \half_duty[0][3] ;
    output \half_duty[0][4] ;
    output \half_duty[0][5] ;
    output \half_duty[0][6] ;
    output \half_duty[0][7] ;
    output \half_duty_new[1] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[5] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input n16247;
    input n16246;
    input n16245;
    input n16244;
    input n16243;
    input n16242;
    input n16241;
    input n15724;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n19120, n28555;
    wire [9:0]half_duty_new_9__N_674;
    wire [22:0]n5334;
    
    wire n23857, n23858, n23856, n23855, n23854;
    wire [10:0]n49;
    
    wire pause_counter_0__N_622;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire n23853, n23852, n23851, n23850, n23849, n23848, n23847, 
        n23846, n23845, n23844, n23843, n23842, n23841, n23840, 
        n23839, n23838, n23837, n23836, n23835, n23834, n23833, 
        n23832, n23831, n23830, n23829, n23828, n23827, n23826, 
        n23825, n23824, n23823, n23822, n23821, n23820, n23819, 
        n23818, n23817, n23517, pwm_out_0__N_596, n23516, n10, n23515, 
        n9, n23514, n8;
    wire [10:0]pwm_out_0__N_597;
    
    wire n23513, n7, n23512, n6, n23511, n5, n23510, n4, n23509, 
        n3, n23508, n2, n23507, n1, n27545, pause_counter_0, n20, 
        n19, n6_adj_3872, n23984, n23983, n23982, n23981, n23980, 
        n23979, n23978, n23977, n23976, n23975, n14, n22, n21, 
        n23, n15, n14_adj_3873, n20_adj_3874, n18, n19_adj_3875, 
        n17, n23859;
    
    SB_DFFE pwm_out_0__39 (.Q(INHA_c_0), .C(CLK_c), .E(n28555), .D(n19120));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 add_1623_22_lut (.I0(GND_net), .I1(n5334[20]), .I2(pwm_setpoint[20]), 
            .I3(n23857), .O(half_duty_new_9__N_674[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1623_22 (.CI(n23857), .I0(n5334[20]), .I1(pwm_setpoint[20]), 
            .CO(n23858));
    SB_LUT4 add_1623_21_lut (.I0(GND_net), .I1(n5334[19]), .I2(pwm_setpoint[19]), 
            .I3(n23856), .O(half_duty_new_9__N_674[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1623_21 (.CI(n23856), .I0(n5334[19]), .I1(pwm_setpoint[19]), 
            .CO(n23857));
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_674[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 add_1623_20_lut (.I0(GND_net), .I1(n5334[18]), .I2(pwm_setpoint[18]), 
            .I3(n23855), .O(half_duty_new_9__N_674[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1623_20 (.CI(n23855), .I0(n5334[18]), .I1(pwm_setpoint[18]), 
            .CO(n23856));
    SB_LUT4 add_1623_19_lut (.I0(GND_net), .I1(n5334[17]), .I2(pwm_setpoint[17]), 
            .I3(n23854), .O(half_duty_new_9__N_674[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR count_0__1192__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[7]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY add_1623_19 (.CI(n23854), .I0(n5334[17]), .I1(pwm_setpoint[17]), 
            .CO(n23855));
    SB_DFFESR count_0__1192__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[6]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1192__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[5]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 add_1623_18_lut (.I0(GND_net), .I1(n5334[16]), .I2(pwm_setpoint[16]), 
            .I3(n23853), .O(half_duty_new_9__N_674[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1623_18 (.CI(n23853), .I0(n5334[16]), .I1(pwm_setpoint[16]), 
            .CO(n23854));
    SB_LUT4 add_1623_17_lut (.I0(GND_net), .I1(n5334[15]), .I2(pwm_setpoint[15]), 
            .I3(n23852), .O(half_duty_new_9__N_674[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1623_17 (.CI(n23852), .I0(n5334[15]), .I1(pwm_setpoint[15]), 
            .CO(n23853));
    SB_CARRY add_1623_16 (.CI(n23851), .I0(n5334[14]), .I1(pwm_setpoint[14]), 
            .CO(n23852));
    SB_CARRY add_1623_15 (.CI(n23850), .I0(n5334[13]), .I1(pwm_setpoint[13]), 
            .CO(n23851));
    SB_CARRY add_1623_14 (.CI(n23849), .I0(n5334[12]), .I1(pwm_setpoint[12]), 
            .CO(n23850));
    SB_CARRY add_1623_13 (.CI(n23848), .I0(n5334[11]), .I1(pwm_setpoint[11]), 
            .CO(n23849));
    SB_CARRY add_1623_12 (.CI(n23847), .I0(n5334[10]), .I1(pwm_setpoint[10]), 
            .CO(n23848));
    SB_CARRY add_1623_11 (.CI(n23846), .I0(n5334[9]), .I1(pwm_setpoint[9]), 
            .CO(n23847));
    SB_CARRY add_1623_10 (.CI(n23845), .I0(n5334[8]), .I1(pwm_setpoint[8]), 
            .CO(n23846));
    SB_CARRY add_1623_9 (.CI(n23844), .I0(n5334[7]), .I1(pwm_setpoint[7]), 
            .CO(n23845));
    SB_CARRY add_1623_8 (.CI(n23843), .I0(n5334[6]), .I1(pwm_setpoint[6]), 
            .CO(n23844));
    SB_CARRY add_1623_7 (.CI(n23842), .I0(n5334[5]), .I1(pwm_setpoint[5]), 
            .CO(n23843));
    SB_CARRY add_1623_6 (.CI(n23841), .I0(n5334[4]), .I1(pwm_setpoint[4]), 
            .CO(n23842));
    SB_CARRY add_1623_5 (.CI(n23840), .I0(n5334[3]), .I1(pwm_setpoint[3]), 
            .CO(n23841));
    SB_CARRY add_1623_4 (.CI(n23839), .I0(n5334[2]), .I1(pwm_setpoint[2]), 
            .CO(n23840));
    SB_CARRY add_1623_3 (.CI(n23838), .I0(n5334[1]), .I1(pwm_setpoint[1]), 
            .CO(n23839));
    SB_CARRY add_1623_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n23838));
    SB_LUT4 add_1630_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n23837), .O(n5334[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1630_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n23836), .O(n5334[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_22 (.CI(n23836), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n23837));
    SB_LUT4 add_1630_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n23835), .O(n5334[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_21 (.CI(n23835), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n23836));
    SB_LUT4 add_1630_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n23834), .O(n5334[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_20 (.CI(n23834), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n23835));
    SB_LUT4 add_1630_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n23833), .O(n5334[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_19 (.CI(n23833), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n23834));
    SB_LUT4 add_1630_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n23832), .O(n5334[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_18 (.CI(n23832), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n23833));
    SB_LUT4 add_1630_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n23831), .O(n5334[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_17 (.CI(n23831), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n23832));
    SB_LUT4 add_1630_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n23830), .O(n5334[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_16 (.CI(n23830), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n23831));
    SB_LUT4 add_1630_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n23829), .O(n5334[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_15 (.CI(n23829), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n23830));
    SB_LUT4 add_1630_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n23828), .O(n5334[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_14 (.CI(n23828), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n23829));
    SB_LUT4 add_1630_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n23827), .O(n5334[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_13 (.CI(n23827), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n23828));
    SB_LUT4 add_1630_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n23826), .O(n5334[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_12 (.CI(n23826), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n23827));
    SB_LUT4 add_1630_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n23825), .O(n5334[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_11 (.CI(n23825), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n23826));
    SB_LUT4 add_1630_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n23824), .O(n5334[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_10 (.CI(n23824), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n23825));
    SB_LUT4 add_1630_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n23823), .O(n5334[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_9 (.CI(n23823), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n23824));
    SB_LUT4 add_1630_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n23822), .O(n5334[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_8 (.CI(n23822), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n23823));
    SB_LUT4 add_1630_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n23821), .O(n5334[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_7 (.CI(n23821), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n23822));
    SB_LUT4 add_1630_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n23820), .O(n5334[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_6 (.CI(n23820), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n23821));
    SB_LUT4 add_1630_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n23819), .O(n5334[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_5 (.CI(n23819), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n23820));
    SB_LUT4 add_1630_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n23818), .O(n5334[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_4 (.CI(n23818), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n23819));
    SB_LUT4 add_1630_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n23817), .O(n5334[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_3 (.CI(n23817), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n23818));
    SB_LUT4 add_1630_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5334[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1630_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1630_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n23817));
    SB_DFFESR count_0__1192__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[4]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1192__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[3]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1192__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[2]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1192__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[1]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY pwm_out_0__I_20_13 (.CI(n23517), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_596));
    SB_CARRY pwm_out_0__I_20_12 (.CI(n23516), .I0(VCC_net), .I1(VCC_net), 
            .CO(n23517));
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n23515), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_11 (.CI(n23515), .I0(VCC_net), .I1(VCC_net), 
            .CO(n23516));
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n23514), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_10 (.CI(n23514), .I0(GND_net), .I1(VCC_net), 
            .CO(n23515));
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_597[7]), 
            .I3(n23513), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_9 (.CI(n23513), .I0(GND_net), .I1(pwm_out_0__N_597[7]), 
            .CO(n23514));
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_597[6]), 
            .I3(n23512), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n23512), .I0(VCC_net), .I1(pwm_out_0__N_597[6]), 
            .CO(n23513));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_597[5]), 
            .I3(n23511), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_7 (.CI(n23511), .I0(GND_net), .I1(pwm_out_0__N_597[5]), 
            .CO(n23512));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_597[4]), 
            .I3(n23510), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_6 (.CI(n23510), .I0(GND_net), .I1(pwm_out_0__N_597[4]), 
            .CO(n23511));
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_597[3]), 
            .I3(n23509), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_5 (.CI(n23509), .I0(GND_net), .I1(pwm_out_0__N_597[3]), 
            .CO(n23510));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_597[2]), 
            .I3(n23508), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_4 (.CI(n23508), .I0(GND_net), .I1(pwm_out_0__N_597[2]), 
            .CO(n23509));
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_597[1]), 
            .I3(n23507), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_3 (.CI(n23507), .I0(GND_net), .I1(pwm_out_0__N_597[1]), 
            .CO(n23508));
    SB_DFFESR count_0__1192__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[8]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_597[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_597[0]), 
            .CO(n23507));
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n27545));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1192__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[0]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 i8_4_lut (.I0(\count[0] [6]), .I1(\count[0] [0]), .I2(\count[0] [10]), 
            .I3(\count[0] [1]), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i7_4_lut (.I0(pause_counter_0), .I1(\count[0] [9]), .I2(\count[0] [8]), 
            .I3(\count[0] [7]), .O(n19));
    defparam i7_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut (.I0(\count[0] [4]), .I1(n19), .I2(n20), .I3(GND_net), 
            .O(n6_adj_3872));
    defparam i1_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i4_4_lut (.I0(\count[0] [5]), .I1(\count[0] [2]), .I2(\count[0] [3]), 
            .I3(n6_adj_3872), .O(n1138));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_622));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22794_1_lut (.I0(n19120), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n27545));
    defparam i22794_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 count_0__1192_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n23984), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1192_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n23983), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0][5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i7_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[6]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY count_0__1192_add_4_11 (.CI(n23983), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n23984));
    SB_LUT4 count_0__1192_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n23982), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_10 (.CI(n23982), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n23983));
    SB_LUT4 count_0__1192_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n23981), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_9 (.CI(n23981), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n23982));
    SB_LUT4 count_0__1192_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n23980), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_8 (.CI(n23980), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n23981));
    SB_LUT4 count_0__1192_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n23979), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_7 (.CI(n23979), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n23980));
    SB_LUT4 count_0__1192_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n23978), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_6 (.CI(n23978), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n23979));
    SB_LUT4 count_0__1192_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n23977), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_5 (.CI(n23977), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n23978));
    SB_LUT4 count_0__1192_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n23976), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_4 (.CI(n23976), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n23977));
    SB_LUT4 count_0__1192_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n23975), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_3 (.CI(n23975), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n23976));
    SB_DFFESR count_0__1192__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[10]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_674[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_674[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_674[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_674[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(\half_duty_new[5] ), .C(CLK_c), .D(half_duty_new_9__N_674[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_674[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_674[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 count_0__1192_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1192_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1192_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n23975));
    SB_DFFESR count_0__1192__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_622), 
            .D(n49[9]), .R(n1138));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 i1_2_lut (.I0(n6), .I1(pause_counter_0), .I2(GND_net), .I3(GND_net), 
            .O(n14));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(n4), .I1(n7), .I2(n5), .I3(n10), .O(n22));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_843 (.I0(\count[0] [10]), .I1(n9), .I2(n8), .I3(n2), 
            .O(n21));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i8_4_lut_adj_843.LUT_INIT = 16'hfffd;
    SB_LUT4 i10_4_lut (.I0(n1), .I1(pwm_out_0__N_596), .I2(n3), .I3(n14), 
            .O(n23));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i10_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i26015_4_lut (.I0(n23), .I1(n19120), .I2(n21), .I3(n22), 
            .O(n28555));
    defparam i26015_4_lut.LUT_INIT = 16'h3337;
    SB_LUT4 i3_4_lut (.I0(\half_duty[0][5] ), .I1(\half_duty[0][7] ), .I2(\count[0] [5]), 
            .I3(\count[0] [7]), .O(n15));
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut (.I0(\count[0] [10]), .I1(\half_duty[0][6] ), .I2(\count[0] [6]), 
            .I3(GND_net), .O(n14_adj_3873));
    defparam i2_3_lut.LUT_INIT = 16'hbebe;
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n16247));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n16246));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0][5] ), .C(CLK_c), .D(n16245));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n16244));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n16243));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n16242));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n16241));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i8_3_lut (.I0(n15), .I1(\count[0] [9]), .I2(\count[0] [8]), 
            .I3(GND_net), .O(n20_adj_3874));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(\half_duty[0][0] ), .I1(\half_duty[0][4] ), .I2(\count[0] [0]), 
            .I3(\count[0] [4]), .O(n18));
    defparam i6_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_844 (.I0(\half_duty[0][3] ), .I1(n14_adj_3873), 
            .I2(pause_counter_0), .I3(\count[0] [3]), .O(n19_adj_3875));
    defparam i7_4_lut_adj_844.LUT_INIT = 16'hfdfe;
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n15724));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i5_4_lut (.I0(\half_duty[0][2] ), .I1(\half_duty[0][1] ), .I2(\count[0] [2]), 
            .I3(\count[0] [1]), .O(n17));
    defparam i5_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i11_4_lut (.I0(n17), .I1(n19_adj_3875), .I2(n18), .I3(n20_adj_3874), 
            .O(n19120));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_1623_24_lut (.I0(GND_net), .I1(n5334[22]), .I2(pwm_setpoint[22]), 
            .I3(n23859), .O(half_duty_new_9__N_674[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1623_23_lut (.I0(GND_net), .I1(n5334[21]), .I2(pwm_setpoint[21]), 
            .I3(n23858), .O(half_duty_new_9__N_674[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1623_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1623_23 (.CI(n23858), .I0(n5334[21]), .I1(pwm_setpoint[21]), 
            .CO(n23859));
    
endmodule
